module c7552 (N1, N5, N9, N12, N15, N18, N23, N26, N29, N32, N35, N38, N41, N44, N47, N50, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N69, N70, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N94, N97, N100, N103, N106, N109, N110, N111, N112, N113, N114, N115, N118, N121, N124, N127, N130, N133, N134, N135, N138, N141, N144, N147, N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241, N242, N245, N248, N251, N254, N257, N260, N263, N267, N271, N274, N277, N280, N283, N286, N289, N293, N296, N299, N303, N307, N310, N313, N316, N319, N322, N325, N328, N331, N334, N337, N340, N343, N346, N349, N352, N355, N358, N361, N364, N367, N382, B241, N387, N388, N478, N482, N484, N486, N489, N492, N501, N505, N507, N509, N511, N513, N515, N517, N519, N535, N537, N539, N541, N543, N545, N547, N549, N551, N553, N556, N559, N561, N563, N565, N567, N569, N571, N573, N582, N643, N707, N813, N881, N882, N883, N884, N885, N889, N945, N1110, N1111, N1112, N1113, N1114, N1489, N1490, N1781, N10025, N10101, N10102, N10103, N10104, N10109, N10110, N10111, N10112, N10350, N10351, N10352, N10353, N10574, N10575, N10576, N10628, N10632, N10641, N10704, N10706, N10711, N10712, N10713, N10714, N10715, N10716, N10717, N10718, N10729, N10759, N10760, N10761, N10762, N10763, N10827, N10837, N10838, N10839, N10840, N10868, N10869, N10870, N10871, N10905, N10906, N10907, N10908, N11333, N11334, N11340, N11342);

input N1, N5, N9, N12, N15, N18, N23, N26, N29, N32, N35, N38, N41, N44, N47, N50, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N69, N70, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N94, N97, N100, N103, N106, N109, N110, N111, N112, N113, N114, N115, N118, N121, N124, N127, N130, N133, N134, N135, N138, N141, N144, N147, N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241, N242, N245, N248, N251, N254, N257, N260, N263, N267, N271, N274, N277, N280, N283, N286, N289, N293, N296, N299, N303, N307, N310, N313, N316, N319, N322, N325, N328, N331, N334, N337, N340, N343, N346, N349, N352, N355, N358, N361, N364, N367, N382;

output B241, N387, N388, N478, N482, N484, N486, N489, N492, N501, N505, N507, N509, N511, N513, N515, N517, N519, N535, N537, N539, N541, N543, N545, N547, N549, N551, N553, N556, N559, N561, N563, N565, N567, N569, N571, N573, N582, N643, N707, N813, N881, N882, N883, N884, N885, N889, N945, N1110, N1111, N1112, N1113, N1114, N1489, N1490, N1781, N10025, N10101, N10102, N10103, N10104, N10109, N10110, N10111, N10112, N10350, N10351, N10352, N10353, N10574, N10575, N10576, N10628, N10632, N10641, N10704, N10706, N10711, N10712, N10713, N10714, N10715, N10716, N10717, N10718, N10729, N10759, N10760, N10761, N10762, N10763, N10827, N10837, N10838, N10839, N10840, N10868, N10869, N10870, N10871, N10905, N10906, N10907, N10908, N11333, N11334, N11340, N11342;

wire N467,N469,N494,N528,N575,N578,N585,N590,N593,N596,N599,N604,N609,N614,N625,N628,N632,N636,N641,N642,N644,N651,N657,N660,N666,N672,N673,N674,N676,N682,N688,N689,N695,N700,N705,N706,N708,N715,N721,N727,N733,N734,N742,N748,N749,N750,N758,N759,N762,N768,N774,N780,N786,N794,N800,N806,N812,N814,N821,N827,N833,N839,N845,N853,N859,N865,N871,N886,N887,N957,N1028,N1029,N1109,N1115,N1116,N1119,N1125,N1132,N1136,N1141,N1147,N1154,N1160,N1167,N1174,N1175,N1182,N1189,N1194,N1199,N1206,N1211,N1218,N1222,N1227,N1233,N1240,N1244,N1249,N1256,N1263,N1270,N1277,N1284,N1287,N1290,N1293,N1296,N1299,N1302,N1305,N1308,N1311,N1314,N1317,N1320,N1323,N1326,N1329,N1332,N1335,N1338,N1341,N1344,N1347,N1350,N1353,N1356,N1359,N1362,N1365,N1368,N1371,N1374,N1377,N1380,N1383,N1386,N1389,N1392,N1395,N1398,N1401,N1404,N1407,N1410,N1413,N1416,N1419,N1422,N1425,N1428,N1431,N1434,N1437,N1440,N1443,N1446,N1449,N1452,N1455,N1458,N1461,N1464,N1467,N1470,N1473,N1476,N1479,N1482,N1485,N1537,N1551,N1649,N1703,N1708,N1713,N1721,N1758,N1782,N1783,N1789,N1793,N1794,N1795,N1796,N1797,N1798,N1799,N1805,N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,N1819,N1820,N1821,N1822,N1828,N1829,N1830,N1832,N1833,N1834,N1835,N1839,N1840,N1841,N1842,N1843,N1845,N1851,N1857,N1858,N1859,N1860,N1861,N1862,N1863,N1864,N1865,N1866,N1867,N1868,N1869,N1870,N1871,N1872,N1873,N1874,N1875,N1876,N1877,N1878,N1879,N1880,N1881,N1882,N1883,N1884,N1885,N1892,N1899,N1906,N1913,N1919,N1926,N1927,N1928,N1929,N1930,N1931,N1932,N1933,N1934,N1935,N1936,N1937,N1938,N1939,N1940,N1941,N1942,N1943,N1944,N1945,N1946,N1947,N1953,N1957,N1958,N1959,N1960,N1961,N1962,N1963,N1965,N1966,N1967,N1968,N1969,N1970,N1971,N1972,N1973,N1974,N1975,N1976,N1977,N1983,N1989,N1990,N1991,N1992,N1993,N1994,N1995,N1996,N1997,N2003,N2010,N2011,N2012,N2013,N2014,N2015,N2016,N2017,N2018,N2019,N2020,N2021,N2022,N2023,N2024,N2031,N2038,N2045,N2052,N2058,N2064,N2065,N2066,N2067,N2068,N2069,N2070,N2071,N2072,N2073,N2074,N2081,N2086,N2107,N2108,N2110,N2111,N2112,N2113,N2114,N2115,N2117,N2171,N2172,N2230,N2231,N2235,N2239,N2240,N2241,N2242,N2243,N2244,N2245,N2246,N2247,N2248,N2249,N2250,N2251,N2252,N2253,N2254,N2255,N2256,N2257,N2267,N2268,N2269,N2274,N2275,N2277,N2278,N2279,N2280,N2281,N2282,N2283,N2284,N2285,N2286,N2287,N2293,N2299,N2300,N2301,N2302,N2303,N2304,N2305,N2306,N2307,N2308,N2309,N2315,N2321,N2322,N2323,N2324,N2325,N2326,N2327,N2328,N2329,N2330,N2331,N2337,N2338,N2339,N2340,N2341,N2342,N2343,N2344,N2345,N2346,N2347,N2348,N2349,N2350,N2351,N2352,N2353,N2354,N2355,N2356,N2357,N2358,N2359,N2360,N2361,N2362,N2363,N2364,N2365,N2366,N2367,N2368,N2374,N2375,N2376,N2377,N2378,N2379,N2380,N2381,N2382,N2383,N2384,N2390,N2396,N2397,N2398,N2399,N2400,N2401,N2402,N2403,N2404,N2405,N2406,N2412,N2418,N2419,N2420,N2421,N2422,N2423,N2424,N2425,N2426,N2427,N2428,N2429,N2430,N2431,N2432,N2433,N2434,N2435,N2436,N2437,N2441,N2442,N2446,N2450,N2454,N2458,N2462,N2466,N2470,N2474,N2478,N2482,N2488,N2496,N2502,N2508,N2523,N2533,N2537,N2538,N2542,N2546,N2550,N2554,N2561,N2567,N2573,N2604,N2607,N2611,N2615,N2619,N2626,N2632,N2638,N2644,N2650,N2653,N2654,N2658,N2662,N2666,N2670,N2674,N2680,N2688,N2692,N2696,N2700,N2704,N2728,N2729,N2733,N2737,N2741,N2745,N2749,N2753,N2757,N2761,N2765,N2766,N2769,N2772,N2775,N2778,N2781,N2784,N2787,N2790,N2793,N2796,N2866,N2867,N2868,N2869,N2878,N2913,N2914,N2915,N2916,N2917,N2918,N2919,N2920,N2921,N2922,N2923,N2924,N2925,N2926,N2927,N2928,N2929,N2930,N2931,N2932,N2933,N2934,N2935,N2936,N2937,N2988,N3005,N3006,N3007,N3008,N3009,N3020,N3021,N3022,N3023,N3024,N3025,N3026,N3027,N3028,N3029,N3032,N3033,N3034,N3035,N3036,N3037,N3038,N3039,N3040,N3041,N3061,N3064,N3067,N3070,N3073,N3080,N3096,N3097,N3101,N3107,N3114,N3122,N3126,N3130,N3131,N3134,N3135,N3136,N3137,N3140,N3144,N3149,N3155,N3159,N3167,N3168,N3169,N3173,N3178,N3184,N3185,N3189,N3195,N3202,N3210,N3211,N3215,N3221,N3228,N3229,N3232,N3236,N3241,N3247,N3251,N3255,N3259,N3263,N3267,N3273,N3281,N3287,N3293,N3299,N3303,N3307,N3311,N3315,N3322,N3328,N3334,N3340,N3343,N3349,N3355,N3361,N3362,N3363,N3364,N3365,N3366,N3367,N3368,N3369,N3370,N3371,N3372,N3373,N3374,N3375,N3379,N3380,N3381,N3384,N3390,N3398,N3404,N3410,N3416,N3420,N3424,N3428,N3432,N3436,N3440,N3444,N3448,N3452,N3453,N3454,N3458,N3462,N3466,N3470,N3474,N3478,N3482,N3486,N3487,N3490,N3493,N3496,N3499,N3502,N3507,N3510,N3515,N3518,N3521,N3524,N3527,N3530,N3535,N3539,N3542,N3545,N3548,N3551,N3552,N3553,N3557,N3560,N3563,N3566,N3569,N3570,N3571,N3574,N3577,N3580,N3583,N3586,N3589,N3592,N3595,N3598,N3601,N3604,N3607,N3610,N3613,N3616,N3619,N3622,N3625,N3628,N3631,N3634,N3637,N3640,N3643,N3646,N3649,N3652,N3655,N3658,N3661,N3664,N3667,N3670,N3673,N3676,N3679,N3682,N3685,N3688,N3691,N3694,N3697,N3700,N3703,N3706,N3709,N3712,N3715,N3718,N3721,N3724,N3727,N3730,N3733,N3736,N3739,N3742,N3745,N3748,N3751,N3754,N3757,N3760,N3763,N3766,N3769,N3772,N3775,N3778,N3781,N3782,N3783,N3786,N3789,N3792,N3795,N3798,N3801,N3804,N3807,N3810,N3813,N3816,N3819,N3822,N3825,N3828,N3831,N3834,N3837,N3840,N3843,N3846,N3849,N3852,N3855,N3858,N3861,N3864,N3867,N3870,N3873,N3876,N3879,N3882,N3885,N3888,N3891,N3953,N3954,N3955,N3956,N3958,N3964,N4193,N4303,N4308,N4313,N4326,N4327,N4333,N4334,N4411,N4412,N4463,N4464,N4465,N4466,N4467,N4468,N4469,N4470,N4471,N4472,N4473,N4474,N4475,N4476,N4477,N4478,N4479,N4480,N4481,N4482,N4483,N4484,N4485,N4486,N4487,N4488,N4489,N4490,N4491,N4492,N4493,N4494,N4495,N4496,N4497,N4498,N4499,N4500,N4501,N4502,N4503,N4504,N4505,N4506,N4507,N4508,N4509,N4510,N4511,N4512,N4513,N4514,N4515,N4516,N4517,N4518,N4519,N4520,N4521,N4522,N4523,N4524,N4525,N4526,N4527,N4528,N4529,N4530,N4531,N4532,N4533,N4534,N4535,N4536,N4537,N4538,N4539,N4540,N4541,N4542,N4543,N4544,N4545,N4549,N4555,N4562,N4563,N4566,N4570,N4575,N4576,N4577,N4581,N4586,N4592,N4593,N4597,N4603,N4610,N4611,N4612,N4613,N4614,N4615,N4616,N4617,N4618,N4619,N4620,N4621,N4622,N4623,N4624,N4625,N4626,N4627,N4628,N4629,N4630,N4631,N4632,N4633,N4634,N4635,N4636,N4637,N4638,N4639,N4640,N4641,N4642,N4643,N4644,N4645,N4646,N4647,N4648,N4649,N4650,N4651,N4652,N4653,N4656,N4657,N4661,N4667,N4674,N4675,N4678,N4682,N4687,N4693,N4694,N4695,N4696,N4697,N4698,N4699,N4700,N4701,N4702,N4706,N4711,N4717,N4718,N4722,N4728,N4735,N4743,N4744,N4745,N4746,N4747,N4748,N4749,N4750,N4751,N4752,N4753,N4754,N4755,N4756,N4757,N4758,N4759,N4760,N4761,N4762,N4763,N4764,N4765,N4766,N4767,N4768,N4769,N4775,N4776,N4777,N4778,N4779,N4780,N4781,N4782,N4783,N4784,N4789,N4790,N4793,N4794,N4795,N4796,N4799,N4800,N4801,N4802,N4803,N4806,N4809,N4810,N4813,N4814,N4817,N4820,N4823,N4826,N4829,N4832,N4835,N4838,N4841,N4844,N4847,N4850,N4853,N4856,N4859,N4862,N4865,N4868,N4871,N4874,N4877,N4880,N4883,N4886,N4889,N4892,N4895,N4898,N4901,N4904,N4907,N4910,N4913,N4916,N4919,N4922,N4925,N4928,N4931,N4934,N4937,N4940,N4943,N4946,N4949,N4952,N4955,N4958,N4961,N4964,N4967,N4970,N4973,N4976,N4979,N4982,N4985,N4988,N4991,N4994,N4997,N5000,N5003,N5006,N5009,N5012,N5015,N5018,N5021,N5024,N5027,N5030,N5033,N5036,N5039,N5042,N5045,N5046,N5047,N5048,N5049,N5052,N5055,N5058,N5061,N5064,N5065,N5066,N5067,N5068,N5071,N5074,N5077,N5080,N5083,N5086,N5089,N5092,N5095,N5098,N5101,N5104,N5107,N5110,N5111,N5112,N5113,N5114,N5117,N5120,N5123,N5126,N5129,N5132,N5135,N5138,N5141,N5144,N5147,N5150,N5153,N5156,N5159,N5162,N5165,N5166,N5167,N5168,N5169,N5170,N5171,N5172,N5173,N5174,N5175,N5176,N5177,N5178,N5179,N5180,N5181,N5182,N5183,N5184,N5185,N5186,N5187,N5188,N5189,N5190,N5191,N5192,N5193,N5196,N5197,N5198,N5199,N5200,N5201,N5202,N5203,N5204,N5205,N5206,N5207,N5208,N5209,N5210,N5211,N5212,N5213,N5283,N5284,N5285,N5286,N5287,N5288,N5289,N5290,N5291,N5292,N5293,N5294,N5295,N5296,N5297,N5298,N5299,N5300,N5314,N5315,N5316,N5317,N5318,N5319,N5320,N5321,N5322,N5323,N5324,N5363,N5364,N5365,N5366,N5367,N5425,N5426,N5427,N5429,N5430,N5431,N5432,N5433,N5451,N5452,N5453,N5454,N5455,N5456,N5457,N5469,N5474,N5475,N5476,N5477,N5571,N5572,N5573,N5574,N5584,N5585,N5586,N5587,N5602,N5603,N5604,N5605,N5631,N5632,N5640,N5654,N5670,N5683,N5690,N5697,N5707,N5718,N5728,N5735,N5736,N5740,N5744,N5747,N5751,N5755,N5758,N5762,N5766,N5769,N5770,N5771,N5778,N5789,N5799,N5807,N5821,N5837,N5850,N5856,N5863,N5870,N5881,N5892,N5898,N5905,N5915,N5926,N5936,N5943,N5944,N5945,N5946,N5947,N5948,N5949,N5950,N5951,N5952,N5953,N5954,N5955,N5956,N5957,N5958,N5959,N5960,N5966,N5967,N5968,N5969,N5970,N5971,N5972,N5973,N5974,N5975,N5976,N5977,N5978,N5979,N5980,N5981,N5989,N5990,N5991,N5996,N6000,N6003,N6009,N6014,N6018,N6021,N6022,N6023,N6024,N6025,N6026,N6027,N6028,N6029,N6030,N6031,N6032,N6033,N6034,N6035,N6036,N6037,N6038,N6039,N6040,N6041,N6047,N6052,N6056,N6059,N6060,N6061,N6062,N6063,N6064,N6065,N6066,N6067,N6068,N6069,N6070,N6071,N6072,N6073,N6074,N6075,N6076,N6077,N6078,N6079,N6083,N6087,N6090,N6091,N6092,N6093,N6094,N6095,N6096,N6097,N6098,N6099,N6100,N6101,N6102,N6103,N6104,N6105,N6106,N6107,N6108,N6109,N6110,N6111,N6112,N6113,N6114,N6115,N6116,N6117,N6118,N6119,N6120,N6121,N6122,N6123,N6124,N6125,N6126,N6127,N6131,N6135,N6136,N6137,N6141,N6145,N6148,N6149,N6150,N6151,N6152,N6153,N6154,N6155,N6156,N6157,N6158,N6159,N6160,N6161,N6162,N6163,N6164,N6165,N6166,N6170,N6174,N6177,N6181,N6182,N6183,N6184,N6185,N6186,N6187,N6188,N6189,N6190,N6191,N6192,N6193,N6194,N6195,N6196,N6199,N6202,N6203,N6204,N6207,N6210,N6213,N6214,N6217,N6220,N6223,N6224,N6225,N6226,N6227,N6228,N6229,N6230,N6231,N6232,N6235,N6236,N6239,N6240,N6241,N6242,N6243,N6246,N6249,N6252,N6255,N6256,N6257,N6258,N6259,N6260,N6261,N6262,N6263,N6266,N6540,N6541,N6542,N6543,N6544,N6545,N6546,N6547,N6555,N6556,N6557,N6558,N6559,N6560,N6561,N6569,N6594,N6595,N6596,N6597,N6598,N6599,N6600,N6601,N6602,N6603,N6604,N6605,N6606,N6621,N6622,N6623,N6624,N6625,N6626,N6627,N6628,N6629,N6639,N6640,N6641,N6642,N6643,N6644,N6645,N6646,N6647,N6648,N6649,N6650,N6651,N6652,N6653,N6654,N6655,N6656,N6657,N6658,N6659,N6660,N6661,N6668,N6677,N6678,N6679,N6680,N6681,N6682,N6683,N6684,N6685,N6686,N6687,N6688,N6689,N6690,N6702,N6703,N6704,N6705,N6706,N6707,N6708,N6709,N6710,N6711,N6712,N6729,N6730,N6731,N6732,N6733,N6734,N6735,N6736,N6741,N6742,N6743,N6744,N6751,N6752,N6753,N6754,N6755,N6756,N6757,N6758,N6761,N6762,N6766,N6767,N6768,N6769,N6770,N6771,N6772,N6773,N6774,N6775,N6776,N6777,N6778,N6779,N6780,N6781,N6782,N6783,N6784,N6787,N6788,N6789,N6790,N6791,N6792,N6793,N6794,N6795,N6796,N6797,N6800,N6803,N6806,N6809,N6812,N6815,N6818,N6821,N6824,N6827,N6830,N6833,N6836,N6837,N6838,N6839,N6840,N6841,N6842,N6843,N6844,N6845,N6848,N6849,N6850,N6851,N6852,N6853,N6854,N6855,N6856,N6857,N6858,N6859,N6860,N6861,N6862,N6863,N6864,N6865,N6866,N6867,N6870,N6871,N6872,N6873,N6874,N6875,N6876,N6877,N6878,N6879,N6880,N6881,N6884,N6885,N6886,N6887,N6888,N6889,N6890,N6891,N6892,N6893,N6894,N6901,N6912,N6923,N6929,N6936,N6946,N6957,N6967,N6968,N6969,N6970,N6977,N6988,N6998,N7006,N7020,N7036,N7049,N7055,N7056,N7057,N7060,N7061,N7062,N7063,N7064,N7065,N7066,N7067,N7068,N7073,N7077,N7080,N7086,N7091,N7095,N7098,N7099,N7100,N7103,N7104,N7105,N7106,N7107,N7114,N7125,N7136,N7142,N7149,N7159,N7170,N7180,N7187,N7188,N7191,N7194,N7198,N7202,N7205,N7209,N7213,N7216,N7219,N7222,N7229,N7240,N7250,N7258,N7272,N7288,N7301,N7307,N7314,N7318,N7322,N7325,N7328,N7331,N7334,N7337,N7340,N7343,N7346,N7351,N7355,N7358,N7364,N7369,N7373,N7376,N7377,N7378,N7381,N7384,N7387,N7391,N7394,N7398,N7402,N7405,N7408,N7411,N7414,N7417,N7420,N7423,N7426,N7429,N7432,N7435,N7438,N7441,N7444,N7447,N7450,N7453,N7456,N7459,N7462,N7465,N7468,N7471,N7474,N7477,N7478,N7479,N7482,N7485,N7488,N7491,N7494,N7497,N7500,N7503,N7506,N7509,N7512,N7515,N7518,N7521,N7524,N7527,N7530,N7533,N7536,N7539,N7542,N7545,N7548,N7551,N7552,N7553,N7556,N7557,N7558,N7559,N7560,N7563,N7566,N7569,N7572,N7573,N7574,N7577,N7580,N7581,N7582,N7585,N7588,N7591,N7609,N7613,N7620,N7649,N7650,N7655,N7659,N7668,N7671,N7744,N7822,N7825,N7826,N7852,N8114,N8117,N8131,N8134,N8144,N8145,N8146,N8156,N8166,N8169,N8183,N8186,N8196,N8200,N8204,N8208,N8216,N8217,N8218,N8219,N8232,N8233,N8242,N8243,N8244,N8245,N8246,N8247,N8248,N8249,N8250,N8251,N8252,N8253,N8254,N8260,N8261,N8262,N8269,N8274,N8275,N8276,N8277,N8278,N8279,N8280,N8281,N8282,N8283,N8284,N8285,N8288,N8294,N8295,N8296,N8297,N8298,N8307,N8315,N8317,N8319,N8321,N8322,N8323,N8324,N8325,N8326,N8333,N8337,N8338,N8339,N8340,N8341,N8342,N8343,N8344,N8345,N8346,N8347,N8348,N8349,N8350,N8351,N8352,N8353,N8354,N8355,N8356,N8357,N8358,N8365,N8369,N8370,N8371,N8372,N8373,N8374,N8375,N8376,N8377,N8378,N8379,N8380,N8381,N8382,N8383,N8384,N8385,N8386,N8387,N8388,N8389,N8390,N8391,N8392,N8393,N8394,N8404,N8405,N8409,N8410,N8411,N8412,N8415,N8416,N8417,N8418,N8421,N8430,N8433,N8434,N8435,N8436,N8437,N8438,N8439,N8440,N8441,N8442,N8443,N8444,N8447,N8448,N8449,N8450,N8451,N8452,N8453,N8454,N8455,N8456,N8457,N8460,N8463,N8466,N8469,N8470,N8471,N8474,N8477,N8480,N8483,N8484,N8485,N8488,N8489,N8490,N8491,N8492,N8493,N8494,N8495,N8496,N8497,N8500,N8501,N8502,N8503,N8504,N8505,N8506,N8507,N8508,N8509,N8510,N8511,N8512,N8513,N8514,N8515,N8516,N8517,N8518,N8519,N8522,N8525,N8528,N8531,N8534,N8537,N8538,N8539,N8540,N8541,N8545,N8546,N8547,N8548,N8551,N8552,N8553,N8554,N8555,N8558,N8561,N8564,N8565,N8566,N8569,N8572,N8575,N8578,N8579,N8580,N8583,N8586,N8589,N8592,N8595,N8598,N8601,N8604,N8607,N8608,N8609,N8610,N8615,N8616,N8617,N8618,N8619,N8624,N8625,N8626,N8627,N8632,N8633,N8634,N8637,N8638,N8639,N8644,N8645,N8646,N8647,N8648,N8653,N8654,N8655,N8660,N8663,N8666,N8669,N8672,N8675,N8678,N8681,N8684,N8687,N8690,N8693,N8696,N8699,N8702,N8705,N8708,N8711,N8714,N8717,N8718,N8721,N8724,N8727,N8730,N8733,N8734,N8735,N8738,N8741,N8744,N8747,N8750,N8753,N8754,N8755,N8756,N8757,N8760,N8763,N8766,N8769,N8772,N8775,N8778,N8781,N8784,N8787,N8790,N8793,N8796,N8799,N8802,N8805,N8808,N8811,N8814,N8815,N8816,N8817,N8818,N8840,N8857,N8861,N8862,N8863,N8864,N8865,N8866,N8871,N8874,N8878,N8879,N8880,N8881,N8882,N8883,N8884,N8885,N8886,N8887,N8888,N8898,N8902,N8920,N8924,N8927,N8931,N8943,N8950,N8956,N8959,N8960,N8963,N8966,N8991,N8992,N8995,N8996,N9001,N9005,N9024,N9025,N9029,N9035,N9053,N9054,N9064,N9065,N9066,N9067,N9068,N9071,N9072,N9073,N9074,N9077,N9079,N9082,N9083,N9086,N9087,N9088,N9089,N9092,N9093,N9094,N9095,N9098,N9099,N9103,N9107,N9111,N9117,N9127,N9146,N9149,N9159,N9160,N9161,N9165,N9169,N9173,N9179,N9180,N9181,N9182,N9183,N9193,N9203,N9206,N9220,N9223,N9234,N9235,N9236,N9237,N9238,N9242,N9243,N9244,N9245,N9246,N9247,N9248,N9249,N9250,N9251,N9252,N9256,N9257,N9258,N9259,N9260,N9261,N9262,N9265,N9268,N9271,N9272,N9273,N9274,N9275,N9276,N9280,N9285,N9286,N9287,N9288,N9290,N9292,N9294,N9296,N9297,N9298,N9299,N9300,N9301,N9307,N9314,N9315,N9318,N9319,N9320,N9321,N9322,N9323,N9324,N9326,N9332,N9339,N9344,N9352,N9354,N9356,N9358,N9359,N9360,N9361,N9362,N9363,N9364,N9365,N9366,N9367,N9368,N9369,N9370,N9371,N9372,N9375,N9381,N9382,N9383,N9384,N9385,N9392,N9393,N9394,N9395,N9396,N9397,N9398,N9399,N9400,N9401,N9402,N9407,N9408,N9412,N9413,N9414,N9415,N9416,N9417,N9418,N9419,N9420,N9421,N9422,N9423,N9426,N9429,N9432,N9435,N9442,N9445,N9454,N9455,N9456,N9459,N9460,N9461,N9462,N9465,N9466,N9467,N9468,N9473,N9476,N9477,N9478,N9485,N9488,N9493,N9494,N9495,N9498,N9499,N9500,N9505,N9506,N9507,N9508,N9509,N9514,N9515,N9516,N9517,N9520,N9526,N9531,N9539,N9540,N9541,N9543,N9551,N9555,N9556,N9557,N9560,N9561,N9562,N9563,N9564,N9565,N9566,N9567,N9568,N9569,N9570,N9571,N9575,N9579,N9581,N9582,N9585,N9591,N9592,N9593,N9594,N9595,N9596,N9597,N9598,N9599,N9600,N9601,N9602,N9603,N9604,N9605,N9608,N9611,N9612,N9613,N9614,N9615,N9616,N9617,N9618,N9621,N9622,N9623,N9624,N9626,N9629,N9632,N9635,N9642,N9645,N9646,N9649,N9650,N9653,N9656,N9659,N9660,N9661,N9662,N9663,N9666,N9667,N9670,N9671,N9674,N9675,N9678,N9679,N9682,N9685,N9690,N9691,N9692,N9695,N9698,N9702,N9707,N9710,N9711,N9714,N9715,N9716,N9717,N9720,N9721,N9722,N9723,N9726,N9727,N9732,N9733,N9734,N9735,N9736,N9737,N9738,N9739,N9740,N9741,N9742,N9754,N9758,N9762,N9763,N9764,N9765,N9766,N9767,N9768,N9769,N9773,N9774,N9775,N9779,N9784,N9785,N9786,N9790,N9791,N9795,N9796,N9797,N9798,N9799,N9800,N9801,N9802,N9803,N9805,N9806,N9809,N9813,N9814,N9815,N9816,N9817,N9820,N9825,N9826,N9827,N9828,N9829,N9830,N9835,N9836,N9837,N9838,N9846,N9847,N9862,N9863,N9866,N9873,N9876,N9890,N9891,N9892,N9893,N9894,N9895,N9896,N9897,N9898,N9899,N9900,N9901,N9902,N9903,N9904,N9905,N9906,N9907,N9908,N9909,N9910,N9911,N9917,N9923,N9924,N9925,N9932,N9935,N9938,N9939,N9945,N9946,N9947,N9948,N9949,N9953,N9954,N9955,N9956,N9957,N9958,N9959,N9960,N9961,N9964,N9967,N9968,N9969,N9970,N9971,N9972,N9973,N9974,N9975,N9976,N9977,N9978,N9979,N9982,N9983,N9986,N9989,N9992,N9995,N9996,N9997,N9998,N9999,N10002,N10003,N10006,N10007,N10010,N10013,N10014,N10015,N10016,N10017,N10018,N10019,N10020,N10021,N10022,N10023,N10024,N10026,N10028,N10032,N10033,N10034,N10035,N10036,N10037,N10038,N10039,N10040,N10041,N10042,N10043,N10050,N10053,N10054,N10055,N10056,N10057,N10058,N10059,N10060,N10061,N10062,N10067,N10070,N10073,N10076,N10077,N10082,N10083,N10084,N10085,N10086,N10093,N10094,N10105,N10106,N10107,N10108,N10113,N10114,N10115,N10116,N10119,N10124,N10130,N10131,N10132,N10133,N10134,N10135,N10136,N10137,N10138,N10139,N10140,N10141,N10148,N10155,N10156,N10157,N10158,N10159,N10160,N10161,N10162,N10163,N10164,N10165,N10170,N10173,N10176,N10177,N10178,N10179,N10180,N10183,N10186,N10189,N10192,N10195,N10196,N10197,N10200,N10203,N10204,N10205,N10206,N10212,N10213,N10230,N10231,N10232,N10233,N10234,N10237,N10238,N10239,N10240,N10241,N10242,N10247,N10248,N10259,N10264,N10265,N10266,N10267,N10268,N10269,N10270,N10271,N10272,N10273,N10278,N10279,N10280,N10281,N10282,N10283,N10287,N10288,N10289,N10290,N10291,N10292,N10293,N10294,N10295,N10296,N10299,N10300,N10301,N10306,N10307,N10308,N10311,N10314,N10315,N10316,N10317,N10318,N10321,N10324,N10325,N10326,N10327,N10328,N10329,N10330,N10331,N10332,N10333,N10334,N10337,N10338,N10339,N10340,N10341,N10344,N10354,N10357,N10360,N10367,N10375,N10381,N10388,N10391,N10399,N10402,N10406,N10409,N10412,N10415,N10419,N10422,N10425,N10428,N10431,N10432,N10437,N10438,N10439,N10440,N10441,N10444,N10445,N10450,N10451,N10455,N10456,N10465,N10466,N10479,N10497,N10509,N10512,N10515,N10516,N10517,N10518,N10519,N10522,N10525,N10528,N10531,N10534,N10535,N10536,N10539,N10542,N10543,N10544,N10545,N10546,N10547,N10548,N10549,N10550,N10551,N10552,N10553,N10554,N10555,N10556,N10557,N10558,N10559,N10560,N10561,N10562,N10563,N10564,N10565,N10566,N10567,N10568,N10569,N10570,N10571,N10572,N10573,N10577,N10581,N10582,N10583,N10587,N10588,N10589,N10594,N10595,N10596,N10597,N10598,N10602,N10609,N10610,N10621,N10626,N10627,N10629,N10631,N10637,N10638,N10639,N10640,N10642,N10643,N10644,N10645,N10647,N10648,N10649,N10652,N10659,N10662,N10665,N10668,N10671,N10672,N10673,N10674,N10675,N10678,N10681,N10682,N10683,N10684,N10685,N10686,N10687,N10688,N10689,N10690,N10691,N10694,N10695,N10696,N10697,N10698,N10701,N10705,N10707,N10708,N10709,N10710,N10719,N10720,N10730,N10731,N10737,N10738,N10739,N10746,N10747,N10748,N10749,N10750,N10753,N10754,N10764,N10765,N10766,N10767,N10768,N10769,N10770,N10771,N10772,N10773,N10774,N10775,N10776,N10778,N10781,N10784,N10789,N10792,N10796,N10797,N10798,N10799,N10800,N10803,N10806,N10809,N10812,N10815,N10816,N10817,N10820,N10823,N10824,N10825,N10826,N10832,N10833,N10834,N10835,N10836,N10845,N10846,N10857,N10862,N10863,N10864,N10865,N10866,N10867,N10872,N10873,N10874,N10875,N10876,N10879,N10882,N10883,N10884,N10885,N10886,N10887,N10888,N10889,N10890,N10891,N10892,N10895,N10896,N10897,N10898,N10899,N10902,N10909,N10910,N10915,N10916,N10917,N10918,N10919,N10922,N10923,N10928,N10931,N10934,N10935,N10936,N10937,N10938,N10941,N10944,N10947,N10950,N10953,N10954,N10955,N10958,N10961,N10962,N10963,N10964,N10969,N10970,N10981,N10986,N10987,N10988,N10989,N10990,N10991,N10992,N10995,N10998,N10999,N11000,N11001,N11002,N11003,N11004,N11005,N11006,N11007,N11008,N11011,N11012,N11013,N11014,N11015,N11018,N11023,N11024,N11027,N11028,N11029,N11030,N11031,N11034,N11035,N11040,N11041,N11042,N11043,N11044,N11047,N11050,N11053,N11056,N11059,N11062,N11065,N11066,N11067,N11070,N11073,N11074,N11075,N11076,N11077,N11078,N11095,N11098,N11099,N11100,N11103,N11106,N11107,N11108,N11109,N11110,N11111,N11112,N11113,N11114,N11115,N11116,N11117,N11118,N11119,N11120,N11121,N11122,N11123,N11124,N11127,N11130,N11137,N11138,N11139,N11140,N11141,N11142,N11143,N11144,N11145,N11152,N11153,N11154,N11155,N11156,N11159,N11162,N11165,N11168,N11171,N11174,N11177,N11180,N11183,N11184,N11185,N11186,N11187,N11188,N11205,N11210,N11211,N11212,N11213,N11214,N11215,N11216,N11217,N11218,N11219,N11220,N11222,N11223,N11224,N11225,N11226,N11227,N11228,N11229,N11231,N11232,N11233,N11236,N11239,N11242,N11243,N11244,N11245,N11246,N11250,N11252,N11257,N11260,N11261,N11262,N11263,N11264,N11265,N11267,N11268,N11269,N11270,N11272,N11277,N11278,N11279,N11280,N11282,N11283,N11284,N11285,N11286,N11288,N11289,N11290,N11291,N11292,N11293,N11294,N11295,N11296,N11297,N11298,N11299,N11302,N11307,N11308,N11309,N11312,N11313,N11314,N11315,N11316,N11317,N11320,N11321,N11323,N11327,N11328,N11329,N11331,N11335,N11336,N11337,N11338,N11339,N11341;

nb1s1 U1 ( .Q(N387), .DIN(N1) );
nb1s1 U2 ( .Q(N388), .DIN(N1) );
hi1s1 U3 ( .Q(N467), .DIN(N57) );
and2s1 U4 ( .Q(N469), .DIN1(N134), .DIN2(N133) );
nb1s1 U5 ( .Q(N478), .DIN(N248) );
nb1s1 U6 ( .Q(N482), .DIN(N254) );
nb1s1 U7 ( .Q(N484), .DIN(N257) );
nb1s1 U8 ( .Q(N486), .DIN(N260) );
nb1s1 U9 ( .Q(N489), .DIN(N263) );
nb1s1 U10 ( .Q(N492), .DIN(N267) );
and4s1 U11 ( .Q(N494), .DIN1(N162), .DIN2(N172), .DIN3(N188), .DIN4(N199) );
nb1s1 U12 ( .Q(N501), .DIN(N274) );
nb1s1 U13 ( .Q(N505), .DIN(N280) );
nb1s1 U14 ( .Q(N507), .DIN(N283) );
nb1s1 U15 ( .Q(N509), .DIN(N286) );
nb1s1 U16 ( .Q(N511), .DIN(N289) );
nb1s1 U17 ( .Q(N513), .DIN(N293) );
nb1s1 U18 ( .Q(N515), .DIN(N296) );
nb1s1 U19 ( .Q(N517), .DIN(N299) );
nb1s1 U20 ( .Q(N519), .DIN(N303) );
and4s1 U21 ( .Q(N528), .DIN1(N150), .DIN2(N184), .DIN3(N228), .DIN4(N240) );
nb1s1 U22 ( .Q(N535), .DIN(N307) );
nb1s1 U23 ( .Q(N537), .DIN(N310) );
nb1s1 U24 ( .Q(N539), .DIN(N313) );
nb1s1 U25 ( .Q(N541), .DIN(N316) );
nb1s1 U26 ( .Q(N543), .DIN(N319) );
nb1s1 U27 ( .Q(N545), .DIN(N322) );
nb1s1 U28 ( .Q(N547), .DIN(N325) );
nb1s1 U29 ( .Q(N549), .DIN(N328) );
nb1s1 U30 ( .Q(N551), .DIN(N331) );
nb1s1 U31 ( .Q(N553), .DIN(N334) );
nb1s1 U32 ( .Q(N556), .DIN(N337) );
nb1s1 U33 ( .Q(N559), .DIN(N343) );
nb1s1 U34 ( .Q(N561), .DIN(N346) );
nb1s1 U35 ( .Q(N563), .DIN(N349) );
nb1s1 U36 ( .Q(N565), .DIN(N352) );
nb1s1 U37 ( .Q(N567), .DIN(N355) );
nb1s1 U38 ( .Q(N569), .DIN(N358) );
nb1s1 U39 ( .Q(N571), .DIN(N361) );
nb1s1 U40 ( .Q(N573), .DIN(N364) );
and4s1 U41 ( .Q(N575), .DIN1(N183), .DIN2(N182), .DIN3(N185), .DIN4(N186) );
and4s1 U42 ( .Q(N578), .DIN1(N210), .DIN2(N152), .DIN3(N218), .DIN4(N230) );
hi1s1 U43 ( .Q(N582), .DIN(N15) );
hi1s1 U44 ( .Q(N585), .DIN(N5) );
nb1s1 U45 ( .Q(N590), .DIN(N1) );
hi1s1 U46 ( .Q(N593), .DIN(N5) );
hi1s1 U47 ( .Q(N596), .DIN(N5) );
hi1s1 U48 ( .Q(N599), .DIN(N289) );
hi1s1 U49 ( .Q(N604), .DIN(N299) );
hi1s1 U50 ( .Q(N609), .DIN(N303) );
nb1s1 U51 ( .Q(N614), .DIN(N38) );
nb1s1 U52 ( .Q(N625), .DIN(N15) );
nnd2s1 U53 ( .Q(N628), .DIN1(N12), .DIN2(N9) );
nnd2s1 U54 ( .Q(N632), .DIN1(N12), .DIN2(N9) );
nb1s1 U55 ( .Q(N636), .DIN(N38) );
hi1s1 U56 ( .Q(N641), .DIN(N245) );
hi1s1 U57 ( .Q(N642), .DIN(N248) );
nb1s1 U58 ( .Q(N643), .DIN(N251) );
hi1s1 U59 ( .Q(N644), .DIN(N251) );
hi1s1 U60 ( .Q(N651), .DIN(N254) );
nb1s1 U61 ( .Q(N657), .DIN(N106) );
hi1s1 U62 ( .Q(N660), .DIN(N257) );
hi1s1 U63 ( .Q(N666), .DIN(N260) );
hi1s1 U64 ( .Q(N672), .DIN(N263) );
hi1s1 U65 ( .Q(N673), .DIN(N267) );
hi1s1 U66 ( .Q(N674), .DIN(N106) );
nb1s1 U67 ( .Q(N676), .DIN(N18) );
nb1s1 U68 ( .Q(N682), .DIN(N18) );
and2s1 U69 ( .Q(N688), .DIN1(N382), .DIN2(N263) );
nb1s1 U70 ( .Q(N689), .DIN(N18) );
hi1s1 U71 ( .Q(N695), .DIN(N18) );
nnd2s1 U72 ( .Q(N700), .DIN1(N382), .DIN2(N267) );
hi1s1 U73 ( .Q(N705), .DIN(N271) );
hi1s1 U74 ( .Q(N706), .DIN(N274) );
nb1s1 U75 ( .Q(N707), .DIN(N277) );
hi1s1 U76 ( .Q(N708), .DIN(N277) );
hi1s1 U77 ( .Q(N715), .DIN(N280) );
hi1s1 U78 ( .Q(N721), .DIN(N283) );
hi1s1 U79 ( .Q(N727), .DIN(N286) );
hi1s1 U80 ( .Q(N733), .DIN(N289) );
hi1s1 U81 ( .Q(N734), .DIN(N293) );
hi1s1 U82 ( .Q(N742), .DIN(N296) );
hi1s1 U83 ( .Q(N748), .DIN(N299) );
hi1s1 U84 ( .Q(N749), .DIN(N303) );
nb1s1 U85 ( .Q(N750), .DIN(N367) );
hi1s1 U86 ( .Q(N758), .DIN(N307) );
hi1s1 U87 ( .Q(N759), .DIN(N310) );
hi1s1 U88 ( .Q(N762), .DIN(N313) );
hi1s1 U89 ( .Q(N768), .DIN(N316) );
hi1s1 U90 ( .Q(N774), .DIN(N319) );
hi1s1 U91 ( .Q(N780), .DIN(N322) );
hi1s1 U92 ( .Q(N786), .DIN(N325) );
hi1s1 U93 ( .Q(N794), .DIN(N328) );
hi1s1 U94 ( .Q(N800), .DIN(N331) );
hi1s1 U95 ( .Q(N806), .DIN(N334) );
hi1s1 U96 ( .Q(N812), .DIN(N337) );
nb1s1 U97 ( .Q(N813), .DIN(N340) );
hi1s1 U98 ( .Q(N814), .DIN(N340) );
hi1s1 U99 ( .Q(N821), .DIN(N343) );
hi1s1 U100 ( .Q(N827), .DIN(N346) );
hi1s1 U101 ( .Q(N833), .DIN(N349) );
hi1s1 U102 ( .Q(N839), .DIN(N352) );
hi1s1 U103 ( .Q(N845), .DIN(N355) );
hi1s1 U104 ( .Q(N853), .DIN(N358) );
hi1s1 U105 ( .Q(N859), .DIN(N361) );
hi1s1 U106 ( .Q(N865), .DIN(N364) );
nb1s1 U107 ( .Q(N871), .DIN(N367) );
nnd2s1 U108 ( .Q(N881), .DIN1(N467), .DIN2(N585) );
hi1s1 U109 ( .Q(N882), .DIN(N528) );
hi1s1 U110 ( .Q(N883), .DIN(N578) );
hi1s1 U111 ( .Q(N884), .DIN(N575) );
hi1s1 U112 ( .Q(N885), .DIN(N494) );
and2s1 U113 ( .Q(N886), .DIN1(N528), .DIN2(N578) );
and2s1 U114 ( .Q(N887), .DIN1(N575), .DIN2(N494) );
nb1s1 U115 ( .Q(N889), .DIN(N590) );
nb1s1 U116 ( .Q(N945), .DIN(N657) );
hi1s1 U117 ( .Q(N957), .DIN(N688) );
and2s1 U118 ( .Q(N1028), .DIN1(N382), .DIN2(N641) );
nnd2s1 U119 ( .Q(N1029), .DIN1(N382), .DIN2(N705) );
and2s1 U120 ( .Q(N1109), .DIN1(N469), .DIN2(N596) );
nnd2s1 U121 ( .Q(N1110), .DIN1(N242), .DIN2(N593) );
hi1s1 U122 ( .Q(N1111), .DIN(N625) );
nnd2s1 U123 ( .Q(N1112), .DIN1(N242), .DIN2(N593) );
nnd2s1 U124 ( .Q(N1113), .DIN1(N469), .DIN2(N596) );
hi1s1 U125 ( .Q(N1114), .DIN(N625) );
hi1s1 U126 ( .Q(N1115), .DIN(N871) );
nb1s1 U127 ( .Q(N1116), .DIN(N590) );
nb1s1 U128 ( .Q(N1119), .DIN(N628) );
nb1s1 U129 ( .Q(N1125), .DIN(N682) );
nb1s1 U130 ( .Q(N1132), .DIN(N628) );
nb1s1 U131 ( .Q(N1136), .DIN(N682) );
nb1s1 U132 ( .Q(N1141), .DIN(N628) );
nb1s1 U133 ( .Q(N1147), .DIN(N682) );
nb1s1 U134 ( .Q(N1154), .DIN(N632) );
nb1s1 U135 ( .Q(N1160), .DIN(N676) );
and2s1 U136 ( .Q(N1167), .DIN1(N700), .DIN2(N614) );
and2s1 U137 ( .Q(N1174), .DIN1(N700), .DIN2(N614) );
nb1s1 U138 ( .Q(N1175), .DIN(N682) );
nb1s1 U139 ( .Q(N1182), .DIN(N676) );
hi1s1 U140 ( .Q(N1189), .DIN(N657) );
hi1s1 U141 ( .Q(N1194), .DIN(N676) );
hi1s1 U142 ( .Q(N1199), .DIN(N682) );
hi1s1 U143 ( .Q(N1206), .DIN(N689) );
nb1s1 U144 ( .Q(N1211), .DIN(N695) );
hi1s1 U145 ( .Q(N1218), .DIN(N750) );
hi1s1 U146 ( .Q(N1222), .DIN(N1028) );
nb1s1 U147 ( .Q(N1227), .DIN(N632) );
nb1s1 U148 ( .Q(N1233), .DIN(N676) );
nb1s1 U149 ( .Q(N1240), .DIN(N632) );
nb1s1 U150 ( .Q(N1244), .DIN(N676) );
nb1s1 U151 ( .Q(N1249), .DIN(N689) );
nb1s1 U152 ( .Q(N1256), .DIN(N689) );
nb1s1 U153 ( .Q(N1263), .DIN(N695) );
nb1s1 U154 ( .Q(N1270), .DIN(N689) );
nb1s1 U155 ( .Q(N1277), .DIN(N689) );
nb1s1 U156 ( .Q(N1284), .DIN(N700) );
nb1s1 U157 ( .Q(N1287), .DIN(N614) );
nb1s1 U158 ( .Q(N1290), .DIN(N666) );
nb1s1 U159 ( .Q(N1293), .DIN(N660) );
nb1s1 U160 ( .Q(N1296), .DIN(N651) );
nb1s1 U161 ( .Q(N1299), .DIN(N614) );
nb1s1 U162 ( .Q(N1302), .DIN(N644) );
nb1s1 U163 ( .Q(N1305), .DIN(N700) );
nb1s1 U164 ( .Q(N1308), .DIN(N614) );
nb1s1 U165 ( .Q(N1311), .DIN(N614) );
nb1s1 U166 ( .Q(N1314), .DIN(N666) );
nb1s1 U167 ( .Q(N1317), .DIN(N660) );
nb1s1 U168 ( .Q(N1320), .DIN(N651) );
nb1s1 U169 ( .Q(N1323), .DIN(N644) );
nb1s1 U170 ( .Q(N1326), .DIN(N609) );
nb1s1 U171 ( .Q(N1329), .DIN(N604) );
nb1s1 U172 ( .Q(N1332), .DIN(N742) );
nb1s1 U173 ( .Q(N1335), .DIN(N599) );
nb1s1 U174 ( .Q(N1338), .DIN(N727) );
nb1s1 U175 ( .Q(N1341), .DIN(N721) );
nb1s1 U176 ( .Q(N1344), .DIN(N715) );
nb1s1 U177 ( .Q(N1347), .DIN(N734) );
nb1s1 U178 ( .Q(N1350), .DIN(N708) );
nb1s1 U179 ( .Q(N1353), .DIN(N609) );
nb1s1 U180 ( .Q(N1356), .DIN(N604) );
nb1s1 U181 ( .Q(N1359), .DIN(N742) );
nb1s1 U182 ( .Q(N1362), .DIN(N734) );
nb1s1 U183 ( .Q(N1365), .DIN(N599) );
nb1s1 U184 ( .Q(N1368), .DIN(N727) );
nb1s1 U185 ( .Q(N1371), .DIN(N721) );
nb1s1 U186 ( .Q(N1374), .DIN(N715) );
nb1s1 U187 ( .Q(N1377), .DIN(N708) );
nb1s1 U188 ( .Q(N1380), .DIN(N806) );
nb1s1 U189 ( .Q(N1383), .DIN(N800) );
nb1s1 U190 ( .Q(N1386), .DIN(N794) );
nb1s1 U191 ( .Q(N1389), .DIN(N786) );
nb1s1 U192 ( .Q(N1392), .DIN(N780) );
nb1s1 U193 ( .Q(N1395), .DIN(N774) );
nb1s1 U194 ( .Q(N1398), .DIN(N768) );
nb1s1 U195 ( .Q(N1401), .DIN(N762) );
nb1s1 U196 ( .Q(N1404), .DIN(N806) );
nb1s1 U197 ( .Q(N1407), .DIN(N800) );
nb1s1 U198 ( .Q(N1410), .DIN(N794) );
nb1s1 U199 ( .Q(N1413), .DIN(N780) );
nb1s1 U200 ( .Q(N1416), .DIN(N774) );
nb1s1 U201 ( .Q(N1419), .DIN(N768) );
nb1s1 U202 ( .Q(N1422), .DIN(N762) );
nb1s1 U203 ( .Q(N1425), .DIN(N786) );
nb1s1 U204 ( .Q(N1428), .DIN(N636) );
nb1s1 U205 ( .Q(N1431), .DIN(N636) );
nb1s1 U206 ( .Q(N1434), .DIN(N865) );
nb1s1 U207 ( .Q(N1437), .DIN(N859) );
nb1s1 U208 ( .Q(N1440), .DIN(N853) );
nb1s1 U209 ( .Q(N1443), .DIN(N845) );
nb1s1 U210 ( .Q(N1446), .DIN(N839) );
nb1s1 U211 ( .Q(N1449), .DIN(N833) );
nb1s1 U212 ( .Q(N1452), .DIN(N827) );
nb1s1 U213 ( .Q(N1455), .DIN(N821) );
nb1s1 U214 ( .Q(N1458), .DIN(N814) );
nb1s1 U215 ( .Q(N1461), .DIN(N865) );
nb1s1 U216 ( .Q(N1464), .DIN(N859) );
nb1s1 U217 ( .Q(N1467), .DIN(N853) );
nb1s1 U218 ( .Q(N1470), .DIN(N839) );
nb1s1 U219 ( .Q(N1473), .DIN(N833) );
nb1s1 U220 ( .Q(N1476), .DIN(N827) );
nb1s1 U221 ( .Q(N1479), .DIN(N821) );
nb1s1 U222 ( .Q(N1482), .DIN(N845) );
nb1s1 U223 ( .Q(N1485), .DIN(N814) );
hi1s1 U224 ( .Q(N1489), .DIN(N1109) );
nb1s1 U225 ( .Q(N1490), .DIN(N1116) );
and2s1 U226 ( .Q(N1537), .DIN1(N957), .DIN2(N614) );
and2s1 U227 ( .Q(N1551), .DIN1(N614), .DIN2(N957) );
and2s1 U228 ( .Q(N1649), .DIN1(N1029), .DIN2(N636) );
nb1s1 U229 ( .Q(N1703), .DIN(N957) );
nor2s1 U230 ( .Q(N1708), .DIN1(N957), .DIN2(N614) );
nb1s1 U231 ( .Q(N1713), .DIN(N957) );
nor2s1 U232 ( .Q(N1721), .DIN1(N614), .DIN2(N957) );
nb1s1 U233 ( .Q(N1758), .DIN(N1029) );
and2s1 U234 ( .Q(N1781), .DIN1(N163), .DIN2(N1116) );
and2s1 U235 ( .Q(N1782), .DIN1(N170), .DIN2(N1125) );
hi1s1 U236 ( .Q(N1783), .DIN(N1125) );
hi1s1 U237 ( .Q(N1789), .DIN(N1136) );
and2s1 U238 ( .Q(N1793), .DIN1(N169), .DIN2(N1125) );
and2s1 U239 ( .Q(N1794), .DIN1(N168), .DIN2(N1125) );
and2s1 U240 ( .Q(N1795), .DIN1(N167), .DIN2(N1125) );
and2s1 U241 ( .Q(N1796), .DIN1(N166), .DIN2(N1136) );
and2s1 U242 ( .Q(N1797), .DIN1(N165), .DIN2(N1136) );
and2s1 U243 ( .Q(N1798), .DIN1(N164), .DIN2(N1136) );
hi1s1 U244 ( .Q(N1799), .DIN(N1147) );
hi1s1 U245 ( .Q(N1805), .DIN(N1160) );
and2s1 U246 ( .Q(N1811), .DIN1(N177), .DIN2(N1147) );
and2s1 U247 ( .Q(N1812), .DIN1(N176), .DIN2(N1147) );
and2s1 U248 ( .Q(N1813), .DIN1(N175), .DIN2(N1147) );
and2s1 U249 ( .Q(N1814), .DIN1(N174), .DIN2(N1147) );
and2s1 U250 ( .Q(N1815), .DIN1(N173), .DIN2(N1147) );
and2s1 U251 ( .Q(N1816), .DIN1(N157), .DIN2(N1160) );
and2s1 U252 ( .Q(N1817), .DIN1(N156), .DIN2(N1160) );
and2s1 U253 ( .Q(N1818), .DIN1(N155), .DIN2(N1160) );
and2s1 U254 ( .Q(N1819), .DIN1(N154), .DIN2(N1160) );
and2s1 U255 ( .Q(N1820), .DIN1(N153), .DIN2(N1160) );
hi1s1 U256 ( .Q(N1821), .DIN(N1284) );
hi1s1 U257 ( .Q(N1822), .DIN(N1287) );
hi1s1 U258 ( .Q(N1828), .DIN(N1290) );
hi1s1 U259 ( .Q(N1829), .DIN(N1293) );
hi1s1 U260 ( .Q(N1830), .DIN(N1296) );
hi1s1 U261 ( .Q(N1832), .DIN(N1299) );
hi1s1 U262 ( .Q(N1833), .DIN(N1302) );
hi1s1 U263 ( .Q(N1834), .DIN(N1305) );
hi1s1 U264 ( .Q(N1835), .DIN(N1308) );
hi1s1 U265 ( .Q(N1839), .DIN(N1311) );
hi1s1 U266 ( .Q(N1840), .DIN(N1314) );
hi1s1 U267 ( .Q(N1841), .DIN(N1317) );
hi1s1 U268 ( .Q(N1842), .DIN(N1320) );
hi1s1 U269 ( .Q(N1843), .DIN(N1323) );
hi1s1 U270 ( .Q(N1845), .DIN(N1175) );
hi1s1 U271 ( .Q(N1851), .DIN(N1182) );
and2s1 U272 ( .Q(N1857), .DIN1(N181), .DIN2(N1175) );
and2s1 U273 ( .Q(N1858), .DIN1(N171), .DIN2(N1175) );
and2s1 U274 ( .Q(N1859), .DIN1(N180), .DIN2(N1175) );
and2s1 U275 ( .Q(N1860), .DIN1(N179), .DIN2(N1175) );
and2s1 U276 ( .Q(N1861), .DIN1(N178), .DIN2(N1175) );
and2s1 U277 ( .Q(N1862), .DIN1(N161), .DIN2(N1182) );
and2s1 U278 ( .Q(N1863), .DIN1(N151), .DIN2(N1182) );
and2s1 U279 ( .Q(N1864), .DIN1(N160), .DIN2(N1182) );
and2s1 U280 ( .Q(N1865), .DIN1(N159), .DIN2(N1182) );
and2s1 U281 ( .Q(N1866), .DIN1(N158), .DIN2(N1182) );
hi1s1 U282 ( .Q(N1867), .DIN(N1326) );
hi1s1 U283 ( .Q(N1868), .DIN(N1329) );
hi1s1 U284 ( .Q(N1869), .DIN(N1332) );
hi1s1 U285 ( .Q(N1870), .DIN(N1335) );
hi1s1 U286 ( .Q(N1871), .DIN(N1338) );
hi1s1 U287 ( .Q(N1872), .DIN(N1341) );
hi1s1 U288 ( .Q(N1873), .DIN(N1344) );
hi1s1 U289 ( .Q(N1874), .DIN(N1347) );
hi1s1 U290 ( .Q(N1875), .DIN(N1350) );
hi1s1 U291 ( .Q(N1876), .DIN(N1353) );
hi1s1 U292 ( .Q(N1877), .DIN(N1356) );
hi1s1 U293 ( .Q(N1878), .DIN(N1359) );
hi1s1 U294 ( .Q(N1879), .DIN(N1362) );
hi1s1 U295 ( .Q(N1880), .DIN(N1365) );
hi1s1 U296 ( .Q(N1881), .DIN(N1368) );
hi1s1 U297 ( .Q(N1882), .DIN(N1371) );
hi1s1 U298 ( .Q(N1883), .DIN(N1374) );
hi1s1 U299 ( .Q(N1884), .DIN(N1377) );
nb1s1 U300 ( .Q(N1885), .DIN(N1199) );
nb1s1 U301 ( .Q(N1892), .DIN(N1194) );
nb1s1 U302 ( .Q(N1899), .DIN(N1199) );
nb1s1 U303 ( .Q(N1906), .DIN(N1194) );
hi1s1 U304 ( .Q(N1913), .DIN(N1211) );
nb1s1 U305 ( .Q(N1919), .DIN(N1194) );
and2s1 U306 ( .Q(N1926), .DIN1(N44), .DIN2(N1211) );
and2s1 U307 ( .Q(N1927), .DIN1(N41), .DIN2(N1211) );
and2s1 U308 ( .Q(N1928), .DIN1(N29), .DIN2(N1211) );
and2s1 U309 ( .Q(N1929), .DIN1(N26), .DIN2(N1211) );
and2s1 U310 ( .Q(N1930), .DIN1(N23), .DIN2(N1211) );
hi1s1 U311 ( .Q(N1931), .DIN(N1380) );
hi1s1 U312 ( .Q(N1932), .DIN(N1383) );
hi1s1 U313 ( .Q(N1933), .DIN(N1386) );
hi1s1 U314 ( .Q(N1934), .DIN(N1389) );
hi1s1 U315 ( .Q(N1935), .DIN(N1392) );
hi1s1 U316 ( .Q(N1936), .DIN(N1395) );
hi1s1 U317 ( .Q(N1937), .DIN(N1398) );
hi1s1 U318 ( .Q(N1938), .DIN(N1401) );
hi1s1 U319 ( .Q(N1939), .DIN(N1404) );
hi1s1 U320 ( .Q(N1940), .DIN(N1407) );
hi1s1 U321 ( .Q(N1941), .DIN(N1410) );
hi1s1 U322 ( .Q(N1942), .DIN(N1413) );
hi1s1 U323 ( .Q(N1943), .DIN(N1416) );
hi1s1 U324 ( .Q(N1944), .DIN(N1419) );
hi1s1 U325 ( .Q(N1945), .DIN(N1422) );
hi1s1 U326 ( .Q(N1946), .DIN(N1425) );
hi1s1 U327 ( .Q(N1947), .DIN(N1233) );
hi1s1 U328 ( .Q(N1953), .DIN(N1244) );
and2s1 U329 ( .Q(N1957), .DIN1(N209), .DIN2(N1233) );
and2s1 U330 ( .Q(N1958), .DIN1(N216), .DIN2(N1233) );
and2s1 U331 ( .Q(N1959), .DIN1(N215), .DIN2(N1233) );
and2s1 U332 ( .Q(N1960), .DIN1(N214), .DIN2(N1233) );
and2s1 U333 ( .Q(N1961), .DIN1(N213), .DIN2(N1244) );
and2s1 U334 ( .Q(N1962), .DIN1(N212), .DIN2(N1244) );
and2s1 U335 ( .Q(N1963), .DIN1(N211), .DIN2(N1244) );
hi1s1 U336 ( .Q(N1965), .DIN(N1428) );
and2s1 U337 ( .Q(N1966), .DIN1(N1222), .DIN2(N636) );
hi1s1 U338 ( .Q(N1967), .DIN(N1431) );
hi1s1 U339 ( .Q(N1968), .DIN(N1434) );
hi1s1 U340 ( .Q(N1969), .DIN(N1437) );
hi1s1 U341 ( .Q(N1970), .DIN(N1440) );
hi1s1 U342 ( .Q(N1971), .DIN(N1443) );
hi1s1 U343 ( .Q(N1972), .DIN(N1446) );
hi1s1 U344 ( .Q(N1973), .DIN(N1449) );
hi1s1 U345 ( .Q(N1974), .DIN(N1452) );
hi1s1 U346 ( .Q(N1975), .DIN(N1455) );
hi1s1 U347 ( .Q(N1976), .DIN(N1458) );
hi1s1 U348 ( .Q(N1977), .DIN(N1249) );
hi1s1 U349 ( .Q(N1983), .DIN(N1256) );
and2s1 U350 ( .Q(N1989), .DIN1(N642), .DIN2(N1249) );
and2s1 U351 ( .Q(N1990), .DIN1(N644), .DIN2(N1249) );
and2s1 U352 ( .Q(N1991), .DIN1(N651), .DIN2(N1249) );
and2s1 U353 ( .Q(N1992), .DIN1(N674), .DIN2(N1249) );
and2s1 U354 ( .Q(N1993), .DIN1(N660), .DIN2(N1249) );
and2s1 U355 ( .Q(N1994), .DIN1(N666), .DIN2(N1256) );
and2s1 U356 ( .Q(N1995), .DIN1(N672), .DIN2(N1256) );
and2s1 U357 ( .Q(N1996), .DIN1(N673), .DIN2(N1256) );
hi1s1 U358 ( .Q(N1997), .DIN(N1263) );
nb1s1 U359 ( .Q(N2003), .DIN(N1194) );
and2s1 U360 ( .Q(N2010), .DIN1(N47), .DIN2(N1263) );
and2s1 U361 ( .Q(N2011), .DIN1(N35), .DIN2(N1263) );
and2s1 U362 ( .Q(N2012), .DIN1(N32), .DIN2(N1263) );
and2s1 U363 ( .Q(N2013), .DIN1(N50), .DIN2(N1263) );
and2s1 U364 ( .Q(N2014), .DIN1(N66), .DIN2(N1263) );
hi1s1 U365 ( .Q(N2015), .DIN(N1461) );
hi1s1 U366 ( .Q(N2016), .DIN(N1464) );
hi1s1 U367 ( .Q(N2017), .DIN(N1467) );
hi1s1 U368 ( .Q(N2018), .DIN(N1470) );
hi1s1 U369 ( .Q(N2019), .DIN(N1473) );
hi1s1 U370 ( .Q(N2020), .DIN(N1476) );
hi1s1 U371 ( .Q(N2021), .DIN(N1479) );
hi1s1 U372 ( .Q(N2022), .DIN(N1482) );
hi1s1 U373 ( .Q(N2023), .DIN(N1485) );
nb1s1 U374 ( .Q(N2024), .DIN(N1206) );
nb1s1 U375 ( .Q(N2031), .DIN(N1206) );
nb1s1 U376 ( .Q(N2038), .DIN(N1206) );
nb1s1 U377 ( .Q(N2045), .DIN(N1206) );
hi1s1 U378 ( .Q(N2052), .DIN(N1270) );
hi1s1 U379 ( .Q(N2058), .DIN(N1277) );
and2s1 U380 ( .Q(N2064), .DIN1(N706), .DIN2(N1270) );
and2s1 U381 ( .Q(N2065), .DIN1(N708), .DIN2(N1270) );
and2s1 U382 ( .Q(N2066), .DIN1(N715), .DIN2(N1270) );
and2s1 U383 ( .Q(N2067), .DIN1(N721), .DIN2(N1270) );
and2s1 U384 ( .Q(N2068), .DIN1(N727), .DIN2(N1270) );
and2s1 U385 ( .Q(N2069), .DIN1(N733), .DIN2(N1277) );
and2s1 U386 ( .Q(N2070), .DIN1(N734), .DIN2(N1277) );
and2s1 U387 ( .Q(N2071), .DIN1(N742), .DIN2(N1277) );
and2s1 U388 ( .Q(N2072), .DIN1(N748), .DIN2(N1277) );
and2s1 U389 ( .Q(N2073), .DIN1(N749), .DIN2(N1277) );
nb1s1 U390 ( .Q(N2074), .DIN(N1189) );
nb1s1 U391 ( .Q(N2081), .DIN(N1189) );
nb1s1 U392 ( .Q(N2086), .DIN(N1222) );
nnd2s1 U393 ( .Q(N2107), .DIN1(N1287), .DIN2(N1821) );
nnd2s1 U394 ( .Q(N2108), .DIN1(N1284), .DIN2(N1822) );
hi1s1 U395 ( .Q(N2110), .DIN(N1703) );
nnd2s1 U396 ( .Q(N2111), .DIN1(N1703), .DIN2(N1832) );
nnd2s1 U397 ( .Q(N2112), .DIN1(N1308), .DIN2(N1834) );
nnd2s1 U398 ( .Q(N2113), .DIN1(N1305), .DIN2(N1835) );
hi1s1 U399 ( .Q(N2114), .DIN(N1713) );
nnd2s1 U400 ( .Q(N2115), .DIN1(N1713), .DIN2(N1839) );
hi1s1 U401 ( .Q(N2117), .DIN(N1721) );
hi1s1 U402 ( .Q(N2171), .DIN(N1758) );
nnd2s1 U403 ( .Q(N2172), .DIN1(N1758), .DIN2(N1965) );
hi1s1 U404 ( .Q(N2230), .DIN(N1708) );
nb1s1 U405 ( .Q(N2231), .DIN(N1537) );
nb1s1 U406 ( .Q(N2235), .DIN(N1551) );
or2s1 U407 ( .Q(N2239), .DIN1(N1783), .DIN2(N1782) );
or2s1 U408 ( .Q(N2240), .DIN1(N1783), .DIN2(N1125) );
or2s1 U409 ( .Q(N2241), .DIN1(N1783), .DIN2(N1793) );
or2s1 U410 ( .Q(N2242), .DIN1(N1783), .DIN2(N1794) );
or2s1 U411 ( .Q(N2243), .DIN1(N1783), .DIN2(N1795) );
or2s1 U412 ( .Q(N2244), .DIN1(N1789), .DIN2(N1796) );
or2s1 U413 ( .Q(N2245), .DIN1(N1789), .DIN2(N1797) );
or2s1 U414 ( .Q(N2246), .DIN1(N1789), .DIN2(N1798) );
or2s1 U415 ( .Q(N2247), .DIN1(N1799), .DIN2(N1811) );
or2s1 U416 ( .Q(N2248), .DIN1(N1799), .DIN2(N1812) );
or2s1 U417 ( .Q(N2249), .DIN1(N1799), .DIN2(N1813) );
or2s1 U418 ( .Q(N2250), .DIN1(N1799), .DIN2(N1814) );
or2s1 U419 ( .Q(N2251), .DIN1(N1799), .DIN2(N1815) );
or2s1 U420 ( .Q(N2252), .DIN1(N1805), .DIN2(N1816) );
or2s1 U421 ( .Q(N2253), .DIN1(N1805), .DIN2(N1817) );
or2s1 U422 ( .Q(N2254), .DIN1(N1805), .DIN2(N1818) );
or2s1 U423 ( .Q(N2255), .DIN1(N1805), .DIN2(N1819) );
or2s1 U424 ( .Q(N2256), .DIN1(N1805), .DIN2(N1820) );
nnd2s1 U425 ( .Q(N2257), .DIN1(N2107), .DIN2(N2108) );
hi1s1 U426 ( .Q(N2267), .DIN(N2074) );
nnd2s1 U427 ( .Q(N2268), .DIN1(N1299), .DIN2(N2110) );
nnd2s1 U428 ( .Q(N2269), .DIN1(N2112), .DIN2(N2113) );
nnd2s1 U429 ( .Q(N2274), .DIN1(N1311), .DIN2(N2114) );
hi1s1 U430 ( .Q(N2275), .DIN(N2081) );
and2s1 U431 ( .Q(N2277), .DIN1(N141), .DIN2(N1845) );
and2s1 U432 ( .Q(N2278), .DIN1(N147), .DIN2(N1845) );
and2s1 U433 ( .Q(N2279), .DIN1(N138), .DIN2(N1845) );
and2s1 U434 ( .Q(N2280), .DIN1(N144), .DIN2(N1845) );
and2s1 U435 ( .Q(N2281), .DIN1(N135), .DIN2(N1845) );
and2s1 U436 ( .Q(N2282), .DIN1(N141), .DIN2(N1851) );
and2s1 U437 ( .Q(N2283), .DIN1(N147), .DIN2(N1851) );
and2s1 U438 ( .Q(N2284), .DIN1(N138), .DIN2(N1851) );
and2s1 U439 ( .Q(N2285), .DIN1(N144), .DIN2(N1851) );
and2s1 U440 ( .Q(N2286), .DIN1(N135), .DIN2(N1851) );
hi1s1 U441 ( .Q(N2287), .DIN(N1885) );
hi1s1 U442 ( .Q(N2293), .DIN(N1892) );
and2s1 U443 ( .Q(N2299), .DIN1(N103), .DIN2(N1885) );
and2s1 U444 ( .Q(N2300), .DIN1(N130), .DIN2(N1885) );
and2s1 U445 ( .Q(N2301), .DIN1(N127), .DIN2(N1885) );
and2s1 U446 ( .Q(N2302), .DIN1(N124), .DIN2(N1885) );
and2s1 U447 ( .Q(N2303), .DIN1(N100), .DIN2(N1885) );
and2s1 U448 ( .Q(N2304), .DIN1(N103), .DIN2(N1892) );
and2s1 U449 ( .Q(N2305), .DIN1(N130), .DIN2(N1892) );
and2s1 U450 ( .Q(N2306), .DIN1(N127), .DIN2(N1892) );
and2s1 U451 ( .Q(N2307), .DIN1(N124), .DIN2(N1892) );
and2s1 U452 ( .Q(N2308), .DIN1(N100), .DIN2(N1892) );
hi1s1 U453 ( .Q(N2309), .DIN(N1899) );
hi1s1 U454 ( .Q(N2315), .DIN(N1906) );
and2s1 U455 ( .Q(N2321), .DIN1(N115), .DIN2(N1899) );
and2s1 U456 ( .Q(N2322), .DIN1(N118), .DIN2(N1899) );
and2s1 U457 ( .Q(N2323), .DIN1(N97), .DIN2(N1899) );
and2s1 U458 ( .Q(N2324), .DIN1(N94), .DIN2(N1899) );
and2s1 U459 ( .Q(N2325), .DIN1(N121), .DIN2(N1899) );
and2s1 U460 ( .Q(N2326), .DIN1(N115), .DIN2(N1906) );
and2s1 U461 ( .Q(N2327), .DIN1(N118), .DIN2(N1906) );
and2s1 U462 ( .Q(N2328), .DIN1(N97), .DIN2(N1906) );
and2s1 U463 ( .Q(N2329), .DIN1(N94), .DIN2(N1906) );
and2s1 U464 ( .Q(N2330), .DIN1(N121), .DIN2(N1906) );
hi1s1 U465 ( .Q(N2331), .DIN(N1919) );
and2s1 U466 ( .Q(N2337), .DIN1(N208), .DIN2(N1913) );
and2s1 U467 ( .Q(N2338), .DIN1(N198), .DIN2(N1913) );
and2s1 U468 ( .Q(N2339), .DIN1(N207), .DIN2(N1913) );
and2s1 U469 ( .Q(N2340), .DIN1(N206), .DIN2(N1913) );
and2s1 U470 ( .Q(N2341), .DIN1(N205), .DIN2(N1913) );
and2s1 U471 ( .Q(N2342), .DIN1(N44), .DIN2(N1919) );
and2s1 U472 ( .Q(N2343), .DIN1(N41), .DIN2(N1919) );
and2s1 U473 ( .Q(N2344), .DIN1(N29), .DIN2(N1919) );
and2s1 U474 ( .Q(N2345), .DIN1(N26), .DIN2(N1919) );
and2s1 U475 ( .Q(N2346), .DIN1(N23), .DIN2(N1919) );
or2s1 U476 ( .Q(N2347), .DIN1(N1947), .DIN2(N1233) );
or2s1 U477 ( .Q(N2348), .DIN1(N1947), .DIN2(N1957) );
or2s1 U478 ( .Q(N2349), .DIN1(N1947), .DIN2(N1958) );
or2s1 U479 ( .Q(N2350), .DIN1(N1947), .DIN2(N1959) );
or2s1 U480 ( .Q(N2351), .DIN1(N1947), .DIN2(N1960) );
or2s1 U481 ( .Q(N2352), .DIN1(N1953), .DIN2(N1961) );
or2s1 U482 ( .Q(N2353), .DIN1(N1953), .DIN2(N1962) );
or2s1 U483 ( .Q(N2354), .DIN1(N1953), .DIN2(N1963) );
nnd2s1 U484 ( .Q(N2355), .DIN1(N1428), .DIN2(N2171) );
hi1s1 U485 ( .Q(N2356), .DIN(N2086) );
nnd2s1 U486 ( .Q(N2357), .DIN1(N2086), .DIN2(N1967) );
and2s1 U487 ( .Q(N2358), .DIN1(N114), .DIN2(N1977) );
and2s1 U488 ( .Q(N2359), .DIN1(N113), .DIN2(N1977) );
and2s1 U489 ( .Q(N2360), .DIN1(N111), .DIN2(N1977) );
and2s1 U490 ( .Q(N2361), .DIN1(N87), .DIN2(N1977) );
and2s1 U491 ( .Q(N2362), .DIN1(N112), .DIN2(N1977) );
and2s1 U492 ( .Q(N2363), .DIN1(N88), .DIN2(N1983) );
and2s1 U493 ( .Q(N2364), .DIN1(N245), .DIN2(N1983) );
and2s1 U494 ( .Q(N2365), .DIN1(N271), .DIN2(N1983) );
and2s1 U495 ( .Q(N2366), .DIN1(N759), .DIN2(N1983) );
and2s1 U496 ( .Q(N2367), .DIN1(N70), .DIN2(N1983) );
hi1s1 U497 ( .Q(N2368), .DIN(N2003) );
and2s1 U498 ( .Q(N2374), .DIN1(N193), .DIN2(N1997) );
and2s1 U499 ( .Q(N2375), .DIN1(N192), .DIN2(N1997) );
and2s1 U500 ( .Q(N2376), .DIN1(N191), .DIN2(N1997) );
and2s1 U501 ( .Q(N2377), .DIN1(N190), .DIN2(N1997) );
and2s1 U502 ( .Q(N2378), .DIN1(N189), .DIN2(N1997) );
and2s1 U503 ( .Q(N2379), .DIN1(N47), .DIN2(N2003) );
and2s1 U504 ( .Q(N2380), .DIN1(N35), .DIN2(N2003) );
and2s1 U505 ( .Q(N2381), .DIN1(N32), .DIN2(N2003) );
and2s1 U506 ( .Q(N2382), .DIN1(N50), .DIN2(N2003) );
and2s1 U507 ( .Q(N2383), .DIN1(N66), .DIN2(N2003) );
hi1s1 U508 ( .Q(N2384), .DIN(N2024) );
hi1s1 U509 ( .Q(N2390), .DIN(N2031) );
and2s1 U510 ( .Q(N2396), .DIN1(N58), .DIN2(N2024) );
and2s1 U511 ( .Q(N2397), .DIN1(N77), .DIN2(N2024) );
and2s1 U512 ( .Q(N2398), .DIN1(N78), .DIN2(N2024) );
and2s1 U513 ( .Q(N2399), .DIN1(N59), .DIN2(N2024) );
and2s1 U514 ( .Q(N2400), .DIN1(N81), .DIN2(N2024) );
and2s1 U515 ( .Q(N2401), .DIN1(N80), .DIN2(N2031) );
and2s1 U516 ( .Q(N2402), .DIN1(N79), .DIN2(N2031) );
and2s1 U517 ( .Q(N2403), .DIN1(N60), .DIN2(N2031) );
and2s1 U518 ( .Q(N2404), .DIN1(N61), .DIN2(N2031) );
and2s1 U519 ( .Q(N2405), .DIN1(N62), .DIN2(N2031) );
hi1s1 U520 ( .Q(N2406), .DIN(N2038) );
hi1s1 U521 ( .Q(N2412), .DIN(N2045) );
and2s1 U522 ( .Q(N2418), .DIN1(N69), .DIN2(N2038) );
and2s1 U523 ( .Q(N2419), .DIN1(N70), .DIN2(N2038) );
and2s1 U524 ( .Q(N2420), .DIN1(N74), .DIN2(N2038) );
and2s1 U525 ( .Q(N2421), .DIN1(N76), .DIN2(N2038) );
and2s1 U526 ( .Q(N2422), .DIN1(N75), .DIN2(N2038) );
and2s1 U527 ( .Q(N2423), .DIN1(N73), .DIN2(N2045) );
and2s1 U528 ( .Q(N2424), .DIN1(N53), .DIN2(N2045) );
and2s1 U529 ( .Q(N2425), .DIN1(N54), .DIN2(N2045) );
and2s1 U530 ( .Q(N2426), .DIN1(N55), .DIN2(N2045) );
and2s1 U531 ( .Q(N2427), .DIN1(N56), .DIN2(N2045) );
and2s1 U532 ( .Q(N2428), .DIN1(N82), .DIN2(N2052) );
and2s1 U533 ( .Q(N2429), .DIN1(N65), .DIN2(N2052) );
and2s1 U534 ( .Q(N2430), .DIN1(N83), .DIN2(N2052) );
and2s1 U535 ( .Q(N2431), .DIN1(N84), .DIN2(N2052) );
and2s1 U536 ( .Q(N2432), .DIN1(N85), .DIN2(N2052) );
and2s1 U537 ( .Q(N2433), .DIN1(N64), .DIN2(N2058) );
and2s1 U538 ( .Q(N2434), .DIN1(N63), .DIN2(N2058) );
and2s1 U539 ( .Q(N2435), .DIN1(N86), .DIN2(N2058) );
and2s1 U540 ( .Q(N2436), .DIN1(N109), .DIN2(N2058) );
and2s1 U541 ( .Q(N2437), .DIN1(N110), .DIN2(N2058) );
and2s1 U542 ( .Q(N2441), .DIN1(N2239), .DIN2(N1119) );
and2s1 U543 ( .Q(N2442), .DIN1(N2240), .DIN2(N1119) );
and2s1 U544 ( .Q(N2446), .DIN1(N2241), .DIN2(N1119) );
and2s1 U545 ( .Q(N2450), .DIN1(N2242), .DIN2(N1119) );
and2s1 U546 ( .Q(N2454), .DIN1(N2243), .DIN2(N1119) );
and2s1 U547 ( .Q(N2458), .DIN1(N2244), .DIN2(N1132) );
and2s1 U548 ( .Q(N2462), .DIN1(N2247), .DIN2(N1141) );
and2s1 U549 ( .Q(N2466), .DIN1(N2248), .DIN2(N1141) );
and2s1 U550 ( .Q(N2470), .DIN1(N2249), .DIN2(N1141) );
and2s1 U551 ( .Q(N2474), .DIN1(N2250), .DIN2(N1141) );
and2s1 U552 ( .Q(N2478), .DIN1(N2251), .DIN2(N1141) );
and2s1 U553 ( .Q(N2482), .DIN1(N2252), .DIN2(N1154) );
and2s1 U554 ( .Q(N2488), .DIN1(N2253), .DIN2(N1154) );
and2s1 U555 ( .Q(N2496), .DIN1(N2254), .DIN2(N1154) );
and2s1 U556 ( .Q(N2502), .DIN1(N2255), .DIN2(N1154) );
and2s1 U557 ( .Q(N2508), .DIN1(N2256), .DIN2(N1154) );
nnd2s1 U558 ( .Q(N2523), .DIN1(N2268), .DIN2(N2111) );
nnd2s1 U559 ( .Q(N2533), .DIN1(N2274), .DIN2(N2115) );
hi1s1 U560 ( .Q(N2537), .DIN(N2235) );
or2s1 U561 ( .Q(N2538), .DIN1(N2278), .DIN2(N1858) );
or2s1 U562 ( .Q(N2542), .DIN1(N2279), .DIN2(N1859) );
or2s1 U563 ( .Q(N2546), .DIN1(N2280), .DIN2(N1860) );
or2s1 U564 ( .Q(N2550), .DIN1(N2281), .DIN2(N1861) );
or2s1 U565 ( .Q(N2554), .DIN1(N2283), .DIN2(N1863) );
or2s1 U566 ( .Q(N2561), .DIN1(N2284), .DIN2(N1864) );
or2s1 U567 ( .Q(N2567), .DIN1(N2285), .DIN2(N1865) );
or2s1 U568 ( .Q(N2573), .DIN1(N2286), .DIN2(N1866) );
or2s1 U569 ( .Q(N2604), .DIN1(N2338), .DIN2(N1927) );
or2s1 U570 ( .Q(N2607), .DIN1(N2339), .DIN2(N1928) );
or2s1 U571 ( .Q(N2611), .DIN1(N2340), .DIN2(N1929) );
or2s1 U572 ( .Q(N2615), .DIN1(N2341), .DIN2(N1930) );
and2s1 U573 ( .Q(N2619), .DIN1(N2348), .DIN2(N1227) );
and2s1 U574 ( .Q(N2626), .DIN1(N2349), .DIN2(N1227) );
and2s1 U575 ( .Q(N2632), .DIN1(N2350), .DIN2(N1227) );
and2s1 U576 ( .Q(N2638), .DIN1(N2351), .DIN2(N1227) );
and2s1 U577 ( .Q(N2644), .DIN1(N2352), .DIN2(N1240) );
nnd2s1 U578 ( .Q(N2650), .DIN1(N2355), .DIN2(N2172) );
nnd2s1 U579 ( .Q(N2653), .DIN1(N1431), .DIN2(N2356) );
or2s1 U580 ( .Q(N2654), .DIN1(N2359), .DIN2(N1990) );
or2s1 U581 ( .Q(N2658), .DIN1(N2360), .DIN2(N1991) );
or2s1 U582 ( .Q(N2662), .DIN1(N2361), .DIN2(N1992) );
or2s1 U583 ( .Q(N2666), .DIN1(N2362), .DIN2(N1993) );
or2s1 U584 ( .Q(N2670), .DIN1(N2363), .DIN2(N1994) );
or2s1 U585 ( .Q(N2674), .DIN1(N2366), .DIN2(N1256) );
or2s1 U586 ( .Q(N2680), .DIN1(N2367), .DIN2(N1256) );
or2s1 U587 ( .Q(N2688), .DIN1(N2374), .DIN2(N2010) );
or2s1 U588 ( .Q(N2692), .DIN1(N2375), .DIN2(N2011) );
or2s1 U589 ( .Q(N2696), .DIN1(N2376), .DIN2(N2012) );
or2s1 U590 ( .Q(N2700), .DIN1(N2377), .DIN2(N2013) );
or2s1 U591 ( .Q(N2704), .DIN1(N2378), .DIN2(N2014) );
and2s1 U592 ( .Q(N2728), .DIN1(N2347), .DIN2(N1227) );
or2s1 U593 ( .Q(N2729), .DIN1(N2429), .DIN2(N2065) );
or2s1 U594 ( .Q(N2733), .DIN1(N2430), .DIN2(N2066) );
or2s1 U595 ( .Q(N2737), .DIN1(N2431), .DIN2(N2067) );
or2s1 U596 ( .Q(N2741), .DIN1(N2432), .DIN2(N2068) );
or2s1 U597 ( .Q(N2745), .DIN1(N2433), .DIN2(N2069) );
or2s1 U598 ( .Q(N2749), .DIN1(N2434), .DIN2(N2070) );
or2s1 U599 ( .Q(N2753), .DIN1(N2435), .DIN2(N2071) );
or2s1 U600 ( .Q(N2757), .DIN1(N2436), .DIN2(N2072) );
or2s1 U601 ( .Q(N2761), .DIN1(N2437), .DIN2(N2073) );
hi1s1 U602 ( .Q(N2765), .DIN(N2231) );
and2s1 U603 ( .Q(N2766), .DIN1(N2354), .DIN2(N1240) );
and2s1 U604 ( .Q(N2769), .DIN1(N2353), .DIN2(N1240) );
and2s1 U605 ( .Q(N2772), .DIN1(N2246), .DIN2(N1132) );
and2s1 U606 ( .Q(N2775), .DIN1(N2245), .DIN2(N1132) );
or2s1 U607 ( .Q(N2778), .DIN1(N2282), .DIN2(N1862) );
or2s1 U608 ( .Q(N2781), .DIN1(N2358), .DIN2(N1989) );
or2s1 U609 ( .Q(N2784), .DIN1(N2365), .DIN2(N1996) );
or2s1 U610 ( .Q(N2787), .DIN1(N2364), .DIN2(N1995) );
or2s1 U611 ( .Q(N2790), .DIN1(N2337), .DIN2(N1926) );
or2s1 U612 ( .Q(N2793), .DIN1(N2277), .DIN2(N1857) );
or2s1 U613 ( .Q(N2796), .DIN1(N2428), .DIN2(N2064) );
and2s1 U614 ( .Q(N2866), .DIN1(N2257), .DIN2(N1537) );
and2s1 U615 ( .Q(N2867), .DIN1(N2257), .DIN2(N1537) );
and2s1 U616 ( .Q(N2868), .DIN1(N2257), .DIN2(N1537) );
and2s1 U617 ( .Q(N2869), .DIN1(N2257), .DIN2(N1537) );
and2s1 U618 ( .Q(N2878), .DIN1(N2269), .DIN2(N1551) );
and2s1 U619 ( .Q(N2913), .DIN1(N204), .DIN2(N2287) );
and2s1 U620 ( .Q(N2914), .DIN1(N203), .DIN2(N2287) );
and2s1 U621 ( .Q(N2915), .DIN1(N202), .DIN2(N2287) );
and2s1 U622 ( .Q(N2916), .DIN1(N201), .DIN2(N2287) );
and2s1 U623 ( .Q(N2917), .DIN1(N200), .DIN2(N2287) );
and2s1 U624 ( .Q(N2918), .DIN1(N235), .DIN2(N2293) );
and2s1 U625 ( .Q(N2919), .DIN1(N234), .DIN2(N2293) );
and2s1 U626 ( .Q(N2920), .DIN1(N233), .DIN2(N2293) );
and2s1 U627 ( .Q(N2921), .DIN1(N232), .DIN2(N2293) );
and2s1 U628 ( .Q(N2922), .DIN1(N231), .DIN2(N2293) );
and2s1 U629 ( .Q(N2923), .DIN1(N197), .DIN2(N2309) );
and2s1 U630 ( .Q(N2924), .DIN1(N187), .DIN2(N2309) );
and2s1 U631 ( .Q(N2925), .DIN1(N196), .DIN2(N2309) );
and2s1 U632 ( .Q(N2926), .DIN1(N195), .DIN2(N2309) );
and2s1 U633 ( .Q(N2927), .DIN1(N194), .DIN2(N2309) );
and2s1 U634 ( .Q(N2928), .DIN1(N227), .DIN2(N2315) );
and2s1 U635 ( .Q(N2929), .DIN1(N217), .DIN2(N2315) );
and2s1 U636 ( .Q(N2930), .DIN1(N226), .DIN2(N2315) );
and2s1 U637 ( .Q(N2931), .DIN1(N225), .DIN2(N2315) );
and2s1 U638 ( .Q(N2932), .DIN1(N224), .DIN2(N2315) );
and2s1 U639 ( .Q(N2933), .DIN1(N239), .DIN2(N2331) );
and2s1 U640 ( .Q(N2934), .DIN1(N229), .DIN2(N2331) );
and2s1 U641 ( .Q(N2935), .DIN1(N238), .DIN2(N2331) );
and2s1 U642 ( .Q(N2936), .DIN1(N237), .DIN2(N2331) );
and2s1 U643 ( .Q(N2937), .DIN1(N236), .DIN2(N2331) );
nnd2s1 U644 ( .Q(N2988), .DIN1(N2653), .DIN2(N2357) );
and2s1 U645 ( .Q(N3005), .DIN1(N223), .DIN2(N2368) );
and2s1 U646 ( .Q(N3006), .DIN1(N222), .DIN2(N2368) );
and2s1 U647 ( .Q(N3007), .DIN1(N221), .DIN2(N2368) );
and2s1 U648 ( .Q(N3008), .DIN1(N220), .DIN2(N2368) );
and2s1 U649 ( .Q(N3009), .DIN1(N219), .DIN2(N2368) );
and2s1 U650 ( .Q(N3020), .DIN1(N812), .DIN2(N2384) );
and2s1 U651 ( .Q(N3021), .DIN1(N814), .DIN2(N2384) );
and2s1 U652 ( .Q(N3022), .DIN1(N821), .DIN2(N2384) );
and2s1 U653 ( .Q(N3023), .DIN1(N827), .DIN2(N2384) );
and2s1 U654 ( .Q(N3024), .DIN1(N833), .DIN2(N2384) );
and2s1 U655 ( .Q(N3025), .DIN1(N839), .DIN2(N2390) );
and2s1 U656 ( .Q(N3026), .DIN1(N845), .DIN2(N2390) );
and2s1 U657 ( .Q(N3027), .DIN1(N853), .DIN2(N2390) );
and2s1 U658 ( .Q(N3028), .DIN1(N859), .DIN2(N2390) );
and2s1 U659 ( .Q(N3029), .DIN1(N865), .DIN2(N2390) );
and2s1 U660 ( .Q(N3032), .DIN1(N758), .DIN2(N2406) );
and2s1 U661 ( .Q(N3033), .DIN1(N759), .DIN2(N2406) );
and2s1 U662 ( .Q(N3034), .DIN1(N762), .DIN2(N2406) );
and2s1 U663 ( .Q(N3035), .DIN1(N768), .DIN2(N2406) );
and2s1 U664 ( .Q(N3036), .DIN1(N774), .DIN2(N2406) );
and2s1 U665 ( .Q(N3037), .DIN1(N780), .DIN2(N2412) );
and2s1 U666 ( .Q(N3038), .DIN1(N786), .DIN2(N2412) );
and2s1 U667 ( .Q(N3039), .DIN1(N794), .DIN2(N2412) );
and2s1 U668 ( .Q(N3040), .DIN1(N800), .DIN2(N2412) );
and2s1 U669 ( .Q(N3041), .DIN1(N806), .DIN2(N2412) );
nb1s1 U670 ( .Q(N3061), .DIN(N2257) );
nb1s1 U671 ( .Q(N3064), .DIN(N2257) );
nb1s1 U672 ( .Q(N3067), .DIN(N2269) );
nb1s1 U673 ( .Q(N3070), .DIN(N2269) );
hi1s1 U674 ( .Q(N3073), .DIN(N2728) );
hi1s1 U675 ( .Q(N3080), .DIN(N2441) );
and2s1 U676 ( .Q(N3096), .DIN1(N666), .DIN2(N2644) );
and2s1 U677 ( .Q(N3097), .DIN1(N660), .DIN2(N2638) );
and2s1 U678 ( .Q(N3101), .DIN1(N1189), .DIN2(N2632) );
and2s1 U679 ( .Q(N3107), .DIN1(N651), .DIN2(N2626) );
and2s1 U680 ( .Q(N3114), .DIN1(N644), .DIN2(N2619) );
and2s1 U681 ( .Q(N3122), .DIN1(N2523), .DIN2(N2257) );
or2s1 U682 ( .Q(N3126), .DIN1(N1167), .DIN2(N2866) );
and2s1 U683 ( .Q(N3130), .DIN1(N2523), .DIN2(N2257) );
or2s1 U684 ( .Q(N3131), .DIN1(N1167), .DIN2(N2869) );
and2s1 U685 ( .Q(N3134), .DIN1(N2523), .DIN2(N2257) );
hi1s1 U686 ( .Q(N3135), .DIN(N2533) );
and2s1 U687 ( .Q(N3136), .DIN1(N666), .DIN2(N2644) );
and2s1 U688 ( .Q(N3137), .DIN1(N660), .DIN2(N2638) );
and2s1 U689 ( .Q(N3140), .DIN1(N1189), .DIN2(N2632) );
and2s1 U690 ( .Q(N3144), .DIN1(N651), .DIN2(N2626) );
and2s1 U691 ( .Q(N3149), .DIN1(N644), .DIN2(N2619) );
and2s1 U692 ( .Q(N3155), .DIN1(N2533), .DIN2(N2269) );
or2s1 U693 ( .Q(N3159), .DIN1(N1174), .DIN2(N2878) );
hi1s1 U694 ( .Q(N3167), .DIN(N2778) );
and2s1 U695 ( .Q(N3168), .DIN1(N609), .DIN2(N2508) );
and2s1 U696 ( .Q(N3169), .DIN1(N604), .DIN2(N2502) );
and2s1 U697 ( .Q(N3173), .DIN1(N742), .DIN2(N2496) );
and2s1 U698 ( .Q(N3178), .DIN1(N734), .DIN2(N2488) );
and2s1 U699 ( .Q(N3184), .DIN1(N599), .DIN2(N2482) );
and2s1 U700 ( .Q(N3185), .DIN1(N727), .DIN2(N2573) );
and2s1 U701 ( .Q(N3189), .DIN1(N721), .DIN2(N2567) );
and2s1 U702 ( .Q(N3195), .DIN1(N715), .DIN2(N2561) );
and2s1 U703 ( .Q(N3202), .DIN1(N708), .DIN2(N2554) );
and2s1 U704 ( .Q(N3210), .DIN1(N609), .DIN2(N2508) );
and2s1 U705 ( .Q(N3211), .DIN1(N604), .DIN2(N2502) );
and2s1 U706 ( .Q(N3215), .DIN1(N742), .DIN2(N2496) );
and2s1 U707 ( .Q(N3221), .DIN1(N2488), .DIN2(N734) );
and2s1 U708 ( .Q(N3228), .DIN1(N599), .DIN2(N2482) );
and2s1 U709 ( .Q(N3229), .DIN1(N727), .DIN2(N2573) );
and2s1 U710 ( .Q(N3232), .DIN1(N721), .DIN2(N2567) );
and2s1 U711 ( .Q(N3236), .DIN1(N715), .DIN2(N2561) );
and2s1 U712 ( .Q(N3241), .DIN1(N708), .DIN2(N2554) );
or2s1 U713 ( .Q(N3247), .DIN1(N2913), .DIN2(N2299) );
or2s1 U714 ( .Q(N3251), .DIN1(N2914), .DIN2(N2300) );
or2s1 U715 ( .Q(N3255), .DIN1(N2915), .DIN2(N2301) );
or2s1 U716 ( .Q(N3259), .DIN1(N2916), .DIN2(N2302) );
or2s1 U717 ( .Q(N3263), .DIN1(N2917), .DIN2(N2303) );
or2s1 U718 ( .Q(N3267), .DIN1(N2918), .DIN2(N2304) );
or2s1 U719 ( .Q(N3273), .DIN1(N2919), .DIN2(N2305) );
or2s1 U720 ( .Q(N3281), .DIN1(N2920), .DIN2(N2306) );
or2s1 U721 ( .Q(N3287), .DIN1(N2921), .DIN2(N2307) );
or2s1 U722 ( .Q(N3293), .DIN1(N2922), .DIN2(N2308) );
or2s1 U723 ( .Q(N3299), .DIN1(N2924), .DIN2(N2322) );
or2s1 U724 ( .Q(N3303), .DIN1(N2925), .DIN2(N2323) );
or2s1 U725 ( .Q(N3307), .DIN1(N2926), .DIN2(N2324) );
or2s1 U726 ( .Q(N3311), .DIN1(N2927), .DIN2(N2325) );
or2s1 U727 ( .Q(N3315), .DIN1(N2929), .DIN2(N2327) );
or2s1 U728 ( .Q(N3322), .DIN1(N2930), .DIN2(N2328) );
or2s1 U729 ( .Q(N3328), .DIN1(N2931), .DIN2(N2329) );
or2s1 U730 ( .Q(N3334), .DIN1(N2932), .DIN2(N2330) );
or2s1 U731 ( .Q(N3340), .DIN1(N2934), .DIN2(N2343) );
or2s1 U732 ( .Q(N3343), .DIN1(N2935), .DIN2(N2344) );
or2s1 U733 ( .Q(N3349), .DIN1(N2936), .DIN2(N2345) );
or2s1 U734 ( .Q(N3355), .DIN1(N2937), .DIN2(N2346) );
and2s1 U735 ( .Q(N3361), .DIN1(N2761), .DIN2(N2478) );
and2s1 U736 ( .Q(N3362), .DIN1(N2757), .DIN2(N2474) );
and2s1 U737 ( .Q(N3363), .DIN1(N2753), .DIN2(N2470) );
and2s1 U738 ( .Q(N3364), .DIN1(N2749), .DIN2(N2466) );
and2s1 U739 ( .Q(N3365), .DIN1(N2745), .DIN2(N2462) );
and2s1 U740 ( .Q(N3366), .DIN1(N2741), .DIN2(N2550) );
and2s1 U741 ( .Q(N3367), .DIN1(N2737), .DIN2(N2546) );
and2s1 U742 ( .Q(N3368), .DIN1(N2733), .DIN2(N2542) );
and2s1 U743 ( .Q(N3369), .DIN1(N2729), .DIN2(N2538) );
and2s1 U744 ( .Q(N3370), .DIN1(N2670), .DIN2(N2458) );
and2s1 U745 ( .Q(N3371), .DIN1(N2666), .DIN2(N2454) );
and2s1 U746 ( .Q(N3372), .DIN1(N2662), .DIN2(N2450) );
and2s1 U747 ( .Q(N3373), .DIN1(N2658), .DIN2(N2446) );
and2s1 U748 ( .Q(N3374), .DIN1(N2654), .DIN2(N2442) );
and2s1 U749 ( .Q(N3375), .DIN1(N2988), .DIN2(N2650) );
and2s1 U750 ( .Q(N3379), .DIN1(N2650), .DIN2(N1966) );
hi1s1 U751 ( .Q(N3380), .DIN(N2781) );
and2s1 U752 ( .Q(N3381), .DIN1(N695), .DIN2(N2604) );
or2s1 U753 ( .Q(N3384), .DIN1(N3005), .DIN2(N2379) );
or2s1 U754 ( .Q(N3390), .DIN1(N3006), .DIN2(N2380) );
or2s1 U755 ( .Q(N3398), .DIN1(N3007), .DIN2(N2381) );
or2s1 U756 ( .Q(N3404), .DIN1(N3008), .DIN2(N2382) );
or2s1 U757 ( .Q(N3410), .DIN1(N3009), .DIN2(N2383) );
or2s1 U758 ( .Q(N3416), .DIN1(N3021), .DIN2(N2397) );
or2s1 U759 ( .Q(N3420), .DIN1(N3022), .DIN2(N2398) );
or2s1 U760 ( .Q(N3424), .DIN1(N3023), .DIN2(N2399) );
or2s1 U761 ( .Q(N3428), .DIN1(N3024), .DIN2(N2400) );
or2s1 U762 ( .Q(N3432), .DIN1(N3025), .DIN2(N2401) );
or2s1 U763 ( .Q(N3436), .DIN1(N3026), .DIN2(N2402) );
or2s1 U764 ( .Q(N3440), .DIN1(N3027), .DIN2(N2403) );
or2s1 U765 ( .Q(N3444), .DIN1(N3028), .DIN2(N2404) );
or2s1 U766 ( .Q(N3448), .DIN1(N3029), .DIN2(N2405) );
hi1s1 U767 ( .Q(N3452), .DIN(N2790) );
hi1s1 U768 ( .Q(N3453), .DIN(N2793) );
or2s1 U769 ( .Q(N3454), .DIN1(N3034), .DIN2(N2420) );
or2s1 U770 ( .Q(N3458), .DIN1(N3035), .DIN2(N2421) );
or2s1 U771 ( .Q(N3462), .DIN1(N3036), .DIN2(N2422) );
or2s1 U772 ( .Q(N3466), .DIN1(N3037), .DIN2(N2423) );
or2s1 U773 ( .Q(N3470), .DIN1(N3038), .DIN2(N2424) );
or2s1 U774 ( .Q(N3474), .DIN1(N3039), .DIN2(N2425) );
or2s1 U775 ( .Q(N3478), .DIN1(N3040), .DIN2(N2426) );
or2s1 U776 ( .Q(N3482), .DIN1(N3041), .DIN2(N2427) );
hi1s1 U777 ( .Q(N3486), .DIN(N2796) );
nb1s1 U778 ( .Q(N3487), .DIN(N2644) );
nb1s1 U779 ( .Q(N3490), .DIN(N2638) );
nb1s1 U780 ( .Q(N3493), .DIN(N2632) );
nb1s1 U781 ( .Q(N3496), .DIN(N2626) );
nb1s1 U782 ( .Q(N3499), .DIN(N2619) );
nb1s1 U783 ( .Q(N3502), .DIN(N2523) );
nor2s1 U784 ( .Q(N3507), .DIN1(N1167), .DIN2(N2868) );
nb1s1 U785 ( .Q(N3510), .DIN(N2523) );
nor2s1 U786 ( .Q(N3515), .DIN1(N644), .DIN2(N2619) );
nb1s1 U787 ( .Q(N3518), .DIN(N2644) );
nb1s1 U788 ( .Q(N3521), .DIN(N2638) );
nb1s1 U789 ( .Q(N3524), .DIN(N2632) );
nb1s1 U790 ( .Q(N3527), .DIN(N2626) );
nb1s1 U791 ( .Q(N3530), .DIN(N2619) );
nb1s1 U792 ( .Q(N3535), .DIN(N2619) );
nb1s1 U793 ( .Q(N3539), .DIN(N2632) );
nb1s1 U794 ( .Q(N3542), .DIN(N2626) );
nb1s1 U795 ( .Q(N3545), .DIN(N2644) );
nb1s1 U796 ( .Q(N3548), .DIN(N2638) );
hi1s1 U797 ( .Q(N3551), .DIN(N2766) );
hi1s1 U798 ( .Q(N3552), .DIN(N2769) );
nb1s1 U799 ( .Q(N3553), .DIN(N2442) );
nb1s1 U800 ( .Q(N3557), .DIN(N2450) );
nb1s1 U801 ( .Q(N3560), .DIN(N2446) );
nb1s1 U802 ( .Q(N3563), .DIN(N2458) );
nb1s1 U803 ( .Q(N3566), .DIN(N2454) );
hi1s1 U804 ( .Q(N3569), .DIN(N2772) );
hi1s1 U805 ( .Q(N3570), .DIN(N2775) );
nb1s1 U806 ( .Q(N3571), .DIN(N2554) );
nb1s1 U807 ( .Q(N3574), .DIN(N2567) );
nb1s1 U808 ( .Q(N3577), .DIN(N2561) );
nb1s1 U809 ( .Q(N3580), .DIN(N2482) );
nb1s1 U810 ( .Q(N3583), .DIN(N2573) );
nb1s1 U811 ( .Q(N3586), .DIN(N2496) );
nb1s1 U812 ( .Q(N3589), .DIN(N2488) );
nb1s1 U813 ( .Q(N3592), .DIN(N2508) );
nb1s1 U814 ( .Q(N3595), .DIN(N2502) );
nb1s1 U815 ( .Q(N3598), .DIN(N2508) );
nb1s1 U816 ( .Q(N3601), .DIN(N2502) );
nb1s1 U817 ( .Q(N3604), .DIN(N2496) );
nb1s1 U818 ( .Q(N3607), .DIN(N2482) );
nb1s1 U819 ( .Q(N3610), .DIN(N2573) );
nb1s1 U820 ( .Q(N3613), .DIN(N2567) );
nb1s1 U821 ( .Q(N3616), .DIN(N2561) );
nb1s1 U822 ( .Q(N3619), .DIN(N2488) );
nb1s1 U823 ( .Q(N3622), .DIN(N2554) );
nor2s1 U824 ( .Q(N3625), .DIN1(N734), .DIN2(N2488) );
nor2s1 U825 ( .Q(N3628), .DIN1(N708), .DIN2(N2554) );
nb1s1 U826 ( .Q(N3631), .DIN(N2508) );
nb1s1 U827 ( .Q(N3634), .DIN(N2502) );
nb1s1 U828 ( .Q(N3637), .DIN(N2496) );
nb1s1 U829 ( .Q(N3640), .DIN(N2488) );
nb1s1 U830 ( .Q(N3643), .DIN(N2482) );
nb1s1 U831 ( .Q(N3646), .DIN(N2573) );
nb1s1 U832 ( .Q(N3649), .DIN(N2567) );
nb1s1 U833 ( .Q(N3652), .DIN(N2561) );
nb1s1 U834 ( .Q(N3655), .DIN(N2554) );
nor2s1 U835 ( .Q(N3658), .DIN1(N2488), .DIN2(N734) );
nb1s1 U836 ( .Q(N3661), .DIN(N2674) );
nb1s1 U837 ( .Q(N3664), .DIN(N2674) );
nb1s1 U838 ( .Q(N3667), .DIN(N2761) );
nb1s1 U839 ( .Q(N3670), .DIN(N2478) );
nb1s1 U840 ( .Q(N3673), .DIN(N2757) );
nb1s1 U841 ( .Q(N3676), .DIN(N2474) );
nb1s1 U842 ( .Q(N3679), .DIN(N2753) );
nb1s1 U843 ( .Q(N3682), .DIN(N2470) );
nb1s1 U844 ( .Q(N3685), .DIN(N2745) );
nb1s1 U845 ( .Q(N3688), .DIN(N2462) );
nb1s1 U846 ( .Q(N3691), .DIN(N2741) );
nb1s1 U847 ( .Q(N3694), .DIN(N2550) );
nb1s1 U848 ( .Q(N3697), .DIN(N2737) );
nb1s1 U849 ( .Q(N3700), .DIN(N2546) );
nb1s1 U850 ( .Q(N3703), .DIN(N2733) );
nb1s1 U851 ( .Q(N3706), .DIN(N2542) );
nb1s1 U852 ( .Q(N3709), .DIN(N2749) );
nb1s1 U853 ( .Q(N3712), .DIN(N2466) );
nb1s1 U854 ( .Q(N3715), .DIN(N2729) );
nb1s1 U855 ( .Q(N3718), .DIN(N2538) );
nb1s1 U856 ( .Q(N3721), .DIN(N2704) );
nb1s1 U857 ( .Q(N3724), .DIN(N2700) );
nb1s1 U858 ( .Q(N3727), .DIN(N2696) );
nb1s1 U859 ( .Q(N3730), .DIN(N2688) );
nb1s1 U860 ( .Q(N3733), .DIN(N2692) );
nb1s1 U861 ( .Q(N3736), .DIN(N2670) );
nb1s1 U862 ( .Q(N3739), .DIN(N2458) );
nb1s1 U863 ( .Q(N3742), .DIN(N2666) );
nb1s1 U864 ( .Q(N3745), .DIN(N2454) );
nb1s1 U865 ( .Q(N3748), .DIN(N2662) );
nb1s1 U866 ( .Q(N3751), .DIN(N2450) );
nb1s1 U867 ( .Q(N3754), .DIN(N2658) );
nb1s1 U868 ( .Q(N3757), .DIN(N2446) );
nb1s1 U869 ( .Q(N3760), .DIN(N2654) );
nb1s1 U870 ( .Q(N3763), .DIN(N2442) );
nb1s1 U871 ( .Q(N3766), .DIN(N2654) );
nb1s1 U872 ( .Q(N3769), .DIN(N2662) );
nb1s1 U873 ( .Q(N3772), .DIN(N2658) );
nb1s1 U874 ( .Q(N3775), .DIN(N2670) );
nb1s1 U875 ( .Q(N3778), .DIN(N2666) );
hi1s1 U876 ( .Q(N3781), .DIN(N2784) );
hi1s1 U877 ( .Q(N3782), .DIN(N2787) );
or2s1 U878 ( .Q(N3783), .DIN1(N2928), .DIN2(N2326) );
or2s1 U879 ( .Q(N3786), .DIN1(N2933), .DIN2(N2342) );
or2s1 U880 ( .Q(N3789), .DIN1(N2923), .DIN2(N2321) );
nb1s1 U881 ( .Q(N3792), .DIN(N2688) );
nb1s1 U882 ( .Q(N3795), .DIN(N2696) );
nb1s1 U883 ( .Q(N3798), .DIN(N2692) );
nb1s1 U884 ( .Q(N3801), .DIN(N2704) );
nb1s1 U885 ( .Q(N3804), .DIN(N2700) );
nb1s1 U886 ( .Q(N3807), .DIN(N2604) );
nb1s1 U887 ( .Q(N3810), .DIN(N2611) );
nb1s1 U888 ( .Q(N3813), .DIN(N2607) );
nb1s1 U889 ( .Q(N3816), .DIN(N2615) );
nb1s1 U890 ( .Q(N3819), .DIN(N2538) );
nb1s1 U891 ( .Q(N3822), .DIN(N2546) );
nb1s1 U892 ( .Q(N3825), .DIN(N2542) );
nb1s1 U893 ( .Q(N3828), .DIN(N2462) );
nb1s1 U894 ( .Q(N3831), .DIN(N2550) );
nb1s1 U895 ( .Q(N3834), .DIN(N2470) );
nb1s1 U896 ( .Q(N3837), .DIN(N2466) );
nb1s1 U897 ( .Q(N3840), .DIN(N2478) );
nb1s1 U898 ( .Q(N3843), .DIN(N2474) );
nb1s1 U899 ( .Q(N3846), .DIN(N2615) );
nb1s1 U900 ( .Q(N3849), .DIN(N2611) );
nb1s1 U901 ( .Q(N3852), .DIN(N2607) );
nb1s1 U902 ( .Q(N3855), .DIN(N2680) );
nb1s1 U903 ( .Q(N3858), .DIN(N2729) );
nb1s1 U904 ( .Q(N3861), .DIN(N2737) );
nb1s1 U905 ( .Q(N3864), .DIN(N2733) );
nb1s1 U906 ( .Q(N3867), .DIN(N2745) );
nb1s1 U907 ( .Q(N3870), .DIN(N2741) );
nb1s1 U908 ( .Q(N3873), .DIN(N2753) );
nb1s1 U909 ( .Q(N3876), .DIN(N2749) );
nb1s1 U910 ( .Q(N3879), .DIN(N2761) );
nb1s1 U911 ( .Q(N3882), .DIN(N2757) );
or2s1 U912 ( .Q(N3885), .DIN1(N3033), .DIN2(N2419) );
or2s1 U913 ( .Q(N3888), .DIN1(N3032), .DIN2(N2418) );
or2s1 U914 ( .Q(N3891), .DIN1(N3020), .DIN2(N2396) );
nnd2s1 U915 ( .Q(N3953), .DIN1(N3067), .DIN2(N2117) );
hi1s1 U916 ( .Q(N3954), .DIN(N3067) );
nnd2s1 U917 ( .Q(N3955), .DIN1(N3070), .DIN2(N2537) );
hi1s1 U918 ( .Q(N3956), .DIN(N3070) );
hi1s1 U919 ( .Q(N3958), .DIN(N3073) );
hi1s1 U920 ( .Q(N3964), .DIN(N3080) );
or2s1 U921 ( .Q(N4193), .DIN1(N1649), .DIN2(N3379) );
or3s1 U922 ( .Q(N4303), .DIN1(N1167), .DIN2(N2867), .DIN3(N3130) );
hi1s1 U923 ( .Q(N4308), .DIN(N3061) );
hi1s1 U924 ( .Q(N4313), .DIN(N3064) );
nnd2s1 U925 ( .Q(N4326), .DIN1(N2769), .DIN2(N3551) );
nnd2s1 U926 ( .Q(N4327), .DIN1(N2766), .DIN2(N3552) );
nnd2s1 U927 ( .Q(N4333), .DIN1(N2775), .DIN2(N3569) );
nnd2s1 U928 ( .Q(N4334), .DIN1(N2772), .DIN2(N3570) );
nnd2s1 U929 ( .Q(N4411), .DIN1(N2787), .DIN2(N3781) );
nnd2s1 U930 ( .Q(N4412), .DIN1(N2784), .DIN2(N3782) );
nnd2s1 U931 ( .Q(N4463), .DIN1(N3487), .DIN2(N1828) );
hi1s1 U932 ( .Q(N4464), .DIN(N3487) );
nnd2s1 U933 ( .Q(N4465), .DIN1(N3490), .DIN2(N1829) );
hi1s1 U934 ( .Q(N4466), .DIN(N3490) );
nnd2s1 U935 ( .Q(N4467), .DIN1(N3493), .DIN2(N2267) );
hi1s1 U936 ( .Q(N4468), .DIN(N3493) );
nnd2s1 U937 ( .Q(N4469), .DIN1(N3496), .DIN2(N1830) );
hi1s1 U938 ( .Q(N4470), .DIN(N3496) );
nnd2s1 U939 ( .Q(N4471), .DIN1(N3499), .DIN2(N1833) );
hi1s1 U940 ( .Q(N4472), .DIN(N3499) );
hi1s1 U941 ( .Q(N4473), .DIN(N3122) );
hi1s1 U942 ( .Q(N4474), .DIN(N3126) );
nnd2s1 U943 ( .Q(N4475), .DIN1(N3518), .DIN2(N1840) );
hi1s1 U944 ( .Q(N4476), .DIN(N3518) );
nnd2s1 U945 ( .Q(N4477), .DIN1(N3521), .DIN2(N1841) );
hi1s1 U946 ( .Q(N4478), .DIN(N3521) );
nnd2s1 U947 ( .Q(N4479), .DIN1(N3524), .DIN2(N2275) );
hi1s1 U948 ( .Q(N4480), .DIN(N3524) );
nnd2s1 U949 ( .Q(N4481), .DIN1(N3527), .DIN2(N1842) );
hi1s1 U950 ( .Q(N4482), .DIN(N3527) );
nnd2s1 U951 ( .Q(N4483), .DIN1(N3530), .DIN2(N1843) );
hi1s1 U952 ( .Q(N4484), .DIN(N3530) );
hi1s1 U953 ( .Q(N4485), .DIN(N3155) );
hi1s1 U954 ( .Q(N4486), .DIN(N3159) );
nnd2s1 U955 ( .Q(N4487), .DIN1(N1721), .DIN2(N3954) );
nnd2s1 U956 ( .Q(N4488), .DIN1(N2235), .DIN2(N3956) );
hi1s1 U957 ( .Q(N4489), .DIN(N3535) );
nnd2s1 U958 ( .Q(N4490), .DIN1(N3535), .DIN2(N3958) );
hi1s1 U959 ( .Q(N4491), .DIN(N3539) );
hi1s1 U960 ( .Q(N4492), .DIN(N3542) );
hi1s1 U961 ( .Q(N4493), .DIN(N3545) );
hi1s1 U962 ( .Q(N4494), .DIN(N3548) );
hi1s1 U963 ( .Q(N4495), .DIN(N3553) );
nnd2s1 U964 ( .Q(N4496), .DIN1(N3553), .DIN2(N3964) );
hi1s1 U965 ( .Q(N4497), .DIN(N3557) );
hi1s1 U966 ( .Q(N4498), .DIN(N3560) );
hi1s1 U967 ( .Q(N4499), .DIN(N3563) );
hi1s1 U968 ( .Q(N4500), .DIN(N3566) );
hi1s1 U969 ( .Q(N4501), .DIN(N3571) );
nnd2s1 U970 ( .Q(N4502), .DIN1(N3571), .DIN2(N3167) );
hi1s1 U971 ( .Q(N4503), .DIN(N3574) );
hi1s1 U972 ( .Q(N4504), .DIN(N3577) );
hi1s1 U973 ( .Q(N4505), .DIN(N3580) );
hi1s1 U974 ( .Q(N4506), .DIN(N3583) );
nnd2s1 U975 ( .Q(N4507), .DIN1(N3598), .DIN2(N1867) );
hi1s1 U976 ( .Q(N4508), .DIN(N3598) );
nnd2s1 U977 ( .Q(N4509), .DIN1(N3601), .DIN2(N1868) );
hi1s1 U978 ( .Q(N4510), .DIN(N3601) );
nnd2s1 U979 ( .Q(N4511), .DIN1(N3604), .DIN2(N1869) );
hi1s1 U980 ( .Q(N4512), .DIN(N3604) );
nnd2s1 U981 ( .Q(N4513), .DIN1(N3607), .DIN2(N1870) );
hi1s1 U982 ( .Q(N4514), .DIN(N3607) );
nnd2s1 U983 ( .Q(N4515), .DIN1(N3610), .DIN2(N1871) );
hi1s1 U984 ( .Q(N4516), .DIN(N3610) );
nnd2s1 U985 ( .Q(N4517), .DIN1(N3613), .DIN2(N1872) );
hi1s1 U986 ( .Q(N4518), .DIN(N3613) );
nnd2s1 U987 ( .Q(N4519), .DIN1(N3616), .DIN2(N1873) );
hi1s1 U988 ( .Q(N4520), .DIN(N3616) );
nnd2s1 U989 ( .Q(N4521), .DIN1(N3619), .DIN2(N1874) );
hi1s1 U990 ( .Q(N4522), .DIN(N3619) );
nnd2s1 U991 ( .Q(N4523), .DIN1(N3622), .DIN2(N1875) );
hi1s1 U992 ( .Q(N4524), .DIN(N3622) );
nnd2s1 U993 ( .Q(N4525), .DIN1(N3631), .DIN2(N1876) );
hi1s1 U994 ( .Q(N4526), .DIN(N3631) );
nnd2s1 U995 ( .Q(N4527), .DIN1(N3634), .DIN2(N1877) );
hi1s1 U996 ( .Q(N4528), .DIN(N3634) );
nnd2s1 U997 ( .Q(N4529), .DIN1(N3637), .DIN2(N1878) );
hi1s1 U998 ( .Q(N4530), .DIN(N3637) );
nnd2s1 U999 ( .Q(N4531), .DIN1(N3640), .DIN2(N1879) );
hi1s1 U1000 ( .Q(N4532), .DIN(N3640) );
nnd2s1 U1001 ( .Q(N4533), .DIN1(N3643), .DIN2(N1880) );
hi1s1 U1002 ( .Q(N4534), .DIN(N3643) );
nnd2s1 U1003 ( .Q(N4535), .DIN1(N3646), .DIN2(N1881) );
hi1s1 U1004 ( .Q(N4536), .DIN(N3646) );
nnd2s1 U1005 ( .Q(N4537), .DIN1(N3649), .DIN2(N1882) );
hi1s1 U1006 ( .Q(N4538), .DIN(N3649) );
nnd2s1 U1007 ( .Q(N4539), .DIN1(N3652), .DIN2(N1883) );
hi1s1 U1008 ( .Q(N4540), .DIN(N3652) );
nnd2s1 U1009 ( .Q(N4541), .DIN1(N3655), .DIN2(N1884) );
hi1s1 U1010 ( .Q(N4542), .DIN(N3655) );
hi1s1 U1011 ( .Q(N4543), .DIN(N3658) );
and2s1 U1012 ( .Q(N4544), .DIN1(N806), .DIN2(N3293) );
and2s1 U1013 ( .Q(N4545), .DIN1(N800), .DIN2(N3287) );
and2s1 U1014 ( .Q(N4549), .DIN1(N794), .DIN2(N3281) );
and2s1 U1015 ( .Q(N4555), .DIN1(N3273), .DIN2(N786) );
and2s1 U1016 ( .Q(N4562), .DIN1(N780), .DIN2(N3267) );
and2s1 U1017 ( .Q(N4563), .DIN1(N774), .DIN2(N3355) );
and2s1 U1018 ( .Q(N4566), .DIN1(N768), .DIN2(N3349) );
and2s1 U1019 ( .Q(N4570), .DIN1(N762), .DIN2(N3343) );
hi1s1 U1020 ( .Q(N4575), .DIN(N3661) );
and2s1 U1021 ( .Q(N4576), .DIN1(N806), .DIN2(N3293) );
and2s1 U1022 ( .Q(N4577), .DIN1(N800), .DIN2(N3287) );
and2s1 U1023 ( .Q(N4581), .DIN1(N794), .DIN2(N3281) );
and2s1 U1024 ( .Q(N4586), .DIN1(N786), .DIN2(N3273) );
and2s1 U1025 ( .Q(N4592), .DIN1(N780), .DIN2(N3267) );
and2s1 U1026 ( .Q(N4593), .DIN1(N774), .DIN2(N3355) );
and2s1 U1027 ( .Q(N4597), .DIN1(N768), .DIN2(N3349) );
and2s1 U1028 ( .Q(N4603), .DIN1(N762), .DIN2(N3343) );
hi1s1 U1029 ( .Q(N4610), .DIN(N3664) );
hi1s1 U1030 ( .Q(N4611), .DIN(N3667) );
hi1s1 U1031 ( .Q(N4612), .DIN(N3670) );
hi1s1 U1032 ( .Q(N4613), .DIN(N3673) );
hi1s1 U1033 ( .Q(N4614), .DIN(N3676) );
hi1s1 U1034 ( .Q(N4615), .DIN(N3679) );
hi1s1 U1035 ( .Q(N4616), .DIN(N3682) );
hi1s1 U1036 ( .Q(N4617), .DIN(N3685) );
hi1s1 U1037 ( .Q(N4618), .DIN(N3688) );
hi1s1 U1038 ( .Q(N4619), .DIN(N3691) );
hi1s1 U1039 ( .Q(N4620), .DIN(N3694) );
hi1s1 U1040 ( .Q(N4621), .DIN(N3697) );
hi1s1 U1041 ( .Q(N4622), .DIN(N3700) );
hi1s1 U1042 ( .Q(N4623), .DIN(N3703) );
hi1s1 U1043 ( .Q(N4624), .DIN(N3706) );
hi1s1 U1044 ( .Q(N4625), .DIN(N3709) );
hi1s1 U1045 ( .Q(N4626), .DIN(N3712) );
hi1s1 U1046 ( .Q(N4627), .DIN(N3715) );
hi1s1 U1047 ( .Q(N4628), .DIN(N3718) );
hi1s1 U1048 ( .Q(N4629), .DIN(N3721) );
and2s1 U1049 ( .Q(N4630), .DIN1(N3448), .DIN2(N2704) );
hi1s1 U1050 ( .Q(N4631), .DIN(N3724) );
and2s1 U1051 ( .Q(N4632), .DIN1(N3444), .DIN2(N2700) );
hi1s1 U1052 ( .Q(N4633), .DIN(N3727) );
and2s1 U1053 ( .Q(N4634), .DIN1(N3440), .DIN2(N2696) );
and2s1 U1054 ( .Q(N4635), .DIN1(N3436), .DIN2(N2692) );
hi1s1 U1055 ( .Q(N4636), .DIN(N3730) );
and2s1 U1056 ( .Q(N4637), .DIN1(N3432), .DIN2(N2688) );
and2s1 U1057 ( .Q(N4638), .DIN1(N3428), .DIN2(N3311) );
and2s1 U1058 ( .Q(N4639), .DIN1(N3424), .DIN2(N3307) );
and2s1 U1059 ( .Q(N4640), .DIN1(N3420), .DIN2(N3303) );
and2s1 U1060 ( .Q(N4641), .DIN1(N3416), .DIN2(N3299) );
hi1s1 U1061 ( .Q(N4642), .DIN(N3733) );
hi1s1 U1062 ( .Q(N4643), .DIN(N3736) );
hi1s1 U1063 ( .Q(N4644), .DIN(N3739) );
hi1s1 U1064 ( .Q(N4645), .DIN(N3742) );
hi1s1 U1065 ( .Q(N4646), .DIN(N3745) );
hi1s1 U1066 ( .Q(N4647), .DIN(N3748) );
hi1s1 U1067 ( .Q(N4648), .DIN(N3751) );
hi1s1 U1068 ( .Q(N4649), .DIN(N3754) );
hi1s1 U1069 ( .Q(N4650), .DIN(N3757) );
hi1s1 U1070 ( .Q(N4651), .DIN(N3760) );
hi1s1 U1071 ( .Q(N4652), .DIN(N3763) );
hi1s1 U1072 ( .Q(N4653), .DIN(N3375) );
and2s1 U1073 ( .Q(N4656), .DIN1(N865), .DIN2(N3410) );
and2s1 U1074 ( .Q(N4657), .DIN1(N859), .DIN2(N3404) );
and2s1 U1075 ( .Q(N4661), .DIN1(N853), .DIN2(N3398) );
and2s1 U1076 ( .Q(N4667), .DIN1(N3390), .DIN2(N845) );
and2s1 U1077 ( .Q(N4674), .DIN1(N839), .DIN2(N3384) );
and2s1 U1078 ( .Q(N4675), .DIN1(N833), .DIN2(N3334) );
and2s1 U1079 ( .Q(N4678), .DIN1(N827), .DIN2(N3328) );
and2s1 U1080 ( .Q(N4682), .DIN1(N821), .DIN2(N3322) );
and2s1 U1081 ( .Q(N4687), .DIN1(N814), .DIN2(N3315) );
hi1s1 U1082 ( .Q(N4693), .DIN(N3766) );
nnd2s1 U1083 ( .Q(N4694), .DIN1(N3766), .DIN2(N3380) );
hi1s1 U1084 ( .Q(N4695), .DIN(N3769) );
hi1s1 U1085 ( .Q(N4696), .DIN(N3772) );
hi1s1 U1086 ( .Q(N4697), .DIN(N3775) );
hi1s1 U1087 ( .Q(N4698), .DIN(N3778) );
hi1s1 U1088 ( .Q(N4699), .DIN(N3783) );
hi1s1 U1089 ( .Q(N4700), .DIN(N3786) );
and2s1 U1090 ( .Q(N4701), .DIN1(N865), .DIN2(N3410) );
and2s1 U1091 ( .Q(N4702), .DIN1(N859), .DIN2(N3404) );
and2s1 U1092 ( .Q(N4706), .DIN1(N853), .DIN2(N3398) );
and2s1 U1093 ( .Q(N4711), .DIN1(N845), .DIN2(N3390) );
and2s1 U1094 ( .Q(N4717), .DIN1(N839), .DIN2(N3384) );
and2s1 U1095 ( .Q(N4718), .DIN1(N833), .DIN2(N3334) );
and2s1 U1096 ( .Q(N4722), .DIN1(N827), .DIN2(N3328) );
and2s1 U1097 ( .Q(N4728), .DIN1(N821), .DIN2(N3322) );
and2s1 U1098 ( .Q(N4735), .DIN1(N814), .DIN2(N3315) );
hi1s1 U1099 ( .Q(N4743), .DIN(N3789) );
hi1s1 U1100 ( .Q(N4744), .DIN(N3792) );
hi1s1 U1101 ( .Q(N4745), .DIN(N3807) );
nnd2s1 U1102 ( .Q(N4746), .DIN1(N3807), .DIN2(N3452) );
hi1s1 U1103 ( .Q(N4747), .DIN(N3810) );
hi1s1 U1104 ( .Q(N4748), .DIN(N3813) );
hi1s1 U1105 ( .Q(N4749), .DIN(N3816) );
hi1s1 U1106 ( .Q(N4750), .DIN(N3819) );
nnd2s1 U1107 ( .Q(N4751), .DIN1(N3819), .DIN2(N3453) );
hi1s1 U1108 ( .Q(N4752), .DIN(N3822) );
hi1s1 U1109 ( .Q(N4753), .DIN(N3825) );
hi1s1 U1110 ( .Q(N4754), .DIN(N3828) );
hi1s1 U1111 ( .Q(N4755), .DIN(N3831) );
and2s1 U1112 ( .Q(N4756), .DIN1(N3482), .DIN2(N3263) );
and2s1 U1113 ( .Q(N4757), .DIN1(N3478), .DIN2(N3259) );
and2s1 U1114 ( .Q(N4758), .DIN1(N3474), .DIN2(N3255) );
and2s1 U1115 ( .Q(N4759), .DIN1(N3470), .DIN2(N3251) );
and2s1 U1116 ( .Q(N4760), .DIN1(N3466), .DIN2(N3247) );
hi1s1 U1117 ( .Q(N4761), .DIN(N3846) );
and2s1 U1118 ( .Q(N4762), .DIN1(N3462), .DIN2(N2615) );
hi1s1 U1119 ( .Q(N4763), .DIN(N3849) );
and2s1 U1120 ( .Q(N4764), .DIN1(N3458), .DIN2(N2611) );
hi1s1 U1121 ( .Q(N4765), .DIN(N3852) );
and2s1 U1122 ( .Q(N4766), .DIN1(N3454), .DIN2(N2607) );
and2s1 U1123 ( .Q(N4767), .DIN1(N2680), .DIN2(N3381) );
hi1s1 U1124 ( .Q(N4768), .DIN(N3855) );
and2s1 U1125 ( .Q(N4769), .DIN1(N3340), .DIN2(N695) );
hi1s1 U1126 ( .Q(N4775), .DIN(N3858) );
nnd2s1 U1127 ( .Q(N4776), .DIN1(N3858), .DIN2(N3486) );
hi1s1 U1128 ( .Q(N4777), .DIN(N3861) );
hi1s1 U1129 ( .Q(N4778), .DIN(N3864) );
hi1s1 U1130 ( .Q(N4779), .DIN(N3867) );
hi1s1 U1131 ( .Q(N4780), .DIN(N3870) );
hi1s1 U1132 ( .Q(N4781), .DIN(N3885) );
hi1s1 U1133 ( .Q(N4782), .DIN(N3888) );
hi1s1 U1134 ( .Q(N4783), .DIN(N3891) );
or2s1 U1135 ( .Q(N4784), .DIN1(N3131), .DIN2(N3134) );
hi1s1 U1136 ( .Q(N4789), .DIN(N3502) );
hi1s1 U1137 ( .Q(N4790), .DIN(N3131) );
hi1s1 U1138 ( .Q(N4793), .DIN(N3507) );
hi1s1 U1139 ( .Q(N4794), .DIN(N3510) );
hi1s1 U1140 ( .Q(N4795), .DIN(N3515) );
nb1s1 U1141 ( .Q(N4796), .DIN(N3114) );
hi1s1 U1142 ( .Q(N4799), .DIN(N3586) );
hi1s1 U1143 ( .Q(N4800), .DIN(N3589) );
hi1s1 U1144 ( .Q(N4801), .DIN(N3592) );
hi1s1 U1145 ( .Q(N4802), .DIN(N3595) );
nnd2s1 U1146 ( .Q(N4803), .DIN1(N4326), .DIN2(N4327) );
nnd2s1 U1147 ( .Q(N4806), .DIN1(N4333), .DIN2(N4334) );
hi1s1 U1148 ( .Q(N4809), .DIN(N3625) );
nb1s1 U1149 ( .Q(N4810), .DIN(N3178) );
hi1s1 U1150 ( .Q(N4813), .DIN(N3628) );
nb1s1 U1151 ( .Q(N4814), .DIN(N3202) );
nb1s1 U1152 ( .Q(N4817), .DIN(N3221) );
nb1s1 U1153 ( .Q(N4820), .DIN(N3293) );
nb1s1 U1154 ( .Q(N4823), .DIN(N3287) );
nb1s1 U1155 ( .Q(N4826), .DIN(N3281) );
nb1s1 U1156 ( .Q(N4829), .DIN(N3273) );
nb1s1 U1157 ( .Q(N4832), .DIN(N3267) );
nb1s1 U1158 ( .Q(N4835), .DIN(N3355) );
nb1s1 U1159 ( .Q(N4838), .DIN(N3349) );
nb1s1 U1160 ( .Q(N4841), .DIN(N3343) );
nor2s1 U1161 ( .Q(N4844), .DIN1(N3273), .DIN2(N786) );
nb1s1 U1162 ( .Q(N4847), .DIN(N3293) );
nb1s1 U1163 ( .Q(N4850), .DIN(N3287) );
nb1s1 U1164 ( .Q(N4853), .DIN(N3281) );
nb1s1 U1165 ( .Q(N4856), .DIN(N3267) );
nb1s1 U1166 ( .Q(N4859), .DIN(N3355) );
nb1s1 U1167 ( .Q(N4862), .DIN(N3349) );
nb1s1 U1168 ( .Q(N4865), .DIN(N3343) );
nb1s1 U1169 ( .Q(N4868), .DIN(N3273) );
nor2s1 U1170 ( .Q(N4871), .DIN1(N786), .DIN2(N3273) );
nb1s1 U1171 ( .Q(N4874), .DIN(N3448) );
nb1s1 U1172 ( .Q(N4877), .DIN(N3444) );
nb1s1 U1173 ( .Q(N4880), .DIN(N3440) );
nb1s1 U1174 ( .Q(N4883), .DIN(N3432) );
nb1s1 U1175 ( .Q(N4886), .DIN(N3428) );
nb1s1 U1176 ( .Q(N4889), .DIN(N3311) );
nb1s1 U1177 ( .Q(N4892), .DIN(N3424) );
nb1s1 U1178 ( .Q(N4895), .DIN(N3307) );
nb1s1 U1179 ( .Q(N4898), .DIN(N3420) );
nb1s1 U1180 ( .Q(N4901), .DIN(N3303) );
nb1s1 U1181 ( .Q(N4904), .DIN(N3436) );
nb1s1 U1182 ( .Q(N4907), .DIN(N3416) );
nb1s1 U1183 ( .Q(N4910), .DIN(N3299) );
nb1s1 U1184 ( .Q(N4913), .DIN(N3410) );
nb1s1 U1185 ( .Q(N4916), .DIN(N3404) );
nb1s1 U1186 ( .Q(N4919), .DIN(N3398) );
nb1s1 U1187 ( .Q(N4922), .DIN(N3390) );
nb1s1 U1188 ( .Q(N4925), .DIN(N3384) );
nb1s1 U1189 ( .Q(N4928), .DIN(N3334) );
nb1s1 U1190 ( .Q(N4931), .DIN(N3328) );
nb1s1 U1191 ( .Q(N4934), .DIN(N3322) );
nb1s1 U1192 ( .Q(N4937), .DIN(N3315) );
nor2s1 U1193 ( .Q(N4940), .DIN1(N3390), .DIN2(N845) );
nb1s1 U1194 ( .Q(N4943), .DIN(N3315) );
nb1s1 U1195 ( .Q(N4946), .DIN(N3328) );
nb1s1 U1196 ( .Q(N4949), .DIN(N3322) );
nb1s1 U1197 ( .Q(N4952), .DIN(N3384) );
nb1s1 U1198 ( .Q(N4955), .DIN(N3334) );
nb1s1 U1199 ( .Q(N4958), .DIN(N3398) );
nb1s1 U1200 ( .Q(N4961), .DIN(N3390) );
nb1s1 U1201 ( .Q(N4964), .DIN(N3410) );
nb1s1 U1202 ( .Q(N4967), .DIN(N3404) );
nb1s1 U1203 ( .Q(N4970), .DIN(N3340) );
nb1s1 U1204 ( .Q(N4973), .DIN(N3349) );
nb1s1 U1205 ( .Q(N4976), .DIN(N3343) );
nb1s1 U1206 ( .Q(N4979), .DIN(N3267) );
nb1s1 U1207 ( .Q(N4982), .DIN(N3355) );
nb1s1 U1208 ( .Q(N4985), .DIN(N3281) );
nb1s1 U1209 ( .Q(N4988), .DIN(N3273) );
nb1s1 U1210 ( .Q(N4991), .DIN(N3293) );
nb1s1 U1211 ( .Q(N4994), .DIN(N3287) );
nnd2s1 U1212 ( .Q(N4997), .DIN1(N4411), .DIN2(N4412) );
nb1s1 U1213 ( .Q(N5000), .DIN(N3410) );
nb1s1 U1214 ( .Q(N5003), .DIN(N3404) );
nb1s1 U1215 ( .Q(N5006), .DIN(N3398) );
nb1s1 U1216 ( .Q(N5009), .DIN(N3384) );
nb1s1 U1217 ( .Q(N5012), .DIN(N3334) );
nb1s1 U1218 ( .Q(N5015), .DIN(N3328) );
nb1s1 U1219 ( .Q(N5018), .DIN(N3322) );
nb1s1 U1220 ( .Q(N5021), .DIN(N3390) );
nb1s1 U1221 ( .Q(N5024), .DIN(N3315) );
nor2s1 U1222 ( .Q(N5027), .DIN1(N845), .DIN2(N3390) );
nor2s1 U1223 ( .Q(N5030), .DIN1(N814), .DIN2(N3315) );
nb1s1 U1224 ( .Q(N5033), .DIN(N3299) );
nb1s1 U1225 ( .Q(N5036), .DIN(N3307) );
nb1s1 U1226 ( .Q(N5039), .DIN(N3303) );
nb1s1 U1227 ( .Q(N5042), .DIN(N3311) );
hi1s1 U1228 ( .Q(N5045), .DIN(N3795) );
hi1s1 U1229 ( .Q(N5046), .DIN(N3798) );
hi1s1 U1230 ( .Q(N5047), .DIN(N3801) );
hi1s1 U1231 ( .Q(N5048), .DIN(N3804) );
nb1s1 U1232 ( .Q(N5049), .DIN(N3247) );
nb1s1 U1233 ( .Q(N5052), .DIN(N3255) );
nb1s1 U1234 ( .Q(N5055), .DIN(N3251) );
nb1s1 U1235 ( .Q(N5058), .DIN(N3263) );
nb1s1 U1236 ( .Q(N5061), .DIN(N3259) );
hi1s1 U1237 ( .Q(N5064), .DIN(N3834) );
hi1s1 U1238 ( .Q(N5065), .DIN(N3837) );
hi1s1 U1239 ( .Q(N5066), .DIN(N3840) );
hi1s1 U1240 ( .Q(N5067), .DIN(N3843) );
nb1s1 U1241 ( .Q(N5068), .DIN(N3482) );
nb1s1 U1242 ( .Q(N5071), .DIN(N3263) );
nb1s1 U1243 ( .Q(N5074), .DIN(N3478) );
nb1s1 U1244 ( .Q(N5077), .DIN(N3259) );
nb1s1 U1245 ( .Q(N5080), .DIN(N3474) );
nb1s1 U1246 ( .Q(N5083), .DIN(N3255) );
nb1s1 U1247 ( .Q(N5086), .DIN(N3466) );
nb1s1 U1248 ( .Q(N5089), .DIN(N3247) );
nb1s1 U1249 ( .Q(N5092), .DIN(N3462) );
nb1s1 U1250 ( .Q(N5095), .DIN(N3458) );
nb1s1 U1251 ( .Q(N5098), .DIN(N3454) );
nb1s1 U1252 ( .Q(N5101), .DIN(N3470) );
nb1s1 U1253 ( .Q(N5104), .DIN(N3251) );
nb1s1 U1254 ( .Q(N5107), .DIN(N3381) );
hi1s1 U1255 ( .Q(N5110), .DIN(N3873) );
hi1s1 U1256 ( .Q(N5111), .DIN(N3876) );
hi1s1 U1257 ( .Q(N5112), .DIN(N3879) );
hi1s1 U1258 ( .Q(N5113), .DIN(N3882) );
nb1s1 U1259 ( .Q(N5114), .DIN(N3458) );
nb1s1 U1260 ( .Q(N5117), .DIN(N3454) );
nb1s1 U1261 ( .Q(N5120), .DIN(N3466) );
nb1s1 U1262 ( .Q(N5123), .DIN(N3462) );
nb1s1 U1263 ( .Q(N5126), .DIN(N3474) );
nb1s1 U1264 ( .Q(N5129), .DIN(N3470) );
nb1s1 U1265 ( .Q(N5132), .DIN(N3482) );
nb1s1 U1266 ( .Q(N5135), .DIN(N3478) );
nb1s1 U1267 ( .Q(N5138), .DIN(N3416) );
nb1s1 U1268 ( .Q(N5141), .DIN(N3424) );
nb1s1 U1269 ( .Q(N5144), .DIN(N3420) );
nb1s1 U1270 ( .Q(N5147), .DIN(N3432) );
nb1s1 U1271 ( .Q(N5150), .DIN(N3428) );
nb1s1 U1272 ( .Q(N5153), .DIN(N3440) );
nb1s1 U1273 ( .Q(N5156), .DIN(N3436) );
nb1s1 U1274 ( .Q(N5159), .DIN(N3448) );
nb1s1 U1275 ( .Q(N5162), .DIN(N3444) );
nnd2s1 U1276 ( .Q(N5165), .DIN1(N4486), .DIN2(N4485) );
nnd2s1 U1277 ( .Q(N5166), .DIN1(N4474), .DIN2(N4473) );
nnd2s1 U1278 ( .Q(N5167), .DIN1(N1290), .DIN2(N4464) );
nnd2s1 U1279 ( .Q(N5168), .DIN1(N1293), .DIN2(N4466) );
nnd2s1 U1280 ( .Q(N5169), .DIN1(N2074), .DIN2(N4468) );
nnd2s1 U1281 ( .Q(N5170), .DIN1(N1296), .DIN2(N4470) );
nnd2s1 U1282 ( .Q(N5171), .DIN1(N1302), .DIN2(N4472) );
nnd2s1 U1283 ( .Q(N5172), .DIN1(N1314), .DIN2(N4476) );
nnd2s1 U1284 ( .Q(N5173), .DIN1(N1317), .DIN2(N4478) );
nnd2s1 U1285 ( .Q(N5174), .DIN1(N2081), .DIN2(N4480) );
nnd2s1 U1286 ( .Q(N5175), .DIN1(N1320), .DIN2(N4482) );
nnd2s1 U1287 ( .Q(N5176), .DIN1(N1323), .DIN2(N4484) );
nnd2s1 U1288 ( .Q(N5177), .DIN1(N3953), .DIN2(N4487) );
nnd2s1 U1289 ( .Q(N5178), .DIN1(N3955), .DIN2(N4488) );
nnd2s1 U1290 ( .Q(N5179), .DIN1(N3073), .DIN2(N4489) );
nnd2s1 U1291 ( .Q(N5180), .DIN1(N3542), .DIN2(N4491) );
nnd2s1 U1292 ( .Q(N5181), .DIN1(N3539), .DIN2(N4492) );
nnd2s1 U1293 ( .Q(N5182), .DIN1(N3548), .DIN2(N4493) );
nnd2s1 U1294 ( .Q(N5183), .DIN1(N3545), .DIN2(N4494) );
nnd2s1 U1295 ( .Q(N5184), .DIN1(N3080), .DIN2(N4495) );
nnd2s1 U1296 ( .Q(N5185), .DIN1(N3560), .DIN2(N4497) );
nnd2s1 U1297 ( .Q(N5186), .DIN1(N3557), .DIN2(N4498) );
nnd2s1 U1298 ( .Q(N5187), .DIN1(N3566), .DIN2(N4499) );
nnd2s1 U1299 ( .Q(N5188), .DIN1(N3563), .DIN2(N4500) );
nnd2s1 U1300 ( .Q(N5189), .DIN1(N2778), .DIN2(N4501) );
nnd2s1 U1301 ( .Q(N5190), .DIN1(N3577), .DIN2(N4503) );
nnd2s1 U1302 ( .Q(N5191), .DIN1(N3574), .DIN2(N4504) );
nnd2s1 U1303 ( .Q(N5192), .DIN1(N3583), .DIN2(N4505) );
nnd2s1 U1304 ( .Q(N5193), .DIN1(N3580), .DIN2(N4506) );
nnd2s1 U1305 ( .Q(N5196), .DIN1(N1326), .DIN2(N4508) );
nnd2s1 U1306 ( .Q(N5197), .DIN1(N1329), .DIN2(N4510) );
nnd2s1 U1307 ( .Q(N5198), .DIN1(N1332), .DIN2(N4512) );
nnd2s1 U1308 ( .Q(N5199), .DIN1(N1335), .DIN2(N4514) );
nnd2s1 U1309 ( .Q(N5200), .DIN1(N1338), .DIN2(N4516) );
nnd2s1 U1310 ( .Q(N5201), .DIN1(N1341), .DIN2(N4518) );
nnd2s1 U1311 ( .Q(N5202), .DIN1(N1344), .DIN2(N4520) );
nnd2s1 U1312 ( .Q(N5203), .DIN1(N1347), .DIN2(N4522) );
nnd2s1 U1313 ( .Q(N5204), .DIN1(N1350), .DIN2(N4524) );
nnd2s1 U1314 ( .Q(N5205), .DIN1(N1353), .DIN2(N4526) );
nnd2s1 U1315 ( .Q(N5206), .DIN1(N1356), .DIN2(N4528) );
nnd2s1 U1316 ( .Q(N5207), .DIN1(N1359), .DIN2(N4530) );
nnd2s1 U1317 ( .Q(N5208), .DIN1(N1362), .DIN2(N4532) );
nnd2s1 U1318 ( .Q(N5209), .DIN1(N1365), .DIN2(N4534) );
nnd2s1 U1319 ( .Q(N5210), .DIN1(N1368), .DIN2(N4536) );
nnd2s1 U1320 ( .Q(N5211), .DIN1(N1371), .DIN2(N4538) );
nnd2s1 U1321 ( .Q(N5212), .DIN1(N1374), .DIN2(N4540) );
nnd2s1 U1322 ( .Q(N5213), .DIN1(N1377), .DIN2(N4542) );
nnd2s1 U1323 ( .Q(N5283), .DIN1(N3670), .DIN2(N4611) );
nnd2s1 U1324 ( .Q(N5284), .DIN1(N3667), .DIN2(N4612) );
nnd2s1 U1325 ( .Q(N5285), .DIN1(N3676), .DIN2(N4613) );
nnd2s1 U1326 ( .Q(N5286), .DIN1(N3673), .DIN2(N4614) );
nnd2s1 U1327 ( .Q(N5287), .DIN1(N3682), .DIN2(N4615) );
nnd2s1 U1328 ( .Q(N5288), .DIN1(N3679), .DIN2(N4616) );
nnd2s1 U1329 ( .Q(N5289), .DIN1(N3688), .DIN2(N4617) );
nnd2s1 U1330 ( .Q(N5290), .DIN1(N3685), .DIN2(N4618) );
nnd2s1 U1331 ( .Q(N5291), .DIN1(N3694), .DIN2(N4619) );
nnd2s1 U1332 ( .Q(N5292), .DIN1(N3691), .DIN2(N4620) );
nnd2s1 U1333 ( .Q(N5293), .DIN1(N3700), .DIN2(N4621) );
nnd2s1 U1334 ( .Q(N5294), .DIN1(N3697), .DIN2(N4622) );
nnd2s1 U1335 ( .Q(N5295), .DIN1(N3706), .DIN2(N4623) );
nnd2s1 U1336 ( .Q(N5296), .DIN1(N3703), .DIN2(N4624) );
nnd2s1 U1337 ( .Q(N5297), .DIN1(N3712), .DIN2(N4625) );
nnd2s1 U1338 ( .Q(N5298), .DIN1(N3709), .DIN2(N4626) );
nnd2s1 U1339 ( .Q(N5299), .DIN1(N3718), .DIN2(N4627) );
nnd2s1 U1340 ( .Q(N5300), .DIN1(N3715), .DIN2(N4628) );
nnd2s1 U1341 ( .Q(N5314), .DIN1(N3739), .DIN2(N4643) );
nnd2s1 U1342 ( .Q(N5315), .DIN1(N3736), .DIN2(N4644) );
nnd2s1 U1343 ( .Q(N5316), .DIN1(N3745), .DIN2(N4645) );
nnd2s1 U1344 ( .Q(N5317), .DIN1(N3742), .DIN2(N4646) );
nnd2s1 U1345 ( .Q(N5318), .DIN1(N3751), .DIN2(N4647) );
nnd2s1 U1346 ( .Q(N5319), .DIN1(N3748), .DIN2(N4648) );
nnd2s1 U1347 ( .Q(N5320), .DIN1(N3757), .DIN2(N4649) );
nnd2s1 U1348 ( .Q(N5321), .DIN1(N3754), .DIN2(N4650) );
nnd2s1 U1349 ( .Q(N5322), .DIN1(N3763), .DIN2(N4651) );
nnd2s1 U1350 ( .Q(N5323), .DIN1(N3760), .DIN2(N4652) );
hi1s1 U1351 ( .Q(N5324), .DIN(N4193) );
nnd2s1 U1352 ( .Q(N5363), .DIN1(N2781), .DIN2(N4693) );
nnd2s1 U1353 ( .Q(N5364), .DIN1(N3772), .DIN2(N4695) );
nnd2s1 U1354 ( .Q(N5365), .DIN1(N3769), .DIN2(N4696) );
nnd2s1 U1355 ( .Q(N5366), .DIN1(N3778), .DIN2(N4697) );
nnd2s1 U1356 ( .Q(N5367), .DIN1(N3775), .DIN2(N4698) );
nnd2s1 U1357 ( .Q(N5425), .DIN1(N2790), .DIN2(N4745) );
nnd2s1 U1358 ( .Q(N5426), .DIN1(N3813), .DIN2(N4747) );
nnd2s1 U1359 ( .Q(N5427), .DIN1(N3810), .DIN2(N4748) );
nnd2s1 U1360 ( .Q(N5429), .DIN1(N2793), .DIN2(N4750) );
nnd2s1 U1361 ( .Q(N5430), .DIN1(N3825), .DIN2(N4752) );
nnd2s1 U1362 ( .Q(N5431), .DIN1(N3822), .DIN2(N4753) );
nnd2s1 U1363 ( .Q(N5432), .DIN1(N3831), .DIN2(N4754) );
nnd2s1 U1364 ( .Q(N5433), .DIN1(N3828), .DIN2(N4755) );
nnd2s1 U1365 ( .Q(N5451), .DIN1(N2796), .DIN2(N4775) );
nnd2s1 U1366 ( .Q(N5452), .DIN1(N3864), .DIN2(N4777) );
nnd2s1 U1367 ( .Q(N5453), .DIN1(N3861), .DIN2(N4778) );
nnd2s1 U1368 ( .Q(N5454), .DIN1(N3870), .DIN2(N4779) );
nnd2s1 U1369 ( .Q(N5455), .DIN1(N3867), .DIN2(N4780) );
nnd2s1 U1370 ( .Q(N5456), .DIN1(N3888), .DIN2(N4781) );
nnd2s1 U1371 ( .Q(N5457), .DIN1(N3885), .DIN2(N4782) );
hi1s1 U1372 ( .Q(N5469), .DIN(N4303) );
nnd2s1 U1373 ( .Q(N5474), .DIN1(N3589), .DIN2(N4799) );
nnd2s1 U1374 ( .Q(N5475), .DIN1(N3586), .DIN2(N4800) );
nnd2s1 U1375 ( .Q(N5476), .DIN1(N3595), .DIN2(N4801) );
nnd2s1 U1376 ( .Q(N5477), .DIN1(N3592), .DIN2(N4802) );
nnd2s1 U1377 ( .Q(N5571), .DIN1(N3798), .DIN2(N5045) );
nnd2s1 U1378 ( .Q(N5572), .DIN1(N3795), .DIN2(N5046) );
nnd2s1 U1379 ( .Q(N5573), .DIN1(N3804), .DIN2(N5047) );
nnd2s1 U1380 ( .Q(N5574), .DIN1(N3801), .DIN2(N5048) );
nnd2s1 U1381 ( .Q(N5584), .DIN1(N3837), .DIN2(N5064) );
nnd2s1 U1382 ( .Q(N5585), .DIN1(N3834), .DIN2(N5065) );
nnd2s1 U1383 ( .Q(N5586), .DIN1(N3843), .DIN2(N5066) );
nnd2s1 U1384 ( .Q(N5587), .DIN1(N3840), .DIN2(N5067) );
nnd2s1 U1385 ( .Q(N5602), .DIN1(N3876), .DIN2(N5110) );
nnd2s1 U1386 ( .Q(N5603), .DIN1(N3873), .DIN2(N5111) );
nnd2s1 U1387 ( .Q(N5604), .DIN1(N3882), .DIN2(N5112) );
nnd2s1 U1388 ( .Q(N5605), .DIN1(N3879), .DIN2(N5113) );
nnd2s1 U1389 ( .Q(N5631), .DIN1(N5324), .DIN2(N4653) );
nnd2s1 U1390 ( .Q(N5632), .DIN1(N4463), .DIN2(N5167) );
nnd2s1 U1391 ( .Q(N5640), .DIN1(N4465), .DIN2(N5168) );
nnd2s1 U1392 ( .Q(N5654), .DIN1(N4467), .DIN2(N5169) );
nnd2s1 U1393 ( .Q(N5670), .DIN1(N4469), .DIN2(N5170) );
nnd2s1 U1394 ( .Q(N5683), .DIN1(N4471), .DIN2(N5171) );
nnd2s1 U1395 ( .Q(N5690), .DIN1(N4475), .DIN2(N5172) );
nnd2s1 U1396 ( .Q(N5697), .DIN1(N4477), .DIN2(N5173) );
nnd2s1 U1397 ( .Q(N5707), .DIN1(N4479), .DIN2(N5174) );
nnd2s1 U1398 ( .Q(N5718), .DIN1(N4481), .DIN2(N5175) );
nnd2s1 U1399 ( .Q(N5728), .DIN1(N4483), .DIN2(N5176) );
hi1s1 U1400 ( .Q(N5735), .DIN(N5177) );
nnd2s1 U1401 ( .Q(N5736), .DIN1(N5179), .DIN2(N4490) );
nnd2s1 U1402 ( .Q(N5740), .DIN1(N5180), .DIN2(N5181) );
nnd2s1 U1403 ( .Q(N5744), .DIN1(N5182), .DIN2(N5183) );
nnd2s1 U1404 ( .Q(N5747), .DIN1(N5184), .DIN2(N4496) );
nnd2s1 U1405 ( .Q(N5751), .DIN1(N5185), .DIN2(N5186) );
nnd2s1 U1406 ( .Q(N5755), .DIN1(N5187), .DIN2(N5188) );
nnd2s1 U1407 ( .Q(N5758), .DIN1(N5189), .DIN2(N4502) );
nnd2s1 U1408 ( .Q(N5762), .DIN1(N5190), .DIN2(N5191) );
nnd2s1 U1409 ( .Q(N5766), .DIN1(N5192), .DIN2(N5193) );
hi1s1 U1410 ( .Q(N5769), .DIN(N4803) );
hi1s1 U1411 ( .Q(N5770), .DIN(N4806) );
nnd2s1 U1412 ( .Q(N5771), .DIN1(N4507), .DIN2(N5196) );
nnd2s1 U1413 ( .Q(N5778), .DIN1(N4509), .DIN2(N5197) );
nnd2s1 U1414 ( .Q(N5789), .DIN1(N4511), .DIN2(N5198) );
nnd2s1 U1415 ( .Q(N5799), .DIN1(N4513), .DIN2(N5199) );
nnd2s1 U1416 ( .Q(N5807), .DIN1(N4515), .DIN2(N5200) );
nnd2s1 U1417 ( .Q(N5821), .DIN1(N4517), .DIN2(N5201) );
nnd2s1 U1418 ( .Q(N5837), .DIN1(N4519), .DIN2(N5202) );
nnd2s1 U1419 ( .Q(N5850), .DIN1(N4521), .DIN2(N5203) );
nnd2s1 U1420 ( .Q(N5856), .DIN1(N4523), .DIN2(N5204) );
nnd2s1 U1421 ( .Q(N5863), .DIN1(N4525), .DIN2(N5205) );
nnd2s1 U1422 ( .Q(N5870), .DIN1(N4527), .DIN2(N5206) );
nnd2s1 U1423 ( .Q(N5881), .DIN1(N4529), .DIN2(N5207) );
nnd2s1 U1424 ( .Q(N5892), .DIN1(N4531), .DIN2(N5208) );
nnd2s1 U1425 ( .Q(N5898), .DIN1(N4533), .DIN2(N5209) );
nnd2s1 U1426 ( .Q(N5905), .DIN1(N4535), .DIN2(N5210) );
nnd2s1 U1427 ( .Q(N5915), .DIN1(N4537), .DIN2(N5211) );
nnd2s1 U1428 ( .Q(N5926), .DIN1(N4539), .DIN2(N5212) );
nnd2s1 U1429 ( .Q(N5936), .DIN1(N4541), .DIN2(N5213) );
hi1s1 U1430 ( .Q(N5943), .DIN(N4817) );
nnd2s1 U1431 ( .Q(N5944), .DIN1(N4820), .DIN2(N1931) );
hi1s1 U1432 ( .Q(N5945), .DIN(N4820) );
nnd2s1 U1433 ( .Q(N5946), .DIN1(N4823), .DIN2(N1932) );
hi1s1 U1434 ( .Q(N5947), .DIN(N4823) );
nnd2s1 U1435 ( .Q(N5948), .DIN1(N4826), .DIN2(N1933) );
hi1s1 U1436 ( .Q(N5949), .DIN(N4826) );
nnd2s1 U1437 ( .Q(N5950), .DIN1(N4829), .DIN2(N1934) );
hi1s1 U1438 ( .Q(N5951), .DIN(N4829) );
nnd2s1 U1439 ( .Q(N5952), .DIN1(N4832), .DIN2(N1935) );
hi1s1 U1440 ( .Q(N5953), .DIN(N4832) );
nnd2s1 U1441 ( .Q(N5954), .DIN1(N4835), .DIN2(N1936) );
hi1s1 U1442 ( .Q(N5955), .DIN(N4835) );
nnd2s1 U1443 ( .Q(N5956), .DIN1(N4838), .DIN2(N1937) );
hi1s1 U1444 ( .Q(N5957), .DIN(N4838) );
nnd2s1 U1445 ( .Q(N5958), .DIN1(N4841), .DIN2(N1938) );
hi1s1 U1446 ( .Q(N5959), .DIN(N4841) );
and2s1 U1447 ( .Q(N5960), .DIN1(N2674), .DIN2(N4769) );
hi1s1 U1448 ( .Q(N5966), .DIN(N4844) );
nnd2s1 U1449 ( .Q(N5967), .DIN1(N4847), .DIN2(N1939) );
hi1s1 U1450 ( .Q(N5968), .DIN(N4847) );
nnd2s1 U1451 ( .Q(N5969), .DIN1(N4850), .DIN2(N1940) );
hi1s1 U1452 ( .Q(N5970), .DIN(N4850) );
nnd2s1 U1453 ( .Q(N5971), .DIN1(N4853), .DIN2(N1941) );
hi1s1 U1454 ( .Q(N5972), .DIN(N4853) );
nnd2s1 U1455 ( .Q(N5973), .DIN1(N4856), .DIN2(N1942) );
hi1s1 U1456 ( .Q(N5974), .DIN(N4856) );
nnd2s1 U1457 ( .Q(N5975), .DIN1(N4859), .DIN2(N1943) );
hi1s1 U1458 ( .Q(N5976), .DIN(N4859) );
nnd2s1 U1459 ( .Q(N5977), .DIN1(N4862), .DIN2(N1944) );
hi1s1 U1460 ( .Q(N5978), .DIN(N4862) );
nnd2s1 U1461 ( .Q(N5979), .DIN1(N4865), .DIN2(N1945) );
hi1s1 U1462 ( .Q(N5980), .DIN(N4865) );
and2s1 U1463 ( .Q(N5981), .DIN1(N2674), .DIN2(N4769) );
nnd2s1 U1464 ( .Q(N5989), .DIN1(N4868), .DIN2(N1946) );
hi1s1 U1465 ( .Q(N5990), .DIN(N4868) );
nnd2s1 U1466 ( .Q(N5991), .DIN1(N5283), .DIN2(N5284) );
nnd2s1 U1467 ( .Q(N5996), .DIN1(N5285), .DIN2(N5286) );
nnd2s1 U1468 ( .Q(N6000), .DIN1(N5287), .DIN2(N5288) );
nnd2s1 U1469 ( .Q(N6003), .DIN1(N5289), .DIN2(N5290) );
nnd2s1 U1470 ( .Q(N6009), .DIN1(N5291), .DIN2(N5292) );
nnd2s1 U1471 ( .Q(N6014), .DIN1(N5293), .DIN2(N5294) );
nnd2s1 U1472 ( .Q(N6018), .DIN1(N5295), .DIN2(N5296) );
nnd2s1 U1473 ( .Q(N6021), .DIN1(N5297), .DIN2(N5298) );
nnd2s1 U1474 ( .Q(N6022), .DIN1(N5299), .DIN2(N5300) );
hi1s1 U1475 ( .Q(N6023), .DIN(N4874) );
nnd2s1 U1476 ( .Q(N6024), .DIN1(N4874), .DIN2(N4629) );
hi1s1 U1477 ( .Q(N6025), .DIN(N4877) );
nnd2s1 U1478 ( .Q(N6026), .DIN1(N4877), .DIN2(N4631) );
hi1s1 U1479 ( .Q(N6027), .DIN(N4880) );
nnd2s1 U1480 ( .Q(N6028), .DIN1(N4880), .DIN2(N4633) );
hi1s1 U1481 ( .Q(N6029), .DIN(N4883) );
nnd2s1 U1482 ( .Q(N6030), .DIN1(N4883), .DIN2(N4636) );
hi1s1 U1483 ( .Q(N6031), .DIN(N4886) );
hi1s1 U1484 ( .Q(N6032), .DIN(N4889) );
hi1s1 U1485 ( .Q(N6033), .DIN(N4892) );
hi1s1 U1486 ( .Q(N6034), .DIN(N4895) );
hi1s1 U1487 ( .Q(N6035), .DIN(N4898) );
hi1s1 U1488 ( .Q(N6036), .DIN(N4901) );
hi1s1 U1489 ( .Q(N6037), .DIN(N4904) );
nnd2s1 U1490 ( .Q(N6038), .DIN1(N4904), .DIN2(N4642) );
hi1s1 U1491 ( .Q(N6039), .DIN(N4907) );
hi1s1 U1492 ( .Q(N6040), .DIN(N4910) );
nnd2s1 U1493 ( .Q(N6041), .DIN1(N5314), .DIN2(N5315) );
nnd2s1 U1494 ( .Q(N6047), .DIN1(N5316), .DIN2(N5317) );
nnd2s1 U1495 ( .Q(N6052), .DIN1(N5318), .DIN2(N5319) );
nnd2s1 U1496 ( .Q(N6056), .DIN1(N5320), .DIN2(N5321) );
nnd2s1 U1497 ( .Q(N6059), .DIN1(N5322), .DIN2(N5323) );
nnd2s1 U1498 ( .Q(N6060), .DIN1(N4913), .DIN2(N1968) );
hi1s1 U1499 ( .Q(N6061), .DIN(N4913) );
nnd2s1 U1500 ( .Q(N6062), .DIN1(N4916), .DIN2(N1969) );
hi1s1 U1501 ( .Q(N6063), .DIN(N4916) );
nnd2s1 U1502 ( .Q(N6064), .DIN1(N4919), .DIN2(N1970) );
hi1s1 U1503 ( .Q(N6065), .DIN(N4919) );
nnd2s1 U1504 ( .Q(N6066), .DIN1(N4922), .DIN2(N1971) );
hi1s1 U1505 ( .Q(N6067), .DIN(N4922) );
nnd2s1 U1506 ( .Q(N6068), .DIN1(N4925), .DIN2(N1972) );
hi1s1 U1507 ( .Q(N6069), .DIN(N4925) );
nnd2s1 U1508 ( .Q(N6070), .DIN1(N4928), .DIN2(N1973) );
hi1s1 U1509 ( .Q(N6071), .DIN(N4928) );
nnd2s1 U1510 ( .Q(N6072), .DIN1(N4931), .DIN2(N1974) );
hi1s1 U1511 ( .Q(N6073), .DIN(N4931) );
nnd2s1 U1512 ( .Q(N6074), .DIN1(N4934), .DIN2(N1975) );
hi1s1 U1513 ( .Q(N6075), .DIN(N4934) );
nnd2s1 U1514 ( .Q(N6076), .DIN1(N4937), .DIN2(N1976) );
hi1s1 U1515 ( .Q(N6077), .DIN(N4937) );
hi1s1 U1516 ( .Q(N6078), .DIN(N4940) );
nnd2s1 U1517 ( .Q(N6079), .DIN1(N5363), .DIN2(N4694) );
nnd2s1 U1518 ( .Q(N6083), .DIN1(N5364), .DIN2(N5365) );
nnd2s1 U1519 ( .Q(N6087), .DIN1(N5366), .DIN2(N5367) );
hi1s1 U1520 ( .Q(N6090), .DIN(N4943) );
nnd2s1 U1521 ( .Q(N6091), .DIN1(N4943), .DIN2(N4699) );
hi1s1 U1522 ( .Q(N6092), .DIN(N4946) );
hi1s1 U1523 ( .Q(N6093), .DIN(N4949) );
hi1s1 U1524 ( .Q(N6094), .DIN(N4952) );
hi1s1 U1525 ( .Q(N6095), .DIN(N4955) );
hi1s1 U1526 ( .Q(N6096), .DIN(N4970) );
nnd2s1 U1527 ( .Q(N6097), .DIN1(N4970), .DIN2(N4700) );
hi1s1 U1528 ( .Q(N6098), .DIN(N4973) );
hi1s1 U1529 ( .Q(N6099), .DIN(N4976) );
hi1s1 U1530 ( .Q(N6100), .DIN(N4979) );
hi1s1 U1531 ( .Q(N6101), .DIN(N4982) );
hi1s1 U1532 ( .Q(N6102), .DIN(N4997) );
nnd2s1 U1533 ( .Q(N6103), .DIN1(N5000), .DIN2(N2015) );
hi1s1 U1534 ( .Q(N6104), .DIN(N5000) );
nnd2s1 U1535 ( .Q(N6105), .DIN1(N5003), .DIN2(N2016) );
hi1s1 U1536 ( .Q(N6106), .DIN(N5003) );
nnd2s1 U1537 ( .Q(N6107), .DIN1(N5006), .DIN2(N2017) );
hi1s1 U1538 ( .Q(N6108), .DIN(N5006) );
nnd2s1 U1539 ( .Q(N6109), .DIN1(N5009), .DIN2(N2018) );
hi1s1 U1540 ( .Q(N6110), .DIN(N5009) );
nnd2s1 U1541 ( .Q(N6111), .DIN1(N5012), .DIN2(N2019) );
hi1s1 U1542 ( .Q(N6112), .DIN(N5012) );
nnd2s1 U1543 ( .Q(N6113), .DIN1(N5015), .DIN2(N2020) );
hi1s1 U1544 ( .Q(N6114), .DIN(N5015) );
nnd2s1 U1545 ( .Q(N6115), .DIN1(N5018), .DIN2(N2021) );
hi1s1 U1546 ( .Q(N6116), .DIN(N5018) );
nnd2s1 U1547 ( .Q(N6117), .DIN1(N5021), .DIN2(N2022) );
hi1s1 U1548 ( .Q(N6118), .DIN(N5021) );
nnd2s1 U1549 ( .Q(N6119), .DIN1(N5024), .DIN2(N2023) );
hi1s1 U1550 ( .Q(N6120), .DIN(N5024) );
hi1s1 U1551 ( .Q(N6121), .DIN(N5033) );
nnd2s1 U1552 ( .Q(N6122), .DIN1(N5033), .DIN2(N4743) );
hi1s1 U1553 ( .Q(N6123), .DIN(N5036) );
hi1s1 U1554 ( .Q(N6124), .DIN(N5039) );
nnd2s1 U1555 ( .Q(N6125), .DIN1(N5042), .DIN2(N4744) );
hi1s1 U1556 ( .Q(N6126), .DIN(N5042) );
nnd2s1 U1557 ( .Q(N6127), .DIN1(N5425), .DIN2(N4746) );
nnd2s1 U1558 ( .Q(N6131), .DIN1(N5426), .DIN2(N5427) );
hi1s1 U1559 ( .Q(N6135), .DIN(N5049) );
nnd2s1 U1560 ( .Q(N6136), .DIN1(N5049), .DIN2(N4749) );
nnd2s1 U1561 ( .Q(N6137), .DIN1(N5429), .DIN2(N4751) );
nnd2s1 U1562 ( .Q(N6141), .DIN1(N5430), .DIN2(N5431) );
nnd2s1 U1563 ( .Q(N6145), .DIN1(N5432), .DIN2(N5433) );
hi1s1 U1564 ( .Q(N6148), .DIN(N5068) );
hi1s1 U1565 ( .Q(N6149), .DIN(N5071) );
hi1s1 U1566 ( .Q(N6150), .DIN(N5074) );
hi1s1 U1567 ( .Q(N6151), .DIN(N5077) );
hi1s1 U1568 ( .Q(N6152), .DIN(N5080) );
hi1s1 U1569 ( .Q(N6153), .DIN(N5083) );
hi1s1 U1570 ( .Q(N6154), .DIN(N5086) );
hi1s1 U1571 ( .Q(N6155), .DIN(N5089) );
hi1s1 U1572 ( .Q(N6156), .DIN(N5092) );
nnd2s1 U1573 ( .Q(N6157), .DIN1(N5092), .DIN2(N4761) );
hi1s1 U1574 ( .Q(N6158), .DIN(N5095) );
nnd2s1 U1575 ( .Q(N6159), .DIN1(N5095), .DIN2(N4763) );
hi1s1 U1576 ( .Q(N6160), .DIN(N5098) );
nnd2s1 U1577 ( .Q(N6161), .DIN1(N5098), .DIN2(N4765) );
hi1s1 U1578 ( .Q(N6162), .DIN(N5101) );
hi1s1 U1579 ( .Q(N6163), .DIN(N5104) );
nnd2s1 U1580 ( .Q(N6164), .DIN1(N5107), .DIN2(N4768) );
hi1s1 U1581 ( .Q(N6165), .DIN(N5107) );
nnd2s1 U1582 ( .Q(N6166), .DIN1(N5451), .DIN2(N4776) );
nnd2s1 U1583 ( .Q(N6170), .DIN1(N5452), .DIN2(N5453) );
nnd2s1 U1584 ( .Q(N6174), .DIN1(N5454), .DIN2(N5455) );
nnd2s1 U1585 ( .Q(N6177), .DIN1(N5456), .DIN2(N5457) );
hi1s1 U1586 ( .Q(N6181), .DIN(N5114) );
hi1s1 U1587 ( .Q(N6182), .DIN(N5117) );
hi1s1 U1588 ( .Q(N6183), .DIN(N5120) );
hi1s1 U1589 ( .Q(N6184), .DIN(N5123) );
hi1s1 U1590 ( .Q(N6185), .DIN(N5138) );
nnd2s1 U1591 ( .Q(N6186), .DIN1(N5138), .DIN2(N4783) );
hi1s1 U1592 ( .Q(N6187), .DIN(N5141) );
hi1s1 U1593 ( .Q(N6188), .DIN(N5144) );
hi1s1 U1594 ( .Q(N6189), .DIN(N5147) );
hi1s1 U1595 ( .Q(N6190), .DIN(N5150) );
hi1s1 U1596 ( .Q(N6191), .DIN(N4784) );
nnd2s1 U1597 ( .Q(N6192), .DIN1(N4784), .DIN2(N2230) );
hi1s1 U1598 ( .Q(N6193), .DIN(N4790) );
nnd2s1 U1599 ( .Q(N6194), .DIN1(N4790), .DIN2(N2765) );
hi1s1 U1600 ( .Q(N6195), .DIN(N4796) );
nnd2s1 U1601 ( .Q(N6196), .DIN1(N5476), .DIN2(N5477) );
nnd2s1 U1602 ( .Q(N6199), .DIN1(N5474), .DIN2(N5475) );
hi1s1 U1603 ( .Q(N6202), .DIN(N4810) );
hi1s1 U1604 ( .Q(N6203), .DIN(N4814) );
nb1s1 U1605 ( .Q(N6204), .DIN(N4769) );
nb1s1 U1606 ( .Q(N6207), .DIN(N4555) );
nb1s1 U1607 ( .Q(N6210), .DIN(N4769) );
hi1s1 U1608 ( .Q(N6213), .DIN(N4871) );
nb1s1 U1609 ( .Q(N6214), .DIN(N4586) );
nor2s1 U1610 ( .Q(N6217), .DIN1(N2674), .DIN2(N4769) );
nb1s1 U1611 ( .Q(N6220), .DIN(N4667) );
hi1s1 U1612 ( .Q(N6223), .DIN(N4958) );
hi1s1 U1613 ( .Q(N6224), .DIN(N4961) );
hi1s1 U1614 ( .Q(N6225), .DIN(N4964) );
hi1s1 U1615 ( .Q(N6226), .DIN(N4967) );
hi1s1 U1616 ( .Q(N6227), .DIN(N4985) );
hi1s1 U1617 ( .Q(N6228), .DIN(N4988) );
hi1s1 U1618 ( .Q(N6229), .DIN(N4991) );
hi1s1 U1619 ( .Q(N6230), .DIN(N4994) );
hi1s1 U1620 ( .Q(N6231), .DIN(N5027) );
nb1s1 U1621 ( .Q(N6232), .DIN(N4711) );
hi1s1 U1622 ( .Q(N6235), .DIN(N5030) );
nb1s1 U1623 ( .Q(N6236), .DIN(N4735) );
hi1s1 U1624 ( .Q(N6239), .DIN(N5052) );
hi1s1 U1625 ( .Q(N6240), .DIN(N5055) );
hi1s1 U1626 ( .Q(N6241), .DIN(N5058) );
hi1s1 U1627 ( .Q(N6242), .DIN(N5061) );
nnd2s1 U1628 ( .Q(N6243), .DIN1(N5573), .DIN2(N5574) );
nnd2s1 U1629 ( .Q(N6246), .DIN1(N5571), .DIN2(N5572) );
nnd2s1 U1630 ( .Q(N6249), .DIN1(N5586), .DIN2(N5587) );
nnd2s1 U1631 ( .Q(N6252), .DIN1(N5584), .DIN2(N5585) );
hi1s1 U1632 ( .Q(N6255), .DIN(N5126) );
hi1s1 U1633 ( .Q(N6256), .DIN(N5129) );
hi1s1 U1634 ( .Q(N6257), .DIN(N5132) );
hi1s1 U1635 ( .Q(N6258), .DIN(N5135) );
hi1s1 U1636 ( .Q(N6259), .DIN(N5153) );
hi1s1 U1637 ( .Q(N6260), .DIN(N5156) );
hi1s1 U1638 ( .Q(N6261), .DIN(N5159) );
hi1s1 U1639 ( .Q(N6262), .DIN(N5162) );
nnd2s1 U1640 ( .Q(N6263), .DIN1(N5604), .DIN2(N5605) );
nnd2s1 U1641 ( .Q(N6266), .DIN1(N5602), .DIN2(N5603) );
nnd2s1 U1642 ( .Q(N6540), .DIN1(N1380), .DIN2(N5945) );
nnd2s1 U1643 ( .Q(N6541), .DIN1(N1383), .DIN2(N5947) );
nnd2s1 U1644 ( .Q(N6542), .DIN1(N1386), .DIN2(N5949) );
nnd2s1 U1645 ( .Q(N6543), .DIN1(N1389), .DIN2(N5951) );
nnd2s1 U1646 ( .Q(N6544), .DIN1(N1392), .DIN2(N5953) );
nnd2s1 U1647 ( .Q(N6545), .DIN1(N1395), .DIN2(N5955) );
nnd2s1 U1648 ( .Q(N6546), .DIN1(N1398), .DIN2(N5957) );
nnd2s1 U1649 ( .Q(N6547), .DIN1(N1401), .DIN2(N5959) );
nnd2s1 U1650 ( .Q(N6555), .DIN1(N1404), .DIN2(N5968) );
nnd2s1 U1651 ( .Q(N6556), .DIN1(N1407), .DIN2(N5970) );
nnd2s1 U1652 ( .Q(N6557), .DIN1(N1410), .DIN2(N5972) );
nnd2s1 U1653 ( .Q(N6558), .DIN1(N1413), .DIN2(N5974) );
nnd2s1 U1654 ( .Q(N6559), .DIN1(N1416), .DIN2(N5976) );
nnd2s1 U1655 ( .Q(N6560), .DIN1(N1419), .DIN2(N5978) );
nnd2s1 U1656 ( .Q(N6561), .DIN1(N1422), .DIN2(N5980) );
nnd2s1 U1657 ( .Q(N6569), .DIN1(N1425), .DIN2(N5990) );
nnd2s1 U1658 ( .Q(N6594), .DIN1(N3721), .DIN2(N6023) );
nnd2s1 U1659 ( .Q(N6595), .DIN1(N3724), .DIN2(N6025) );
nnd2s1 U1660 ( .Q(N6596), .DIN1(N3727), .DIN2(N6027) );
nnd2s1 U1661 ( .Q(N6597), .DIN1(N3730), .DIN2(N6029) );
nnd2s1 U1662 ( .Q(N6598), .DIN1(N4889), .DIN2(N6031) );
nnd2s1 U1663 ( .Q(N6599), .DIN1(N4886), .DIN2(N6032) );
nnd2s1 U1664 ( .Q(N6600), .DIN1(N4895), .DIN2(N6033) );
nnd2s1 U1665 ( .Q(N6601), .DIN1(N4892), .DIN2(N6034) );
nnd2s1 U1666 ( .Q(N6602), .DIN1(N4901), .DIN2(N6035) );
nnd2s1 U1667 ( .Q(N6603), .DIN1(N4898), .DIN2(N6036) );
nnd2s1 U1668 ( .Q(N6604), .DIN1(N3733), .DIN2(N6037) );
nnd2s1 U1669 ( .Q(N6605), .DIN1(N4910), .DIN2(N6039) );
nnd2s1 U1670 ( .Q(N6606), .DIN1(N4907), .DIN2(N6040) );
nnd2s1 U1671 ( .Q(N6621), .DIN1(N1434), .DIN2(N6061) );
nnd2s1 U1672 ( .Q(N6622), .DIN1(N1437), .DIN2(N6063) );
nnd2s1 U1673 ( .Q(N6623), .DIN1(N1440), .DIN2(N6065) );
nnd2s1 U1674 ( .Q(N6624), .DIN1(N1443), .DIN2(N6067) );
nnd2s1 U1675 ( .Q(N6625), .DIN1(N1446), .DIN2(N6069) );
nnd2s1 U1676 ( .Q(N6626), .DIN1(N1449), .DIN2(N6071) );
nnd2s1 U1677 ( .Q(N6627), .DIN1(N1452), .DIN2(N6073) );
nnd2s1 U1678 ( .Q(N6628), .DIN1(N1455), .DIN2(N6075) );
nnd2s1 U1679 ( .Q(N6629), .DIN1(N1458), .DIN2(N6077) );
nnd2s1 U1680 ( .Q(N6639), .DIN1(N3783), .DIN2(N6090) );
nnd2s1 U1681 ( .Q(N6640), .DIN1(N4949), .DIN2(N6092) );
nnd2s1 U1682 ( .Q(N6641), .DIN1(N4946), .DIN2(N6093) );
nnd2s1 U1683 ( .Q(N6642), .DIN1(N4955), .DIN2(N6094) );
nnd2s1 U1684 ( .Q(N6643), .DIN1(N4952), .DIN2(N6095) );
nnd2s1 U1685 ( .Q(N6644), .DIN1(N3786), .DIN2(N6096) );
nnd2s1 U1686 ( .Q(N6645), .DIN1(N4976), .DIN2(N6098) );
nnd2s1 U1687 ( .Q(N6646), .DIN1(N4973), .DIN2(N6099) );
nnd2s1 U1688 ( .Q(N6647), .DIN1(N4982), .DIN2(N6100) );
nnd2s1 U1689 ( .Q(N6648), .DIN1(N4979), .DIN2(N6101) );
nnd2s1 U1690 ( .Q(N6649), .DIN1(N1461), .DIN2(N6104) );
nnd2s1 U1691 ( .Q(N6650), .DIN1(N1464), .DIN2(N6106) );
nnd2s1 U1692 ( .Q(N6651), .DIN1(N1467), .DIN2(N6108) );
nnd2s1 U1693 ( .Q(N6652), .DIN1(N1470), .DIN2(N6110) );
nnd2s1 U1694 ( .Q(N6653), .DIN1(N1473), .DIN2(N6112) );
nnd2s1 U1695 ( .Q(N6654), .DIN1(N1476), .DIN2(N6114) );
nnd2s1 U1696 ( .Q(N6655), .DIN1(N1479), .DIN2(N6116) );
nnd2s1 U1697 ( .Q(N6656), .DIN1(N1482), .DIN2(N6118) );
nnd2s1 U1698 ( .Q(N6657), .DIN1(N1485), .DIN2(N6120) );
nnd2s1 U1699 ( .Q(N6658), .DIN1(N3789), .DIN2(N6121) );
nnd2s1 U1700 ( .Q(N6659), .DIN1(N5039), .DIN2(N6123) );
nnd2s1 U1701 ( .Q(N6660), .DIN1(N5036), .DIN2(N6124) );
nnd2s1 U1702 ( .Q(N6661), .DIN1(N3792), .DIN2(N6126) );
nnd2s1 U1703 ( .Q(N6668), .DIN1(N3816), .DIN2(N6135) );
nnd2s1 U1704 ( .Q(N6677), .DIN1(N5071), .DIN2(N6148) );
nnd2s1 U1705 ( .Q(N6678), .DIN1(N5068), .DIN2(N6149) );
nnd2s1 U1706 ( .Q(N6679), .DIN1(N5077), .DIN2(N6150) );
nnd2s1 U1707 ( .Q(N6680), .DIN1(N5074), .DIN2(N6151) );
nnd2s1 U1708 ( .Q(N6681), .DIN1(N5083), .DIN2(N6152) );
nnd2s1 U1709 ( .Q(N6682), .DIN1(N5080), .DIN2(N6153) );
nnd2s1 U1710 ( .Q(N6683), .DIN1(N5089), .DIN2(N6154) );
nnd2s1 U1711 ( .Q(N6684), .DIN1(N5086), .DIN2(N6155) );
nnd2s1 U1712 ( .Q(N6685), .DIN1(N3846), .DIN2(N6156) );
nnd2s1 U1713 ( .Q(N6686), .DIN1(N3849), .DIN2(N6158) );
nnd2s1 U1714 ( .Q(N6687), .DIN1(N3852), .DIN2(N6160) );
nnd2s1 U1715 ( .Q(N6688), .DIN1(N5104), .DIN2(N6162) );
nnd2s1 U1716 ( .Q(N6689), .DIN1(N5101), .DIN2(N6163) );
nnd2s1 U1717 ( .Q(N6690), .DIN1(N3855), .DIN2(N6165) );
nnd2s1 U1718 ( .Q(N6702), .DIN1(N5117), .DIN2(N6181) );
nnd2s1 U1719 ( .Q(N6703), .DIN1(N5114), .DIN2(N6182) );
nnd2s1 U1720 ( .Q(N6704), .DIN1(N5123), .DIN2(N6183) );
nnd2s1 U1721 ( .Q(N6705), .DIN1(N5120), .DIN2(N6184) );
nnd2s1 U1722 ( .Q(N6706), .DIN1(N3891), .DIN2(N6185) );
nnd2s1 U1723 ( .Q(N6707), .DIN1(N5144), .DIN2(N6187) );
nnd2s1 U1724 ( .Q(N6708), .DIN1(N5141), .DIN2(N6188) );
nnd2s1 U1725 ( .Q(N6709), .DIN1(N5150), .DIN2(N6189) );
nnd2s1 U1726 ( .Q(N6710), .DIN1(N5147), .DIN2(N6190) );
nnd2s1 U1727 ( .Q(N6711), .DIN1(N1708), .DIN2(N6191) );
nnd2s1 U1728 ( .Q(N6712), .DIN1(N2231), .DIN2(N6193) );
nnd2s1 U1729 ( .Q(N6729), .DIN1(N4961), .DIN2(N6223) );
nnd2s1 U1730 ( .Q(N6730), .DIN1(N4958), .DIN2(N6224) );
nnd2s1 U1731 ( .Q(N6731), .DIN1(N4967), .DIN2(N6225) );
nnd2s1 U1732 ( .Q(N6732), .DIN1(N4964), .DIN2(N6226) );
nnd2s1 U1733 ( .Q(N6733), .DIN1(N4988), .DIN2(N6227) );
nnd2s1 U1734 ( .Q(N6734), .DIN1(N4985), .DIN2(N6228) );
nnd2s1 U1735 ( .Q(N6735), .DIN1(N4994), .DIN2(N6229) );
nnd2s1 U1736 ( .Q(N6736), .DIN1(N4991), .DIN2(N6230) );
nnd2s1 U1737 ( .Q(N6741), .DIN1(N5055), .DIN2(N6239) );
nnd2s1 U1738 ( .Q(N6742), .DIN1(N5052), .DIN2(N6240) );
nnd2s1 U1739 ( .Q(N6743), .DIN1(N5061), .DIN2(N6241) );
nnd2s1 U1740 ( .Q(N6744), .DIN1(N5058), .DIN2(N6242) );
nnd2s1 U1741 ( .Q(N6751), .DIN1(N5129), .DIN2(N6255) );
nnd2s1 U1742 ( .Q(N6752), .DIN1(N5126), .DIN2(N6256) );
nnd2s1 U1743 ( .Q(N6753), .DIN1(N5135), .DIN2(N6257) );
nnd2s1 U1744 ( .Q(N6754), .DIN1(N5132), .DIN2(N6258) );
nnd2s1 U1745 ( .Q(N6755), .DIN1(N5156), .DIN2(N6259) );
nnd2s1 U1746 ( .Q(N6756), .DIN1(N5153), .DIN2(N6260) );
nnd2s1 U1747 ( .Q(N6757), .DIN1(N5162), .DIN2(N6261) );
nnd2s1 U1748 ( .Q(N6758), .DIN1(N5159), .DIN2(N6262) );
hi1s1 U1749 ( .Q(N6761), .DIN(N5892) );
and5s1 U1750 ( .Q(N6762), .DIN1(N5683), .DIN2(N5670), .DIN3(N5654), .DIN4(N5640), .DIN5(N5632) );
and2s1 U1751 ( .Q(N6766), .DIN1(N5632), .DIN2(N3097) );
and3s1 U1752 ( .Q(N6767), .DIN1(N5640), .DIN2(N5632), .DIN3(N3101) );
and4s1 U1753 ( .Q(N6768), .DIN1(N5654), .DIN2(N5632), .DIN3(N3107), .DIN4(N5640) );
and5s1 U1754 ( .Q(N6769), .DIN1(N5670), .DIN2(N5654), .DIN3(N5632), .DIN4(N3114), .DIN5(N5640) );
and2s1 U1755 ( .Q(N6770), .DIN1(N5640), .DIN2(N3101) );
and3s1 U1756 ( .Q(N6771), .DIN1(N5654), .DIN2(N3107), .DIN3(N5640) );
and4s1 U1757 ( .Q(N6772), .DIN1(N5670), .DIN2(N5654), .DIN3(N3114), .DIN4(N5640) );
and4s1 U1758 ( .Q(N6773), .DIN1(N5683), .DIN2(N5654), .DIN3(N5640), .DIN4(N5670) );
and2s1 U1759 ( .Q(N6774), .DIN1(N5640), .DIN2(N3101) );
and3s1 U1760 ( .Q(N6775), .DIN1(N5654), .DIN2(N3107), .DIN3(N5640) );
and4s1 U1761 ( .Q(N6776), .DIN1(N5670), .DIN2(N5654), .DIN3(N3114), .DIN4(N5640) );
and2s1 U1762 ( .Q(N6777), .DIN1(N5654), .DIN2(N3107) );
and3s1 U1763 ( .Q(N6778), .DIN1(N5670), .DIN2(N5654), .DIN3(N3114) );
and3s1 U1764 ( .Q(N6779), .DIN1(N5683), .DIN2(N5654), .DIN3(N5670) );
and2s1 U1765 ( .Q(N6780), .DIN1(N5654), .DIN2(N3107) );
and3s1 U1766 ( .Q(N6781), .DIN1(N5670), .DIN2(N5654), .DIN3(N3114) );
and2s1 U1767 ( .Q(N6782), .DIN1(N5670), .DIN2(N3114) );
and2s1 U1768 ( .Q(N6783), .DIN1(N5683), .DIN2(N5670) );
and5s1 U1769 ( .Q(N6784), .DIN1(N5697), .DIN2(N5728), .DIN3(N5707), .DIN4(N5690), .DIN5(N5718) );
and2s1 U1770 ( .Q(N6787), .DIN1(N5690), .DIN2(N3137) );
and3s1 U1771 ( .Q(N6788), .DIN1(N5697), .DIN2(N5690), .DIN3(N3140) );
and4s1 U1772 ( .Q(N6789), .DIN1(N5707), .DIN2(N5690), .DIN3(N3144), .DIN4(N5697) );
and5s1 U1773 ( .Q(N6790), .DIN1(N5718), .DIN2(N5707), .DIN3(N5690), .DIN4(N3149), .DIN5(N5697) );
and2s1 U1774 ( .Q(N6791), .DIN1(N5697), .DIN2(N3140) );
and3s1 U1775 ( .Q(N6792), .DIN1(N5707), .DIN2(N3144), .DIN3(N5697) );
and4s1 U1776 ( .Q(N6793), .DIN1(N5718), .DIN2(N5707), .DIN3(N3149), .DIN4(N5697) );
and2s1 U1777 ( .Q(N6794), .DIN1(N3144), .DIN2(N5707) );
and3s1 U1778 ( .Q(N6795), .DIN1(N5718), .DIN2(N5707), .DIN3(N3149) );
and2s1 U1779 ( .Q(N6796), .DIN1(N5718), .DIN2(N3149) );
hi1s1 U1780 ( .Q(N6797), .DIN(N5736) );
hi1s1 U1781 ( .Q(N6800), .DIN(N5740) );
hi1s1 U1782 ( .Q(N6803), .DIN(N5747) );
hi1s1 U1783 ( .Q(N6806), .DIN(N5751) );
hi1s1 U1784 ( .Q(N6809), .DIN(N5758) );
hi1s1 U1785 ( .Q(N6812), .DIN(N5762) );
nb1s1 U1786 ( .Q(N6815), .DIN(N5744) );
nb1s1 U1787 ( .Q(N6818), .DIN(N5744) );
nb1s1 U1788 ( .Q(N6821), .DIN(N5755) );
nb1s1 U1789 ( .Q(N6824), .DIN(N5755) );
nb1s1 U1790 ( .Q(N6827), .DIN(N5766) );
nb1s1 U1791 ( .Q(N6830), .DIN(N5766) );
and4s1 U1792 ( .Q(N6833), .DIN1(N5850), .DIN2(N5789), .DIN3(N5778), .DIN4(N5771) );
and2s1 U1793 ( .Q(N6836), .DIN1(N5771), .DIN2(N3169) );
and3s1 U1794 ( .Q(N6837), .DIN1(N5778), .DIN2(N5771), .DIN3(N3173) );
and4s1 U1795 ( .Q(N6838), .DIN1(N5789), .DIN2(N5771), .DIN3(N3178), .DIN4(N5778) );
and2s1 U1796 ( .Q(N6839), .DIN1(N5778), .DIN2(N3173) );
and3s1 U1797 ( .Q(N6840), .DIN1(N5789), .DIN2(N3178), .DIN3(N5778) );
and3s1 U1798 ( .Q(N6841), .DIN1(N5850), .DIN2(N5789), .DIN3(N5778) );
and2s1 U1799 ( .Q(N6842), .DIN1(N5778), .DIN2(N3173) );
and3s1 U1800 ( .Q(N6843), .DIN1(N5789), .DIN2(N3178), .DIN3(N5778) );
and2s1 U1801 ( .Q(N6844), .DIN1(N5789), .DIN2(N3178) );
and5s1 U1802 ( .Q(N6845), .DIN1(N5856), .DIN2(N5837), .DIN3(N5821), .DIN4(N5807), .DIN5(N5799) );
and2s1 U1803 ( .Q(N6848), .DIN1(N5799), .DIN2(N3185) );
and3s1 U1804 ( .Q(N6849), .DIN1(N5807), .DIN2(N5799), .DIN3(N3189) );
and4s1 U1805 ( .Q(N6850), .DIN1(N5821), .DIN2(N5799), .DIN3(N3195), .DIN4(N5807) );
and5s1 U1806 ( .Q(N6851), .DIN1(N5837), .DIN2(N5821), .DIN3(N5799), .DIN4(N3202), .DIN5(N5807) );
and2s1 U1807 ( .Q(N6852), .DIN1(N5807), .DIN2(N3189) );
and3s1 U1808 ( .Q(N6853), .DIN1(N5821), .DIN2(N3195), .DIN3(N5807) );
and4s1 U1809 ( .Q(N6854), .DIN1(N5837), .DIN2(N5821), .DIN3(N3202), .DIN4(N5807) );
and4s1 U1810 ( .Q(N6855), .DIN1(N5856), .DIN2(N5821), .DIN3(N5807), .DIN4(N5837) );
and2s1 U1811 ( .Q(N6856), .DIN1(N5807), .DIN2(N3189) );
and3s1 U1812 ( .Q(N6857), .DIN1(N5821), .DIN2(N3195), .DIN3(N5807) );
and4s1 U1813 ( .Q(N6858), .DIN1(N5837), .DIN2(N5821), .DIN3(N3202), .DIN4(N5807) );
and2s1 U1814 ( .Q(N6859), .DIN1(N5821), .DIN2(N3195) );
and3s1 U1815 ( .Q(N6860), .DIN1(N5837), .DIN2(N5821), .DIN3(N3202) );
and3s1 U1816 ( .Q(N6861), .DIN1(N5856), .DIN2(N5821), .DIN3(N5837) );
and2s1 U1817 ( .Q(N6862), .DIN1(N5821), .DIN2(N3195) );
and3s1 U1818 ( .Q(N6863), .DIN1(N5837), .DIN2(N5821), .DIN3(N3202) );
and2s1 U1819 ( .Q(N6864), .DIN1(N5837), .DIN2(N3202) );
and2s1 U1820 ( .Q(N6865), .DIN1(N5850), .DIN2(N5789) );
and2s1 U1821 ( .Q(N6866), .DIN1(N5856), .DIN2(N5837) );
and4s1 U1822 ( .Q(N6867), .DIN1(N5870), .DIN2(N5892), .DIN3(N5881), .DIN4(N5863) );
and2s1 U1823 ( .Q(N6870), .DIN1(N5863), .DIN2(N3211) );
and3s1 U1824 ( .Q(N6871), .DIN1(N5870), .DIN2(N5863), .DIN3(N3215) );
and4s1 U1825 ( .Q(N6872), .DIN1(N5881), .DIN2(N5863), .DIN3(N3221), .DIN4(N5870) );
and2s1 U1826 ( .Q(N6873), .DIN1(N5870), .DIN2(N3215) );
and3s1 U1827 ( .Q(N6874), .DIN1(N5881), .DIN2(N3221), .DIN3(N5870) );
and3s1 U1828 ( .Q(N6875), .DIN1(N5892), .DIN2(N5881), .DIN3(N5870) );
and2s1 U1829 ( .Q(N6876), .DIN1(N5870), .DIN2(N3215) );
and3s1 U1830 ( .Q(N6877), .DIN1(N3221), .DIN2(N5881), .DIN3(N5870) );
and2s1 U1831 ( .Q(N6878), .DIN1(N5881), .DIN2(N3221) );
and2s1 U1832 ( .Q(N6879), .DIN1(N5892), .DIN2(N5881) );
and2s1 U1833 ( .Q(N6880), .DIN1(N5881), .DIN2(N3221) );
and5s1 U1834 ( .Q(N6881), .DIN1(N5905), .DIN2(N5936), .DIN3(N5915), .DIN4(N5898), .DIN5(N5926) );
and2s1 U1835 ( .Q(N6884), .DIN1(N5898), .DIN2(N3229) );
and3s1 U1836 ( .Q(N6885), .DIN1(N5905), .DIN2(N5898), .DIN3(N3232) );
and4s1 U1837 ( .Q(N6886), .DIN1(N5915), .DIN2(N5898), .DIN3(N3236), .DIN4(N5905) );
and5s1 U1838 ( .Q(N6887), .DIN1(N5926), .DIN2(N5915), .DIN3(N5898), .DIN4(N3241), .DIN5(N5905) );
and2s1 U1839 ( .Q(N6888), .DIN1(N5905), .DIN2(N3232) );
and3s1 U1840 ( .Q(N6889), .DIN1(N5915), .DIN2(N3236), .DIN3(N5905) );
and4s1 U1841 ( .Q(N6890), .DIN1(N5926), .DIN2(N5915), .DIN3(N3241), .DIN4(N5905) );
and2s1 U1842 ( .Q(N6891), .DIN1(N3236), .DIN2(N5915) );
and3s1 U1843 ( .Q(N6892), .DIN1(N5926), .DIN2(N5915), .DIN3(N3241) );
and2s1 U1844 ( .Q(N6893), .DIN1(N5926), .DIN2(N3241) );
nnd2s1 U1845 ( .Q(N6894), .DIN1(N5944), .DIN2(N6540) );
nnd2s1 U1846 ( .Q(N6901), .DIN1(N5946), .DIN2(N6541) );
nnd2s1 U1847 ( .Q(N6912), .DIN1(N5948), .DIN2(N6542) );
nnd2s1 U1848 ( .Q(N6923), .DIN1(N5950), .DIN2(N6543) );
nnd2s1 U1849 ( .Q(N6929), .DIN1(N5952), .DIN2(N6544) );
nnd2s1 U1850 ( .Q(N6936), .DIN1(N5954), .DIN2(N6545) );
nnd2s1 U1851 ( .Q(N6946), .DIN1(N5956), .DIN2(N6546) );
nnd2s1 U1852 ( .Q(N6957), .DIN1(N5958), .DIN2(N6547) );
nnd2s1 U1853 ( .Q(N6967), .DIN1(N6204), .DIN2(N4575) );
hi1s1 U1854 ( .Q(N6968), .DIN(N6204) );
hi1s1 U1855 ( .Q(N6969), .DIN(N6207) );
nnd2s1 U1856 ( .Q(N6970), .DIN1(N5967), .DIN2(N6555) );
nnd2s1 U1857 ( .Q(N6977), .DIN1(N5969), .DIN2(N6556) );
nnd2s1 U1858 ( .Q(N6988), .DIN1(N5971), .DIN2(N6557) );
nnd2s1 U1859 ( .Q(N6998), .DIN1(N5973), .DIN2(N6558) );
nnd2s1 U1860 ( .Q(N7006), .DIN1(N5975), .DIN2(N6559) );
nnd2s1 U1861 ( .Q(N7020), .DIN1(N5977), .DIN2(N6560) );
nnd2s1 U1862 ( .Q(N7036), .DIN1(N5979), .DIN2(N6561) );
nnd2s1 U1863 ( .Q(N7049), .DIN1(N5989), .DIN2(N6569) );
nnd2s1 U1864 ( .Q(N7055), .DIN1(N6210), .DIN2(N4610) );
hi1s1 U1865 ( .Q(N7056), .DIN(N6210) );
and4s1 U1866 ( .Q(N7057), .DIN1(N6021), .DIN2(N6000), .DIN3(N5996), .DIN4(N5991) );
and2s1 U1867 ( .Q(N7060), .DIN1(N5991), .DIN2(N3362) );
and3s1 U1868 ( .Q(N7061), .DIN1(N5996), .DIN2(N5991), .DIN3(N3363) );
and4s1 U1869 ( .Q(N7062), .DIN1(N6000), .DIN2(N5991), .DIN3(N3364), .DIN4(N5996) );
and5s1 U1870 ( .Q(N7063), .DIN1(N6022), .DIN2(N6018), .DIN3(N6014), .DIN4(N6009), .DIN5(N6003) );
and2s1 U1871 ( .Q(N7064), .DIN1(N6003), .DIN2(N3366) );
and3s1 U1872 ( .Q(N7065), .DIN1(N6009), .DIN2(N6003), .DIN3(N3367) );
and4s1 U1873 ( .Q(N7066), .DIN1(N6014), .DIN2(N6003), .DIN3(N3368), .DIN4(N6009) );
and5s1 U1874 ( .Q(N7067), .DIN1(N6018), .DIN2(N6014), .DIN3(N6003), .DIN4(N3369), .DIN5(N6009) );
nnd2s1 U1875 ( .Q(N7068), .DIN1(N6594), .DIN2(N6024) );
nnd2s1 U1876 ( .Q(N7073), .DIN1(N6595), .DIN2(N6026) );
nnd2s1 U1877 ( .Q(N7077), .DIN1(N6596), .DIN2(N6028) );
nnd2s1 U1878 ( .Q(N7080), .DIN1(N6597), .DIN2(N6030) );
nnd2s1 U1879 ( .Q(N7086), .DIN1(N6598), .DIN2(N6599) );
nnd2s1 U1880 ( .Q(N7091), .DIN1(N6600), .DIN2(N6601) );
nnd2s1 U1881 ( .Q(N7095), .DIN1(N6602), .DIN2(N6603) );
nnd2s1 U1882 ( .Q(N7098), .DIN1(N6604), .DIN2(N6038) );
nnd2s1 U1883 ( .Q(N7099), .DIN1(N6605), .DIN2(N6606) );
and5s1 U1884 ( .Q(N7100), .DIN1(N6059), .DIN2(N6056), .DIN3(N6052), .DIN4(N6047), .DIN5(N6041) );
and2s1 U1885 ( .Q(N7103), .DIN1(N6041), .DIN2(N3371) );
and3s1 U1886 ( .Q(N7104), .DIN1(N6047), .DIN2(N6041), .DIN3(N3372) );
and4s1 U1887 ( .Q(N7105), .DIN1(N6052), .DIN2(N6041), .DIN3(N3373), .DIN4(N6047) );
and5s1 U1888 ( .Q(N7106), .DIN1(N6056), .DIN2(N6052), .DIN3(N6041), .DIN4(N3374), .DIN5(N6047) );
nnd2s1 U1889 ( .Q(N7107), .DIN1(N6060), .DIN2(N6621) );
nnd2s1 U1890 ( .Q(N7114), .DIN1(N6062), .DIN2(N6622) );
nnd2s1 U1891 ( .Q(N7125), .DIN1(N6064), .DIN2(N6623) );
nnd2s1 U1892 ( .Q(N7136), .DIN1(N6066), .DIN2(N6624) );
nnd2s1 U1893 ( .Q(N7142), .DIN1(N6068), .DIN2(N6625) );
nnd2s1 U1894 ( .Q(N7149), .DIN1(N6070), .DIN2(N6626) );
nnd2s1 U1895 ( .Q(N7159), .DIN1(N6072), .DIN2(N6627) );
nnd2s1 U1896 ( .Q(N7170), .DIN1(N6074), .DIN2(N6628) );
nnd2s1 U1897 ( .Q(N7180), .DIN1(N6076), .DIN2(N6629) );
hi1s1 U1898 ( .Q(N7187), .DIN(N6220) );
hi1s1 U1899 ( .Q(N7188), .DIN(N6079) );
hi1s1 U1900 ( .Q(N7191), .DIN(N6083) );
nnd2s1 U1901 ( .Q(N7194), .DIN1(N6639), .DIN2(N6091) );
nnd2s1 U1902 ( .Q(N7198), .DIN1(N6640), .DIN2(N6641) );
nnd2s1 U1903 ( .Q(N7202), .DIN1(N6642), .DIN2(N6643) );
nnd2s1 U1904 ( .Q(N7205), .DIN1(N6644), .DIN2(N6097) );
nnd2s1 U1905 ( .Q(N7209), .DIN1(N6645), .DIN2(N6646) );
nnd2s1 U1906 ( .Q(N7213), .DIN1(N6647), .DIN2(N6648) );
nb1s1 U1907 ( .Q(N7216), .DIN(N6087) );
nb1s1 U1908 ( .Q(N7219), .DIN(N6087) );
nnd2s1 U1909 ( .Q(N7222), .DIN1(N6103), .DIN2(N6649) );
nnd2s1 U1910 ( .Q(N7229), .DIN1(N6105), .DIN2(N6650) );
nnd2s1 U1911 ( .Q(N7240), .DIN1(N6107), .DIN2(N6651) );
nnd2s1 U1912 ( .Q(N7250), .DIN1(N6109), .DIN2(N6652) );
nnd2s1 U1913 ( .Q(N7258), .DIN1(N6111), .DIN2(N6653) );
nnd2s1 U1914 ( .Q(N7272), .DIN1(N6113), .DIN2(N6654) );
nnd2s1 U1915 ( .Q(N7288), .DIN1(N6115), .DIN2(N6655) );
nnd2s1 U1916 ( .Q(N7301), .DIN1(N6117), .DIN2(N6656) );
nnd2s1 U1917 ( .Q(N7307), .DIN1(N6119), .DIN2(N6657) );
nnd2s1 U1918 ( .Q(N7314), .DIN1(N6658), .DIN2(N6122) );
nnd2s1 U1919 ( .Q(N7318), .DIN1(N6659), .DIN2(N6660) );
nnd2s1 U1920 ( .Q(N7322), .DIN1(N6125), .DIN2(N6661) );
hi1s1 U1921 ( .Q(N7325), .DIN(N6127) );
hi1s1 U1922 ( .Q(N7328), .DIN(N6131) );
nnd2s1 U1923 ( .Q(N7331), .DIN1(N6668), .DIN2(N6136) );
hi1s1 U1924 ( .Q(N7334), .DIN(N6137) );
hi1s1 U1925 ( .Q(N7337), .DIN(N6141) );
nb1s1 U1926 ( .Q(N7340), .DIN(N6145) );
nb1s1 U1927 ( .Q(N7343), .DIN(N6145) );
nnd2s1 U1928 ( .Q(N7346), .DIN1(N6677), .DIN2(N6678) );
nnd2s1 U1929 ( .Q(N7351), .DIN1(N6679), .DIN2(N6680) );
nnd2s1 U1930 ( .Q(N7355), .DIN1(N6681), .DIN2(N6682) );
nnd2s1 U1931 ( .Q(N7358), .DIN1(N6683), .DIN2(N6684) );
nnd2s1 U1932 ( .Q(N7364), .DIN1(N6685), .DIN2(N6157) );
nnd2s1 U1933 ( .Q(N7369), .DIN1(N6686), .DIN2(N6159) );
nnd2s1 U1934 ( .Q(N7373), .DIN1(N6687), .DIN2(N6161) );
nnd2s1 U1935 ( .Q(N7376), .DIN1(N6688), .DIN2(N6689) );
nnd2s1 U1936 ( .Q(N7377), .DIN1(N6164), .DIN2(N6690) );
hi1s1 U1937 ( .Q(N7378), .DIN(N6166) );
hi1s1 U1938 ( .Q(N7381), .DIN(N6170) );
hi1s1 U1939 ( .Q(N7384), .DIN(N6177) );
nnd2s1 U1940 ( .Q(N7387), .DIN1(N6702), .DIN2(N6703) );
nnd2s1 U1941 ( .Q(N7391), .DIN1(N6704), .DIN2(N6705) );
nnd2s1 U1942 ( .Q(N7394), .DIN1(N6706), .DIN2(N6186) );
nnd2s1 U1943 ( .Q(N7398), .DIN1(N6707), .DIN2(N6708) );
nnd2s1 U1944 ( .Q(N7402), .DIN1(N6709), .DIN2(N6710) );
nb1s1 U1945 ( .Q(N7405), .DIN(N6174) );
nb1s1 U1946 ( .Q(N7408), .DIN(N6174) );
nb1s1 U1947 ( .Q(N7411), .DIN(N5936) );
nb1s1 U1948 ( .Q(N7414), .DIN(N5898) );
nb1s1 U1949 ( .Q(N7417), .DIN(N5905) );
nb1s1 U1950 ( .Q(N7420), .DIN(N5915) );
nb1s1 U1951 ( .Q(N7423), .DIN(N5926) );
nb1s1 U1952 ( .Q(N7426), .DIN(N5728) );
nb1s1 U1953 ( .Q(N7429), .DIN(N5690) );
nb1s1 U1954 ( .Q(N7432), .DIN(N5697) );
nb1s1 U1955 ( .Q(N7435), .DIN(N5707) );
nb1s1 U1956 ( .Q(N7438), .DIN(N5718) );
nnd2s1 U1957 ( .Q(N7441), .DIN1(N6192), .DIN2(N6711) );
nnd2s1 U1958 ( .Q(N7444), .DIN1(N6194), .DIN2(N6712) );
nb1s1 U1959 ( .Q(N7447), .DIN(N5683) );
nb1s1 U1960 ( .Q(N7450), .DIN(N5670) );
nb1s1 U1961 ( .Q(N7453), .DIN(N5632) );
nb1s1 U1962 ( .Q(N7456), .DIN(N5654) );
nb1s1 U1963 ( .Q(N7459), .DIN(N5640) );
nb1s1 U1964 ( .Q(N7462), .DIN(N5640) );
nb1s1 U1965 ( .Q(N7465), .DIN(N5683) );
nb1s1 U1966 ( .Q(N7468), .DIN(N5670) );
nb1s1 U1967 ( .Q(N7471), .DIN(N5632) );
nb1s1 U1968 ( .Q(N7474), .DIN(N5654) );
hi1s1 U1969 ( .Q(N7477), .DIN(N6196) );
hi1s1 U1970 ( .Q(N7478), .DIN(N6199) );
nb1s1 U1971 ( .Q(N7479), .DIN(N5850) );
nb1s1 U1972 ( .Q(N7482), .DIN(N5789) );
nb1s1 U1973 ( .Q(N7485), .DIN(N5771) );
nb1s1 U1974 ( .Q(N7488), .DIN(N5778) );
nb1s1 U1975 ( .Q(N7491), .DIN(N5850) );
nb1s1 U1976 ( .Q(N7494), .DIN(N5789) );
nb1s1 U1977 ( .Q(N7497), .DIN(N5771) );
nb1s1 U1978 ( .Q(N7500), .DIN(N5778) );
nb1s1 U1979 ( .Q(N7503), .DIN(N5856) );
nb1s1 U1980 ( .Q(N7506), .DIN(N5837) );
nb1s1 U1981 ( .Q(N7509), .DIN(N5799) );
nb1s1 U1982 ( .Q(N7512), .DIN(N5821) );
nb1s1 U1983 ( .Q(N7515), .DIN(N5807) );
nb1s1 U1984 ( .Q(N7518), .DIN(N5807) );
nb1s1 U1985 ( .Q(N7521), .DIN(N5856) );
nb1s1 U1986 ( .Q(N7524), .DIN(N5837) );
nb1s1 U1987 ( .Q(N7527), .DIN(N5799) );
nb1s1 U1988 ( .Q(N7530), .DIN(N5821) );
nb1s1 U1989 ( .Q(N7533), .DIN(N5863) );
nb1s1 U1990 ( .Q(N7536), .DIN(N5863) );
nb1s1 U1991 ( .Q(N7539), .DIN(N5870) );
nb1s1 U1992 ( .Q(N7542), .DIN(N5870) );
nb1s1 U1993 ( .Q(N7545), .DIN(N5881) );
nb1s1 U1994 ( .Q(N7548), .DIN(N5881) );
hi1s1 U1995 ( .Q(N7551), .DIN(N6214) );
hi1s1 U1996 ( .Q(N7552), .DIN(N6217) );
nb1s1 U1997 ( .Q(N7553), .DIN(N5981) );
hi1s1 U1998 ( .Q(N7556), .DIN(N6249) );
hi1s1 U1999 ( .Q(N7557), .DIN(N6252) );
hi1s1 U2000 ( .Q(N7558), .DIN(N6243) );
hi1s1 U2001 ( .Q(N7559), .DIN(N6246) );
nnd2s1 U2002 ( .Q(N7560), .DIN1(N6731), .DIN2(N6732) );
nnd2s1 U2003 ( .Q(N7563), .DIN1(N6729), .DIN2(N6730) );
nnd2s1 U2004 ( .Q(N7566), .DIN1(N6735), .DIN2(N6736) );
nnd2s1 U2005 ( .Q(N7569), .DIN1(N6733), .DIN2(N6734) );
hi1s1 U2006 ( .Q(N7572), .DIN(N6232) );
hi1s1 U2007 ( .Q(N7573), .DIN(N6236) );
nnd2s1 U2008 ( .Q(N7574), .DIN1(N6743), .DIN2(N6744) );
nnd2s1 U2009 ( .Q(N7577), .DIN1(N6741), .DIN2(N6742) );
hi1s1 U2010 ( .Q(N7580), .DIN(N6263) );
hi1s1 U2011 ( .Q(N7581), .DIN(N6266) );
nnd2s1 U2012 ( .Q(N7582), .DIN1(N6753), .DIN2(N6754) );
nnd2s1 U2013 ( .Q(N7585), .DIN1(N6751), .DIN2(N6752) );
nnd2s1 U2014 ( .Q(N7588), .DIN1(N6757), .DIN2(N6758) );
nnd2s1 U2015 ( .Q(N7591), .DIN1(N6755), .DIN2(N6756) );
or5s1 U2016 ( .Q(N7609), .DIN1(N3096), .DIN2(N6766), .DIN3(N6767), .DIN4(N6768), .DIN5(N6769) );
or2s1 U2017 ( .Q(N7613), .DIN1(N3107), .DIN2(N6782) );
or5s1 U2018 ( .Q(N7620), .DIN1(N3136), .DIN2(N6787), .DIN3(N6788), .DIN4(N6789), .DIN5(N6790) );
or4s1 U2019 ( .Q(N7649), .DIN1(N3168), .DIN2(N6836), .DIN3(N6837), .DIN4(N6838) );
or2s1 U2020 ( .Q(N7650), .DIN1(N3173), .DIN2(N6844) );
or5s1 U2021 ( .Q(N7655), .DIN1(N3184), .DIN2(N6848), .DIN3(N6849), .DIN4(N6850), .DIN5(N6851) );
or2s1 U2022 ( .Q(N7659), .DIN1(N3195), .DIN2(N6864) );
or4s1 U2023 ( .Q(N7668), .DIN1(N3210), .DIN2(N6870), .DIN3(N6871), .DIN4(N6872) );
or5s1 U2024 ( .Q(N7671), .DIN1(N3228), .DIN2(N6884), .DIN3(N6885), .DIN4(N6886), .DIN5(N6887) );
nnd2s1 U2025 ( .Q(N7744), .DIN1(N3661), .DIN2(N6968) );
nnd2s1 U2026 ( .Q(N7822), .DIN1(N3664), .DIN2(N7056) );
or4s1 U2027 ( .Q(N7825), .DIN1(N3361), .DIN2(N7060), .DIN3(N7061), .DIN4(N7062) );
or5s1 U2028 ( .Q(N7826), .DIN1(N3365), .DIN2(N7064), .DIN3(N7065), .DIN4(N7066), .DIN5(N7067) );
or5s1 U2029 ( .Q(N7852), .DIN1(N3370), .DIN2(N7103), .DIN3(N7104), .DIN4(N7105), .DIN5(N7106) );
or4s1 U2030 ( .Q(N8114), .DIN1(N3101), .DIN2(N6777), .DIN3(N6778), .DIN4(N6779) );
or5s1 U2031 ( .Q(N8117), .DIN1(N3097), .DIN2(N6770), .DIN3(N6771), .DIN4(N6772), .DIN5(N6773) );
nor3s1 U2032 ( .Q(N8131), .DIN1(N3101), .DIN2(N6780), .DIN3(N6781) );
nor4s1 U2033 ( .Q(N8134), .DIN1(N3097), .DIN2(N6774), .DIN3(N6775), .DIN4(N6776) );
nnd2s1 U2034 ( .Q(N8144), .DIN1(N6199), .DIN2(N7477) );
nnd2s1 U2035 ( .Q(N8145), .DIN1(N6196), .DIN2(N7478) );
or4s1 U2036 ( .Q(N8146), .DIN1(N3169), .DIN2(N6839), .DIN3(N6840), .DIN4(N6841) );
nor3s1 U2037 ( .Q(N8156), .DIN1(N3169), .DIN2(N6842), .DIN3(N6843) );
or4s1 U2038 ( .Q(N8166), .DIN1(N3189), .DIN2(N6859), .DIN3(N6860), .DIN4(N6861) );
or5s1 U2039 ( .Q(N8169), .DIN1(N3185), .DIN2(N6852), .DIN3(N6853), .DIN4(N6854), .DIN5(N6855) );
nor3s1 U2040 ( .Q(N8183), .DIN1(N3189), .DIN2(N6862), .DIN3(N6863) );
nor4s1 U2041 ( .Q(N8186), .DIN1(N3185), .DIN2(N6856), .DIN3(N6857), .DIN4(N6858) );
or4s1 U2042 ( .Q(N8196), .DIN1(N3211), .DIN2(N6873), .DIN3(N6874), .DIN4(N6875) );
nor3s1 U2043 ( .Q(N8200), .DIN1(N3211), .DIN2(N6876), .DIN3(N6877) );
or3s1 U2044 ( .Q(N8204), .DIN1(N3215), .DIN2(N6878), .DIN3(N6879) );
nor2s1 U2045 ( .Q(N8208), .DIN1(N3215), .DIN2(N6880) );
nnd2s1 U2046 ( .Q(N8216), .DIN1(N6252), .DIN2(N7556) );
nnd2s1 U2047 ( .Q(N8217), .DIN1(N6249), .DIN2(N7557) );
nnd2s1 U2048 ( .Q(N8218), .DIN1(N6246), .DIN2(N7558) );
nnd2s1 U2049 ( .Q(N8219), .DIN1(N6243), .DIN2(N7559) );
nnd2s1 U2050 ( .Q(N8232), .DIN1(N6266), .DIN2(N7580) );
nnd2s1 U2051 ( .Q(N8233), .DIN1(N6263), .DIN2(N7581) );
hi1s1 U2052 ( .Q(N8242), .DIN(N7411) );
hi1s1 U2053 ( .Q(N8243), .DIN(N7414) );
hi1s1 U2054 ( .Q(N8244), .DIN(N7417) );
hi1s1 U2055 ( .Q(N8245), .DIN(N7420) );
hi1s1 U2056 ( .Q(N8246), .DIN(N7423) );
hi1s1 U2057 ( .Q(N8247), .DIN(N7426) );
hi1s1 U2058 ( .Q(N8248), .DIN(N7429) );
hi1s1 U2059 ( .Q(N8249), .DIN(N7432) );
hi1s1 U2060 ( .Q(N8250), .DIN(N7435) );
hi1s1 U2061 ( .Q(N8251), .DIN(N7438) );
hi1s1 U2062 ( .Q(N8252), .DIN(N7136) );
hi1s1 U2063 ( .Q(N8253), .DIN(N6923) );
hi1s1 U2064 ( .Q(N8254), .DIN(N6762) );
hi1s1 U2065 ( .Q(N8260), .DIN(N7459) );
hi1s1 U2066 ( .Q(N8261), .DIN(N7462) );
and2s1 U2067 ( .Q(N8262), .DIN1(N3122), .DIN2(N6762) );
and2s1 U2068 ( .Q(N8269), .DIN1(N3155), .DIN2(N6784) );
hi1s1 U2069 ( .Q(N8274), .DIN(N6815) );
hi1s1 U2070 ( .Q(N8275), .DIN(N6818) );
hi1s1 U2071 ( .Q(N8276), .DIN(N6821) );
hi1s1 U2072 ( .Q(N8277), .DIN(N6824) );
hi1s1 U2073 ( .Q(N8278), .DIN(N6827) );
hi1s1 U2074 ( .Q(N8279), .DIN(N6830) );
and3s1 U2075 ( .Q(N8280), .DIN1(N5740), .DIN2(N5736), .DIN3(N6815) );
and3s1 U2076 ( .Q(N8281), .DIN1(N6800), .DIN2(N6797), .DIN3(N6818) );
and3s1 U2077 ( .Q(N8282), .DIN1(N5751), .DIN2(N5747), .DIN3(N6821) );
and3s1 U2078 ( .Q(N8283), .DIN1(N6806), .DIN2(N6803), .DIN3(N6824) );
and3s1 U2079 ( .Q(N8284), .DIN1(N5762), .DIN2(N5758), .DIN3(N6827) );
and3s1 U2080 ( .Q(N8285), .DIN1(N6812), .DIN2(N6809), .DIN3(N6830) );
hi1s1 U2081 ( .Q(N8288), .DIN(N6845) );
hi1s1 U2082 ( .Q(N8294), .DIN(N7488) );
hi1s1 U2083 ( .Q(N8295), .DIN(N7500) );
hi1s1 U2084 ( .Q(N8296), .DIN(N7515) );
hi1s1 U2085 ( .Q(N8297), .DIN(N7518) );
and2s1 U2086 ( .Q(N8298), .DIN1(N6833), .DIN2(N6845) );
and2s1 U2087 ( .Q(N8307), .DIN1(N6867), .DIN2(N6881) );
hi1s1 U2088 ( .Q(N8315), .DIN(N7533) );
hi1s1 U2089 ( .Q(N8317), .DIN(N7536) );
hi1s1 U2090 ( .Q(N8319), .DIN(N7539) );
hi1s1 U2091 ( .Q(N8321), .DIN(N7542) );
nnd2s1 U2092 ( .Q(N8322), .DIN1(N7545), .DIN2(N4543) );
hi1s1 U2093 ( .Q(N8323), .DIN(N7545) );
nnd2s1 U2094 ( .Q(N8324), .DIN1(N7548), .DIN2(N5943) );
hi1s1 U2095 ( .Q(N8325), .DIN(N7548) );
nnd2s1 U2096 ( .Q(N8326), .DIN1(N6967), .DIN2(N7744) );
and4s1 U2097 ( .Q(N8333), .DIN1(N6901), .DIN2(N6923), .DIN3(N6912), .DIN4(N6894) );
and2s1 U2098 ( .Q(N8337), .DIN1(N6894), .DIN2(N4545) );
and3s1 U2099 ( .Q(N8338), .DIN1(N6901), .DIN2(N6894), .DIN3(N4549) );
and4s1 U2100 ( .Q(N8339), .DIN1(N6912), .DIN2(N6894), .DIN3(N4555), .DIN4(N6901) );
and2s1 U2101 ( .Q(N8340), .DIN1(N6901), .DIN2(N4549) );
and3s1 U2102 ( .Q(N8341), .DIN1(N6912), .DIN2(N4555), .DIN3(N6901) );
and3s1 U2103 ( .Q(N8342), .DIN1(N6923), .DIN2(N6912), .DIN3(N6901) );
and2s1 U2104 ( .Q(N8343), .DIN1(N6901), .DIN2(N4549) );
and3s1 U2105 ( .Q(N8344), .DIN1(N4555), .DIN2(N6912), .DIN3(N6901) );
and2s1 U2106 ( .Q(N8345), .DIN1(N6912), .DIN2(N4555) );
and2s1 U2107 ( .Q(N8346), .DIN1(N6923), .DIN2(N6912) );
and2s1 U2108 ( .Q(N8347), .DIN1(N6912), .DIN2(N4555) );
and2s1 U2109 ( .Q(N8348), .DIN1(N6929), .DIN2(N4563) );
and3s1 U2110 ( .Q(N8349), .DIN1(N6936), .DIN2(N6929), .DIN3(N4566) );
and4s1 U2111 ( .Q(N8350), .DIN1(N6946), .DIN2(N6929), .DIN3(N4570), .DIN4(N6936) );
and5s1 U2112 ( .Q(N8351), .DIN1(N6957), .DIN2(N6946), .DIN3(N6929), .DIN4(N5960), .DIN5(N6936) );
and2s1 U2113 ( .Q(N8352), .DIN1(N6936), .DIN2(N4566) );
and3s1 U2114 ( .Q(N8353), .DIN1(N6946), .DIN2(N4570), .DIN3(N6936) );
and4s1 U2115 ( .Q(N8354), .DIN1(N6957), .DIN2(N6946), .DIN3(N5960), .DIN4(N6936) );
and2s1 U2116 ( .Q(N8355), .DIN1(N4570), .DIN2(N6946) );
and3s1 U2117 ( .Q(N8356), .DIN1(N6957), .DIN2(N6946), .DIN3(N5960) );
and2s1 U2118 ( .Q(N8357), .DIN1(N6957), .DIN2(N5960) );
nnd2s1 U2119 ( .Q(N8358), .DIN1(N7055), .DIN2(N7822) );
and4s1 U2120 ( .Q(N8365), .DIN1(N7049), .DIN2(N6988), .DIN3(N6977), .DIN4(N6970) );
and2s1 U2121 ( .Q(N8369), .DIN1(N6970), .DIN2(N4577) );
and3s1 U2122 ( .Q(N8370), .DIN1(N6977), .DIN2(N6970), .DIN3(N4581) );
and4s1 U2123 ( .Q(N8371), .DIN1(N6988), .DIN2(N6970), .DIN3(N4586), .DIN4(N6977) );
and2s1 U2124 ( .Q(N8372), .DIN1(N6977), .DIN2(N4581) );
and3s1 U2125 ( .Q(N8373), .DIN1(N6988), .DIN2(N4586), .DIN3(N6977) );
and3s1 U2126 ( .Q(N8374), .DIN1(N7049), .DIN2(N6988), .DIN3(N6977) );
and2s1 U2127 ( .Q(N8375), .DIN1(N6977), .DIN2(N4581) );
and3s1 U2128 ( .Q(N8376), .DIN1(N6988), .DIN2(N4586), .DIN3(N6977) );
and2s1 U2129 ( .Q(N8377), .DIN1(N6988), .DIN2(N4586) );
and2s1 U2130 ( .Q(N8378), .DIN1(N6998), .DIN2(N4593) );
and3s1 U2131 ( .Q(N8379), .DIN1(N7006), .DIN2(N6998), .DIN3(N4597) );
and4s1 U2132 ( .Q(N8380), .DIN1(N7020), .DIN2(N6998), .DIN3(N4603), .DIN4(N7006) );
and5s1 U2133 ( .Q(N8381), .DIN1(N7036), .DIN2(N7020), .DIN3(N6998), .DIN4(N5981), .DIN5(N7006) );
and2s1 U2134 ( .Q(N8382), .DIN1(N7006), .DIN2(N4597) );
and3s1 U2135 ( .Q(N8383), .DIN1(N7020), .DIN2(N4603), .DIN3(N7006) );
and4s1 U2136 ( .Q(N8384), .DIN1(N7036), .DIN2(N7020), .DIN3(N5981), .DIN4(N7006) );
and2s1 U2137 ( .Q(N8385), .DIN1(N7006), .DIN2(N4597) );
and3s1 U2138 ( .Q(N8386), .DIN1(N7020), .DIN2(N4603), .DIN3(N7006) );
and4s1 U2139 ( .Q(N8387), .DIN1(N7036), .DIN2(N7020), .DIN3(N5981), .DIN4(N7006) );
and2s1 U2140 ( .Q(N8388), .DIN1(N7020), .DIN2(N4603) );
and3s1 U2141 ( .Q(N8389), .DIN1(N7036), .DIN2(N7020), .DIN3(N5981) );
and2s1 U2142 ( .Q(N8390), .DIN1(N7020), .DIN2(N4603) );
and3s1 U2143 ( .Q(N8391), .DIN1(N7036), .DIN2(N7020), .DIN3(N5981) );
and2s1 U2144 ( .Q(N8392), .DIN1(N7036), .DIN2(N5981) );
and2s1 U2145 ( .Q(N8393), .DIN1(N7049), .DIN2(N6988) );
and2s1 U2146 ( .Q(N8394), .DIN1(N7057), .DIN2(N7063) );
and2s1 U2147 ( .Q(N8404), .DIN1(N7057), .DIN2(N7826) );
and4s1 U2148 ( .Q(N8405), .DIN1(N7098), .DIN2(N7077), .DIN3(N7073), .DIN4(N7068) );
and2s1 U2149 ( .Q(N8409), .DIN1(N7068), .DIN2(N4632) );
and3s1 U2150 ( .Q(N8410), .DIN1(N7073), .DIN2(N7068), .DIN3(N4634) );
and4s1 U2151 ( .Q(N8411), .DIN1(N7077), .DIN2(N7068), .DIN3(N4635), .DIN4(N7073) );
and5s1 U2152 ( .Q(N8412), .DIN1(N7099), .DIN2(N7095), .DIN3(N7091), .DIN4(N7086), .DIN5(N7080) );
and2s1 U2153 ( .Q(N8415), .DIN1(N7080), .DIN2(N4638) );
and3s1 U2154 ( .Q(N8416), .DIN1(N7086), .DIN2(N7080), .DIN3(N4639) );
and4s1 U2155 ( .Q(N8417), .DIN1(N7091), .DIN2(N7080), .DIN3(N4640), .DIN4(N7086) );
and5s1 U2156 ( .Q(N8418), .DIN1(N7095), .DIN2(N7091), .DIN3(N7080), .DIN4(N4641), .DIN5(N7086) );
and2s1 U2157 ( .Q(N8421), .DIN1(N3375), .DIN2(N7100) );
and4s1 U2158 ( .Q(N8430), .DIN1(N7114), .DIN2(N7136), .DIN3(N7125), .DIN4(N7107) );
and2s1 U2159 ( .Q(N8433), .DIN1(N7107), .DIN2(N4657) );
and3s1 U2160 ( .Q(N8434), .DIN1(N7114), .DIN2(N7107), .DIN3(N4661) );
and4s1 U2161 ( .Q(N8435), .DIN1(N7125), .DIN2(N7107), .DIN3(N4667), .DIN4(N7114) );
and2s1 U2162 ( .Q(N8436), .DIN1(N7114), .DIN2(N4661) );
and3s1 U2163 ( .Q(N8437), .DIN1(N7125), .DIN2(N4667), .DIN3(N7114) );
and3s1 U2164 ( .Q(N8438), .DIN1(N7136), .DIN2(N7125), .DIN3(N7114) );
and2s1 U2165 ( .Q(N8439), .DIN1(N7114), .DIN2(N4661) );
and3s1 U2166 ( .Q(N8440), .DIN1(N4667), .DIN2(N7125), .DIN3(N7114) );
and2s1 U2167 ( .Q(N8441), .DIN1(N7125), .DIN2(N4667) );
and2s1 U2168 ( .Q(N8442), .DIN1(N7136), .DIN2(N7125) );
and2s1 U2169 ( .Q(N8443), .DIN1(N7125), .DIN2(N4667) );
and5s1 U2170 ( .Q(N8444), .DIN1(N7149), .DIN2(N7180), .DIN3(N7159), .DIN4(N7142), .DIN5(N7170) );
and2s1 U2171 ( .Q(N8447), .DIN1(N7142), .DIN2(N4675) );
and3s1 U2172 ( .Q(N8448), .DIN1(N7149), .DIN2(N7142), .DIN3(N4678) );
and4s1 U2173 ( .Q(N8449), .DIN1(N7159), .DIN2(N7142), .DIN3(N4682), .DIN4(N7149) );
and5s1 U2174 ( .Q(N8450), .DIN1(N7170), .DIN2(N7159), .DIN3(N7142), .DIN4(N4687), .DIN5(N7149) );
and2s1 U2175 ( .Q(N8451), .DIN1(N7149), .DIN2(N4678) );
and3s1 U2176 ( .Q(N8452), .DIN1(N7159), .DIN2(N4682), .DIN3(N7149) );
and4s1 U2177 ( .Q(N8453), .DIN1(N7170), .DIN2(N7159), .DIN3(N4687), .DIN4(N7149) );
and2s1 U2178 ( .Q(N8454), .DIN1(N4682), .DIN2(N7159) );
and3s1 U2179 ( .Q(N8455), .DIN1(N7170), .DIN2(N7159), .DIN3(N4687) );
and2s1 U2180 ( .Q(N8456), .DIN1(N7170), .DIN2(N4687) );
hi1s1 U2181 ( .Q(N8457), .DIN(N7194) );
hi1s1 U2182 ( .Q(N8460), .DIN(N7198) );
hi1s1 U2183 ( .Q(N8463), .DIN(N7205) );
hi1s1 U2184 ( .Q(N8466), .DIN(N7209) );
hi1s1 U2185 ( .Q(N8469), .DIN(N7216) );
hi1s1 U2186 ( .Q(N8470), .DIN(N7219) );
nb1s1 U2187 ( .Q(N8471), .DIN(N7202) );
nb1s1 U2188 ( .Q(N8474), .DIN(N7202) );
nb1s1 U2189 ( .Q(N8477), .DIN(N7213) );
nb1s1 U2190 ( .Q(N8480), .DIN(N7213) );
and3s1 U2191 ( .Q(N8483), .DIN1(N6083), .DIN2(N6079), .DIN3(N7216) );
and3s1 U2192 ( .Q(N8484), .DIN1(N7191), .DIN2(N7188), .DIN3(N7219) );
and4s1 U2193 ( .Q(N8485), .DIN1(N7301), .DIN2(N7240), .DIN3(N7229), .DIN4(N7222) );
and2s1 U2194 ( .Q(N8488), .DIN1(N7222), .DIN2(N4702) );
and3s1 U2195 ( .Q(N8489), .DIN1(N7229), .DIN2(N7222), .DIN3(N4706) );
and4s1 U2196 ( .Q(N8490), .DIN1(N7240), .DIN2(N7222), .DIN3(N4711), .DIN4(N7229) );
and2s1 U2197 ( .Q(N8491), .DIN1(N7229), .DIN2(N4706) );
and3s1 U2198 ( .Q(N8492), .DIN1(N7240), .DIN2(N4711), .DIN3(N7229) );
and3s1 U2199 ( .Q(N8493), .DIN1(N7301), .DIN2(N7240), .DIN3(N7229) );
and2s1 U2200 ( .Q(N8494), .DIN1(N7229), .DIN2(N4706) );
and3s1 U2201 ( .Q(N8495), .DIN1(N7240), .DIN2(N4711), .DIN3(N7229) );
and2s1 U2202 ( .Q(N8496), .DIN1(N7240), .DIN2(N4711) );
and5s1 U2203 ( .Q(N8497), .DIN1(N7307), .DIN2(N7288), .DIN3(N7272), .DIN4(N7258), .DIN5(N7250) );
and2s1 U2204 ( .Q(N8500), .DIN1(N7250), .DIN2(N4718) );
and3s1 U2205 ( .Q(N8501), .DIN1(N7258), .DIN2(N7250), .DIN3(N4722) );
and4s1 U2206 ( .Q(N8502), .DIN1(N7272), .DIN2(N7250), .DIN3(N4728), .DIN4(N7258) );
and5s1 U2207 ( .Q(N8503), .DIN1(N7288), .DIN2(N7272), .DIN3(N7250), .DIN4(N4735), .DIN5(N7258) );
and2s1 U2208 ( .Q(N8504), .DIN1(N7258), .DIN2(N4722) );
and3s1 U2209 ( .Q(N8505), .DIN1(N7272), .DIN2(N4728), .DIN3(N7258) );
and4s1 U2210 ( .Q(N8506), .DIN1(N7288), .DIN2(N7272), .DIN3(N4735), .DIN4(N7258) );
and4s1 U2211 ( .Q(N8507), .DIN1(N7307), .DIN2(N7272), .DIN3(N7258), .DIN4(N7288) );
and2s1 U2212 ( .Q(N8508), .DIN1(N7258), .DIN2(N4722) );
and3s1 U2213 ( .Q(N8509), .DIN1(N7272), .DIN2(N4728), .DIN3(N7258) );
and4s1 U2214 ( .Q(N8510), .DIN1(N7288), .DIN2(N7272), .DIN3(N4735), .DIN4(N7258) );
and2s1 U2215 ( .Q(N8511), .DIN1(N7272), .DIN2(N4728) );
and3s1 U2216 ( .Q(N8512), .DIN1(N7288), .DIN2(N7272), .DIN3(N4735) );
and3s1 U2217 ( .Q(N8513), .DIN1(N7307), .DIN2(N7272), .DIN3(N7288) );
and2s1 U2218 ( .Q(N8514), .DIN1(N7272), .DIN2(N4728) );
and3s1 U2219 ( .Q(N8515), .DIN1(N7288), .DIN2(N7272), .DIN3(N4735) );
and2s1 U2220 ( .Q(N8516), .DIN1(N7288), .DIN2(N4735) );
and2s1 U2221 ( .Q(N8517), .DIN1(N7301), .DIN2(N7240) );
and2s1 U2222 ( .Q(N8518), .DIN1(N7307), .DIN2(N7288) );
hi1s1 U2223 ( .Q(N8519), .DIN(N7314) );
hi1s1 U2224 ( .Q(N8522), .DIN(N7318) );
nb1s1 U2225 ( .Q(N8525), .DIN(N7322) );
nb1s1 U2226 ( .Q(N8528), .DIN(N7322) );
nb1s1 U2227 ( .Q(N8531), .DIN(N7331) );
nb1s1 U2228 ( .Q(N8534), .DIN(N7331) );
hi1s1 U2229 ( .Q(N8537), .DIN(N7340) );
hi1s1 U2230 ( .Q(N8538), .DIN(N7343) );
and3s1 U2231 ( .Q(N8539), .DIN1(N6141), .DIN2(N6137), .DIN3(N7340) );
and3s1 U2232 ( .Q(N8540), .DIN1(N7337), .DIN2(N7334), .DIN3(N7343) );
and4s1 U2233 ( .Q(N8541), .DIN1(N7376), .DIN2(N7355), .DIN3(N7351), .DIN4(N7346) );
and2s1 U2234 ( .Q(N8545), .DIN1(N7346), .DIN2(N4757) );
and3s1 U2235 ( .Q(N8546), .DIN1(N7351), .DIN2(N7346), .DIN3(N4758) );
and4s1 U2236 ( .Q(N8547), .DIN1(N7355), .DIN2(N7346), .DIN3(N4759), .DIN4(N7351) );
and5s1 U2237 ( .Q(N8548), .DIN1(N7377), .DIN2(N7373), .DIN3(N7369), .DIN4(N7364), .DIN5(N7358) );
and2s1 U2238 ( .Q(N8551), .DIN1(N7358), .DIN2(N4762) );
and3s1 U2239 ( .Q(N8552), .DIN1(N7364), .DIN2(N7358), .DIN3(N4764) );
and4s1 U2240 ( .Q(N8553), .DIN1(N7369), .DIN2(N7358), .DIN3(N4766), .DIN4(N7364) );
and5s1 U2241 ( .Q(N8554), .DIN1(N7373), .DIN2(N7369), .DIN3(N7358), .DIN4(N4767), .DIN5(N7364) );
hi1s1 U2242 ( .Q(N8555), .DIN(N7387) );
hi1s1 U2243 ( .Q(N8558), .DIN(N7394) );
hi1s1 U2244 ( .Q(N8561), .DIN(N7398) );
hi1s1 U2245 ( .Q(N8564), .DIN(N7405) );
hi1s1 U2246 ( .Q(N8565), .DIN(N7408) );
nb1s1 U2247 ( .Q(N8566), .DIN(N7391) );
nb1s1 U2248 ( .Q(N8569), .DIN(N7391) );
nb1s1 U2249 ( .Q(N8572), .DIN(N7402) );
nb1s1 U2250 ( .Q(N8575), .DIN(N7402) );
and3s1 U2251 ( .Q(N8578), .DIN1(N6170), .DIN2(N6166), .DIN3(N7405) );
and3s1 U2252 ( .Q(N8579), .DIN1(N7381), .DIN2(N7378), .DIN3(N7408) );
nb1s1 U2253 ( .Q(N8580), .DIN(N7180) );
nb1s1 U2254 ( .Q(N8583), .DIN(N7142) );
nb1s1 U2255 ( .Q(N8586), .DIN(N7149) );
nb1s1 U2256 ( .Q(N8589), .DIN(N7159) );
nb1s1 U2257 ( .Q(N8592), .DIN(N7170) );
nb1s1 U2258 ( .Q(N8595), .DIN(N6929) );
nb1s1 U2259 ( .Q(N8598), .DIN(N6936) );
nb1s1 U2260 ( .Q(N8601), .DIN(N6946) );
nb1s1 U2261 ( .Q(N8604), .DIN(N6957) );
hi1s1 U2262 ( .Q(N8607), .DIN(N7441) );
nnd2s1 U2263 ( .Q(N8608), .DIN1(N7441), .DIN2(N5469) );
hi1s1 U2264 ( .Q(N8609), .DIN(N7444) );
nnd2s1 U2265 ( .Q(N8610), .DIN1(N7444), .DIN2(N4793) );
hi1s1 U2266 ( .Q(N8615), .DIN(N7447) );
hi1s1 U2267 ( .Q(N8616), .DIN(N7450) );
hi1s1 U2268 ( .Q(N8617), .DIN(N7453) );
hi1s1 U2269 ( .Q(N8618), .DIN(N7456) );
hi1s1 U2270 ( .Q(N8619), .DIN(N7474) );
hi1s1 U2271 ( .Q(N8624), .DIN(N7465) );
hi1s1 U2272 ( .Q(N8625), .DIN(N7468) );
hi1s1 U2273 ( .Q(N8626), .DIN(N7471) );
nnd2s1 U2274 ( .Q(N8627), .DIN1(N8144), .DIN2(N8145) );
hi1s1 U2275 ( .Q(N8632), .DIN(N7479) );
hi1s1 U2276 ( .Q(N8633), .DIN(N7482) );
hi1s1 U2277 ( .Q(N8634), .DIN(N7485) );
hi1s1 U2278 ( .Q(N8637), .DIN(N7491) );
hi1s1 U2279 ( .Q(N8638), .DIN(N7494) );
hi1s1 U2280 ( .Q(N8639), .DIN(N7497) );
hi1s1 U2281 ( .Q(N8644), .DIN(N7503) );
hi1s1 U2282 ( .Q(N8645), .DIN(N7506) );
hi1s1 U2283 ( .Q(N8646), .DIN(N7509) );
hi1s1 U2284 ( .Q(N8647), .DIN(N7512) );
hi1s1 U2285 ( .Q(N8648), .DIN(N7530) );
hi1s1 U2286 ( .Q(N8653), .DIN(N7521) );
hi1s1 U2287 ( .Q(N8654), .DIN(N7524) );
hi1s1 U2288 ( .Q(N8655), .DIN(N7527) );
nb1s1 U2289 ( .Q(N8660), .DIN(N6894) );
nb1s1 U2290 ( .Q(N8663), .DIN(N6894) );
nb1s1 U2291 ( .Q(N8666), .DIN(N6901) );
nb1s1 U2292 ( .Q(N8669), .DIN(N6901) );
nb1s1 U2293 ( .Q(N8672), .DIN(N6912) );
nb1s1 U2294 ( .Q(N8675), .DIN(N6912) );
nb1s1 U2295 ( .Q(N8678), .DIN(N7049) );
nb1s1 U2296 ( .Q(N8681), .DIN(N6988) );
nb1s1 U2297 ( .Q(N8684), .DIN(N6970) );
nb1s1 U2298 ( .Q(N8687), .DIN(N6977) );
nb1s1 U2299 ( .Q(N8690), .DIN(N7049) );
nb1s1 U2300 ( .Q(N8693), .DIN(N6988) );
nb1s1 U2301 ( .Q(N8696), .DIN(N6970) );
nb1s1 U2302 ( .Q(N8699), .DIN(N6977) );
nb1s1 U2303 ( .Q(N8702), .DIN(N7036) );
nb1s1 U2304 ( .Q(N8705), .DIN(N6998) );
nb1s1 U2305 ( .Q(N8708), .DIN(N7020) );
nb1s1 U2306 ( .Q(N8711), .DIN(N7006) );
nb1s1 U2307 ( .Q(N8714), .DIN(N7006) );
hi1s1 U2308 ( .Q(N8717), .DIN(N7553) );
nb1s1 U2309 ( .Q(N8718), .DIN(N7036) );
nb1s1 U2310 ( .Q(N8721), .DIN(N6998) );
nb1s1 U2311 ( .Q(N8724), .DIN(N7020) );
nnd2s1 U2312 ( .Q(N8727), .DIN1(N8216), .DIN2(N8217) );
nnd2s1 U2313 ( .Q(N8730), .DIN1(N8218), .DIN2(N8219) );
hi1s1 U2314 ( .Q(N8733), .DIN(N7574) );
hi1s1 U2315 ( .Q(N8734), .DIN(N7577) );
nb1s1 U2316 ( .Q(N8735), .DIN(N7107) );
nb1s1 U2317 ( .Q(N8738), .DIN(N7107) );
nb1s1 U2318 ( .Q(N8741), .DIN(N7114) );
nb1s1 U2319 ( .Q(N8744), .DIN(N7114) );
nb1s1 U2320 ( .Q(N8747), .DIN(N7125) );
nb1s1 U2321 ( .Q(N8750), .DIN(N7125) );
hi1s1 U2322 ( .Q(N8753), .DIN(N7560) );
hi1s1 U2323 ( .Q(N8754), .DIN(N7563) );
hi1s1 U2324 ( .Q(N8755), .DIN(N7566) );
hi1s1 U2325 ( .Q(N8756), .DIN(N7569) );
nb1s1 U2326 ( .Q(N8757), .DIN(N7301) );
nb1s1 U2327 ( .Q(N8760), .DIN(N7240) );
nb1s1 U2328 ( .Q(N8763), .DIN(N7222) );
nb1s1 U2329 ( .Q(N8766), .DIN(N7229) );
nb1s1 U2330 ( .Q(N8769), .DIN(N7301) );
nb1s1 U2331 ( .Q(N8772), .DIN(N7240) );
nb1s1 U2332 ( .Q(N8775), .DIN(N7222) );
nb1s1 U2333 ( .Q(N8778), .DIN(N7229) );
nb1s1 U2334 ( .Q(N8781), .DIN(N7307) );
nb1s1 U2335 ( .Q(N8784), .DIN(N7288) );
nb1s1 U2336 ( .Q(N8787), .DIN(N7250) );
nb1s1 U2337 ( .Q(N8790), .DIN(N7272) );
nb1s1 U2338 ( .Q(N8793), .DIN(N7258) );
nb1s1 U2339 ( .Q(N8796), .DIN(N7258) );
nb1s1 U2340 ( .Q(N8799), .DIN(N7307) );
nb1s1 U2341 ( .Q(N8802), .DIN(N7288) );
nb1s1 U2342 ( .Q(N8805), .DIN(N7250) );
nb1s1 U2343 ( .Q(N8808), .DIN(N7272) );
nnd2s1 U2344 ( .Q(N8811), .DIN1(N8232), .DIN2(N8233) );
hi1s1 U2345 ( .Q(N8814), .DIN(N7588) );
hi1s1 U2346 ( .Q(N8815), .DIN(N7591) );
hi1s1 U2347 ( .Q(N8816), .DIN(N7582) );
hi1s1 U2348 ( .Q(N8817), .DIN(N7585) );
and2s1 U2349 ( .Q(N8818), .DIN1(N7620), .DIN2(N3155) );
and2s1 U2350 ( .Q(N8840), .DIN1(N3122), .DIN2(N7609) );
hi1s1 U2351 ( .Q(N8857), .DIN(N7609) );
and3s1 U2352 ( .Q(N8861), .DIN1(N6797), .DIN2(N5740), .DIN3(N8274) );
and3s1 U2353 ( .Q(N8862), .DIN1(N5736), .DIN2(N6800), .DIN3(N8275) );
and3s1 U2354 ( .Q(N8863), .DIN1(N6803), .DIN2(N5751), .DIN3(N8276) );
and3s1 U2355 ( .Q(N8864), .DIN1(N5747), .DIN2(N6806), .DIN3(N8277) );
and3s1 U2356 ( .Q(N8865), .DIN1(N6809), .DIN2(N5762), .DIN3(N8278) );
and3s1 U2357 ( .Q(N8866), .DIN1(N5758), .DIN2(N6812), .DIN3(N8279) );
hi1s1 U2358 ( .Q(N8871), .DIN(N7655) );
and2s1 U2359 ( .Q(N8874), .DIN1(N6833), .DIN2(N7655) );
and2s1 U2360 ( .Q(N8878), .DIN1(N7671), .DIN2(N6867) );
hi1s1 U2361 ( .Q(N8879), .DIN(N8196) );
nnd2s1 U2362 ( .Q(N8880), .DIN1(N8196), .DIN2(N8315) );
hi1s1 U2363 ( .Q(N8881), .DIN(N8200) );
nnd2s1 U2364 ( .Q(N8882), .DIN1(N8200), .DIN2(N8317) );
hi1s1 U2365 ( .Q(N8883), .DIN(N8204) );
nnd2s1 U2366 ( .Q(N8884), .DIN1(N8204), .DIN2(N8319) );
hi1s1 U2367 ( .Q(N8885), .DIN(N8208) );
nnd2s1 U2368 ( .Q(N8886), .DIN1(N8208), .DIN2(N8321) );
nnd2s1 U2369 ( .Q(N8887), .DIN1(N3658), .DIN2(N8323) );
nnd2s1 U2370 ( .Q(N8888), .DIN1(N4817), .DIN2(N8325) );
or4s1 U2371 ( .Q(N8898), .DIN1(N4544), .DIN2(N8337), .DIN3(N8338), .DIN4(N8339) );
or5s1 U2372 ( .Q(N8902), .DIN1(N4562), .DIN2(N8348), .DIN3(N8349), .DIN4(N8350), .DIN5(N8351) );
or4s1 U2373 ( .Q(N8920), .DIN1(N4576), .DIN2(N8369), .DIN3(N8370), .DIN4(N8371) );
or2s1 U2374 ( .Q(N8924), .DIN1(N4581), .DIN2(N8377) );
or5s1 U2375 ( .Q(N8927), .DIN1(N4592), .DIN2(N8378), .DIN3(N8379), .DIN4(N8380), .DIN5(N8381) );
or2s1 U2376 ( .Q(N8931), .DIN1(N4603), .DIN2(N8392) );
or2s1 U2377 ( .Q(N8943), .DIN1(N7825), .DIN2(N8404) );
or4s1 U2378 ( .Q(N8950), .DIN1(N4630), .DIN2(N8409), .DIN3(N8410), .DIN4(N8411) );
or5s1 U2379 ( .Q(N8956), .DIN1(N4637), .DIN2(N8415), .DIN3(N8416), .DIN4(N8417), .DIN5(N8418) );
hi1s1 U2380 ( .Q(N8959), .DIN(N7852) );
and2s1 U2381 ( .Q(N8960), .DIN1(N3375), .DIN2(N7852) );
or4s1 U2382 ( .Q(N8963), .DIN1(N4656), .DIN2(N8433), .DIN3(N8434), .DIN4(N8435) );
or5s1 U2383 ( .Q(N8966), .DIN1(N4674), .DIN2(N8447), .DIN3(N8448), .DIN4(N8449), .DIN5(N8450) );
and3s1 U2384 ( .Q(N8991), .DIN1(N7188), .DIN2(N6083), .DIN3(N8469) );
and3s1 U2385 ( .Q(N8992), .DIN1(N6079), .DIN2(N7191), .DIN3(N8470) );
or4s1 U2386 ( .Q(N8995), .DIN1(N4701), .DIN2(N8488), .DIN3(N8489), .DIN4(N8490) );
or2s1 U2387 ( .Q(N8996), .DIN1(N4706), .DIN2(N8496) );
or5s1 U2388 ( .Q(N9001), .DIN1(N4717), .DIN2(N8500), .DIN3(N8501), .DIN4(N8502), .DIN5(N8503) );
or2s1 U2389 ( .Q(N9005), .DIN1(N4728), .DIN2(N8516) );
and3s1 U2390 ( .Q(N9024), .DIN1(N7334), .DIN2(N6141), .DIN3(N8537) );
and3s1 U2391 ( .Q(N9025), .DIN1(N6137), .DIN2(N7337), .DIN3(N8538) );
or4s1 U2392 ( .Q(N9029), .DIN1(N4756), .DIN2(N8545), .DIN3(N8546), .DIN4(N8547) );
or5s1 U2393 ( .Q(N9035), .DIN1(N4760), .DIN2(N8551), .DIN3(N8552), .DIN4(N8553), .DIN5(N8554) );
and3s1 U2394 ( .Q(N9053), .DIN1(N7378), .DIN2(N6170), .DIN3(N8564) );
and3s1 U2395 ( .Q(N9054), .DIN1(N6166), .DIN2(N7381), .DIN3(N8565) );
nnd2s1 U2396 ( .Q(N9064), .DIN1(N4303), .DIN2(N8607) );
nnd2s1 U2397 ( .Q(N9065), .DIN1(N3507), .DIN2(N8609) );
hi1s1 U2398 ( .Q(N9066), .DIN(N8114) );
nnd2s1 U2399 ( .Q(N9067), .DIN1(N8114), .DIN2(N4795) );
or2s1 U2400 ( .Q(N9068), .DIN1(N7613), .DIN2(N6783) );
hi1s1 U2401 ( .Q(N9071), .DIN(N8117) );
hi1s1 U2402 ( .Q(N9072), .DIN(N8131) );
nnd2s1 U2403 ( .Q(N9073), .DIN1(N8131), .DIN2(N6195) );
hi1s1 U2404 ( .Q(N9074), .DIN(N7613) );
hi1s1 U2405 ( .Q(N9077), .DIN(N8134) );
or2s1 U2406 ( .Q(N9079), .DIN1(N7650), .DIN2(N6865) );
hi1s1 U2407 ( .Q(N9082), .DIN(N8146) );
hi1s1 U2408 ( .Q(N9083), .DIN(N7650) );
hi1s1 U2409 ( .Q(N9086), .DIN(N8156) );
hi1s1 U2410 ( .Q(N9087), .DIN(N8166) );
nnd2s1 U2411 ( .Q(N9088), .DIN1(N8166), .DIN2(N4813) );
or2s1 U2412 ( .Q(N9089), .DIN1(N7659), .DIN2(N6866) );
hi1s1 U2413 ( .Q(N9092), .DIN(N8169) );
hi1s1 U2414 ( .Q(N9093), .DIN(N8183) );
nnd2s1 U2415 ( .Q(N9094), .DIN1(N8183), .DIN2(N6203) );
hi1s1 U2416 ( .Q(N9095), .DIN(N7659) );
hi1s1 U2417 ( .Q(N9098), .DIN(N8186) );
or4s1 U2418 ( .Q(N9099), .DIN1(N4545), .DIN2(N8340), .DIN3(N8341), .DIN4(N8342) );
nor3s1 U2419 ( .Q(N9103), .DIN1(N4545), .DIN2(N8343), .DIN3(N8344) );
or3s1 U2420 ( .Q(N9107), .DIN1(N4549), .DIN2(N8345), .DIN3(N8346) );
nor2s1 U2421 ( .Q(N9111), .DIN1(N4549), .DIN2(N8347) );
or4s1 U2422 ( .Q(N9117), .DIN1(N4577), .DIN2(N8372), .DIN3(N8373), .DIN4(N8374) );
nor3s1 U2423 ( .Q(N9127), .DIN1(N4577), .DIN2(N8375), .DIN3(N8376) );
nor3s1 U2424 ( .Q(N9146), .DIN1(N4597), .DIN2(N8390), .DIN3(N8391) );
nor4s1 U2425 ( .Q(N9149), .DIN1(N4593), .DIN2(N8385), .DIN3(N8386), .DIN4(N8387) );
nnd2s1 U2426 ( .Q(N9159), .DIN1(N7577), .DIN2(N8733) );
nnd2s1 U2427 ( .Q(N9160), .DIN1(N7574), .DIN2(N8734) );
or4s1 U2428 ( .Q(N9161), .DIN1(N4657), .DIN2(N8436), .DIN3(N8437), .DIN4(N8438) );
nor3s1 U2429 ( .Q(N9165), .DIN1(N4657), .DIN2(N8439), .DIN3(N8440) );
or3s1 U2430 ( .Q(N9169), .DIN1(N4661), .DIN2(N8441), .DIN3(N8442) );
nor2s1 U2431 ( .Q(N9173), .DIN1(N4661), .DIN2(N8443) );
nnd2s1 U2432 ( .Q(N9179), .DIN1(N7563), .DIN2(N8753) );
nnd2s1 U2433 ( .Q(N9180), .DIN1(N7560), .DIN2(N8754) );
nnd2s1 U2434 ( .Q(N9181), .DIN1(N7569), .DIN2(N8755) );
nnd2s1 U2435 ( .Q(N9182), .DIN1(N7566), .DIN2(N8756) );
or4s1 U2436 ( .Q(N9183), .DIN1(N4702), .DIN2(N8491), .DIN3(N8492), .DIN4(N8493) );
nor3s1 U2437 ( .Q(N9193), .DIN1(N4702), .DIN2(N8494), .DIN3(N8495) );
or4s1 U2438 ( .Q(N9203), .DIN1(N4722), .DIN2(N8511), .DIN3(N8512), .DIN4(N8513) );
or5s1 U2439 ( .Q(N9206), .DIN1(N4718), .DIN2(N8504), .DIN3(N8505), .DIN4(N8506), .DIN5(N8507) );
nor3s1 U2440 ( .Q(N9220), .DIN1(N4722), .DIN2(N8514), .DIN3(N8515) );
nor4s1 U2441 ( .Q(N9223), .DIN1(N4718), .DIN2(N8508), .DIN3(N8509), .DIN4(N8510) );
nnd2s1 U2442 ( .Q(N9234), .DIN1(N7591), .DIN2(N8814) );
nnd2s1 U2443 ( .Q(N9235), .DIN1(N7588), .DIN2(N8815) );
nnd2s1 U2444 ( .Q(N9236), .DIN1(N7585), .DIN2(N8816) );
nnd2s1 U2445 ( .Q(N9237), .DIN1(N7582), .DIN2(N8817) );
or2s1 U2446 ( .Q(N9238), .DIN1(N3159), .DIN2(N8818) );
or2s1 U2447 ( .Q(N9242), .DIN1(N3126), .DIN2(N8840) );
nnd2s1 U2448 ( .Q(N9243), .DIN1(N8324), .DIN2(N8888) );
hi1s1 U2449 ( .Q(N9244), .DIN(N8580) );
hi1s1 U2450 ( .Q(N9245), .DIN(N8583) );
hi1s1 U2451 ( .Q(N9246), .DIN(N8586) );
hi1s1 U2452 ( .Q(N9247), .DIN(N8589) );
hi1s1 U2453 ( .Q(N9248), .DIN(N8592) );
hi1s1 U2454 ( .Q(N9249), .DIN(N8595) );
hi1s1 U2455 ( .Q(N9250), .DIN(N8598) );
hi1s1 U2456 ( .Q(N9251), .DIN(N8601) );
hi1s1 U2457 ( .Q(N9252), .DIN(N8604) );
nor2s1 U2458 ( .Q(N9256), .DIN1(N8861), .DIN2(N8280) );
nor2s1 U2459 ( .Q(N9257), .DIN1(N8862), .DIN2(N8281) );
nor2s1 U2460 ( .Q(N9258), .DIN1(N8863), .DIN2(N8282) );
nor2s1 U2461 ( .Q(N9259), .DIN1(N8864), .DIN2(N8283) );
nor2s1 U2462 ( .Q(N9260), .DIN1(N8865), .DIN2(N8284) );
nor2s1 U2463 ( .Q(N9261), .DIN1(N8866), .DIN2(N8285) );
hi1s1 U2464 ( .Q(N9262), .DIN(N8627) );
or2s1 U2465 ( .Q(N9265), .DIN1(N7649), .DIN2(N8874) );
or2s1 U2466 ( .Q(N9268), .DIN1(N7668), .DIN2(N8878) );
nnd2s1 U2467 ( .Q(N9271), .DIN1(N7533), .DIN2(N8879) );
nnd2s1 U2468 ( .Q(N9272), .DIN1(N7536), .DIN2(N8881) );
nnd2s1 U2469 ( .Q(N9273), .DIN1(N7539), .DIN2(N8883) );
nnd2s1 U2470 ( .Q(N9274), .DIN1(N7542), .DIN2(N8885) );
nnd2s1 U2471 ( .Q(N9275), .DIN1(N8322), .DIN2(N8887) );
hi1s1 U2472 ( .Q(N9276), .DIN(N8333) );
and5s1 U2473 ( .Q(N9280), .DIN1(N6936), .DIN2(N8326), .DIN3(N6946), .DIN4(N6929), .DIN5(N6957) );
and5s1 U2474 ( .Q(N9285), .DIN1(N367), .DIN2(N8326), .DIN3(N6946), .DIN4(N6957), .DIN5(N6936) );
and4s1 U2475 ( .Q(N9286), .DIN1(N367), .DIN2(N8326), .DIN3(N6946), .DIN4(N6957) );
and3s1 U2476 ( .Q(N9287), .DIN1(N367), .DIN2(N8326), .DIN3(N6957) );
and2s1 U2477 ( .Q(N9288), .DIN1(N367), .DIN2(N8326) );
hi1s1 U2478 ( .Q(N9290), .DIN(N8660) );
hi1s1 U2479 ( .Q(N9292), .DIN(N8663) );
hi1s1 U2480 ( .Q(N9294), .DIN(N8666) );
hi1s1 U2481 ( .Q(N9296), .DIN(N8669) );
nnd2s1 U2482 ( .Q(N9297), .DIN1(N8672), .DIN2(N5966) );
hi1s1 U2483 ( .Q(N9298), .DIN(N8672) );
nnd2s1 U2484 ( .Q(N9299), .DIN1(N8675), .DIN2(N6969) );
hi1s1 U2485 ( .Q(N9300), .DIN(N8675) );
hi1s1 U2486 ( .Q(N9301), .DIN(N8365) );
and5s1 U2487 ( .Q(N9307), .DIN1(N8358), .DIN2(N7036), .DIN3(N7020), .DIN4(N7006), .DIN5(N6998) );
and4s1 U2488 ( .Q(N9314), .DIN1(N8358), .DIN2(N7020), .DIN3(N7006), .DIN4(N7036) );
and3s1 U2489 ( .Q(N9315), .DIN1(N8358), .DIN2(N7020), .DIN3(N7036) );
and2s1 U2490 ( .Q(N9318), .DIN1(N8358), .DIN2(N7036) );
hi1s1 U2491 ( .Q(N9319), .DIN(N8687) );
hi1s1 U2492 ( .Q(N9320), .DIN(N8699) );
hi1s1 U2493 ( .Q(N9321), .DIN(N8711) );
hi1s1 U2494 ( .Q(N9322), .DIN(N8714) );
hi1s1 U2495 ( .Q(N9323), .DIN(N8727) );
hi1s1 U2496 ( .Q(N9324), .DIN(N8730) );
hi1s1 U2497 ( .Q(N9326), .DIN(N8405) );
and2s1 U2498 ( .Q(N9332), .DIN1(N8405), .DIN2(N8412) );
or2s1 U2499 ( .Q(N9339), .DIN1(N4193), .DIN2(N8960) );
and2s1 U2500 ( .Q(N9344), .DIN1(N8430), .DIN2(N8444) );
hi1s1 U2501 ( .Q(N9352), .DIN(N8735) );
hi1s1 U2502 ( .Q(N9354), .DIN(N8738) );
hi1s1 U2503 ( .Q(N9356), .DIN(N8741) );
hi1s1 U2504 ( .Q(N9358), .DIN(N8744) );
nnd2s1 U2505 ( .Q(N9359), .DIN1(N8747), .DIN2(N6078) );
hi1s1 U2506 ( .Q(N9360), .DIN(N8747) );
nnd2s1 U2507 ( .Q(N9361), .DIN1(N8750), .DIN2(N7187) );
hi1s1 U2508 ( .Q(N9362), .DIN(N8750) );
hi1s1 U2509 ( .Q(N9363), .DIN(N8471) );
hi1s1 U2510 ( .Q(N9364), .DIN(N8474) );
hi1s1 U2511 ( .Q(N9365), .DIN(N8477) );
hi1s1 U2512 ( .Q(N9366), .DIN(N8480) );
nor2s1 U2513 ( .Q(N9367), .DIN1(N8991), .DIN2(N8483) );
nor2s1 U2514 ( .Q(N9368), .DIN1(N8992), .DIN2(N8484) );
and3s1 U2515 ( .Q(N9369), .DIN1(N7198), .DIN2(N7194), .DIN3(N8471) );
and3s1 U2516 ( .Q(N9370), .DIN1(N8460), .DIN2(N8457), .DIN3(N8474) );
and3s1 U2517 ( .Q(N9371), .DIN1(N7209), .DIN2(N7205), .DIN3(N8477) );
and3s1 U2518 ( .Q(N9372), .DIN1(N8466), .DIN2(N8463), .DIN3(N8480) );
hi1s1 U2519 ( .Q(N9375), .DIN(N8497) );
hi1s1 U2520 ( .Q(N9381), .DIN(N8766) );
hi1s1 U2521 ( .Q(N9382), .DIN(N8778) );
hi1s1 U2522 ( .Q(N9383), .DIN(N8793) );
hi1s1 U2523 ( .Q(N9384), .DIN(N8796) );
and2s1 U2524 ( .Q(N9385), .DIN1(N8485), .DIN2(N8497) );
hi1s1 U2525 ( .Q(N9392), .DIN(N8525) );
hi1s1 U2526 ( .Q(N9393), .DIN(N8528) );
hi1s1 U2527 ( .Q(N9394), .DIN(N8531) );
hi1s1 U2528 ( .Q(N9395), .DIN(N8534) );
and3s1 U2529 ( .Q(N9396), .DIN1(N7318), .DIN2(N7314), .DIN3(N8525) );
and3s1 U2530 ( .Q(N9397), .DIN1(N8522), .DIN2(N8519), .DIN3(N8528) );
and3s1 U2531 ( .Q(N9398), .DIN1(N6131), .DIN2(N6127), .DIN3(N8531) );
and3s1 U2532 ( .Q(N9399), .DIN1(N7328), .DIN2(N7325), .DIN3(N8534) );
nor2s1 U2533 ( .Q(N9400), .DIN1(N9024), .DIN2(N8539) );
nor2s1 U2534 ( .Q(N9401), .DIN1(N9025), .DIN2(N8540) );
hi1s1 U2535 ( .Q(N9402), .DIN(N8541) );
nnd2s1 U2536 ( .Q(N9407), .DIN1(N8548), .DIN2(N89) );
and2s1 U2537 ( .Q(N9408), .DIN1(N8541), .DIN2(N8548) );
hi1s1 U2538 ( .Q(N9412), .DIN(N8811) );
hi1s1 U2539 ( .Q(N9413), .DIN(N8566) );
hi1s1 U2540 ( .Q(N9414), .DIN(N8569) );
hi1s1 U2541 ( .Q(N9415), .DIN(N8572) );
hi1s1 U2542 ( .Q(N9416), .DIN(N8575) );
nor2s1 U2543 ( .Q(N9417), .DIN1(N9053), .DIN2(N8578) );
nor2s1 U2544 ( .Q(N9418), .DIN1(N9054), .DIN2(N8579) );
and3s1 U2545 ( .Q(N9419), .DIN1(N7387), .DIN2(N6177), .DIN3(N8566) );
and3s1 U2546 ( .Q(N9420), .DIN1(N8555), .DIN2(N7384), .DIN3(N8569) );
and3s1 U2547 ( .Q(N9421), .DIN1(N7398), .DIN2(N7394), .DIN3(N8572) );
and3s1 U2548 ( .Q(N9422), .DIN1(N8561), .DIN2(N8558), .DIN3(N8575) );
nb1s1 U2549 ( .Q(N9423), .DIN(N8326) );
nnd2s1 U2550 ( .Q(N9426), .DIN1(N9064), .DIN2(N8608) );
nnd2s1 U2551 ( .Q(N9429), .DIN1(N9065), .DIN2(N8610) );
nnd2s1 U2552 ( .Q(N9432), .DIN1(N3515), .DIN2(N9066) );
nnd2s1 U2553 ( .Q(N9435), .DIN1(N4796), .DIN2(N9072) );
nnd2s1 U2554 ( .Q(N9442), .DIN1(N3628), .DIN2(N9087) );
nnd2s1 U2555 ( .Q(N9445), .DIN1(N4814), .DIN2(N9093) );
hi1s1 U2556 ( .Q(N9454), .DIN(N8678) );
hi1s1 U2557 ( .Q(N9455), .DIN(N8681) );
hi1s1 U2558 ( .Q(N9456), .DIN(N8684) );
hi1s1 U2559 ( .Q(N9459), .DIN(N8690) );
hi1s1 U2560 ( .Q(N9460), .DIN(N8693) );
hi1s1 U2561 ( .Q(N9461), .DIN(N8696) );
nb1s1 U2562 ( .Q(N9462), .DIN(N8358) );
hi1s1 U2563 ( .Q(N9465), .DIN(N8702) );
hi1s1 U2564 ( .Q(N9466), .DIN(N8705) );
hi1s1 U2565 ( .Q(N9467), .DIN(N8708) );
hi1s1 U2566 ( .Q(N9468), .DIN(N8724) );
nb1s1 U2567 ( .Q(N9473), .DIN(N8358) );
hi1s1 U2568 ( .Q(N9476), .DIN(N8718) );
hi1s1 U2569 ( .Q(N9477), .DIN(N8721) );
nnd2s1 U2570 ( .Q(N9478), .DIN1(N9159), .DIN2(N9160) );
nnd2s1 U2571 ( .Q(N9485), .DIN1(N9179), .DIN2(N9180) );
nnd2s1 U2572 ( .Q(N9488), .DIN1(N9181), .DIN2(N9182) );
hi1s1 U2573 ( .Q(N9493), .DIN(N8757) );
hi1s1 U2574 ( .Q(N9494), .DIN(N8760) );
hi1s1 U2575 ( .Q(N9495), .DIN(N8763) );
hi1s1 U2576 ( .Q(N9498), .DIN(N8769) );
hi1s1 U2577 ( .Q(N9499), .DIN(N8772) );
hi1s1 U2578 ( .Q(N9500), .DIN(N8775) );
hi1s1 U2579 ( .Q(N9505), .DIN(N8781) );
hi1s1 U2580 ( .Q(N9506), .DIN(N8784) );
hi1s1 U2581 ( .Q(N9507), .DIN(N8787) );
hi1s1 U2582 ( .Q(N9508), .DIN(N8790) );
hi1s1 U2583 ( .Q(N9509), .DIN(N8808) );
hi1s1 U2584 ( .Q(N9514), .DIN(N8799) );
hi1s1 U2585 ( .Q(N9515), .DIN(N8802) );
hi1s1 U2586 ( .Q(N9516), .DIN(N8805) );
nnd2s1 U2587 ( .Q(N9517), .DIN1(N9234), .DIN2(N9235) );
nnd2s1 U2588 ( .Q(N9520), .DIN1(N9236), .DIN2(N9237) );
and2s1 U2589 ( .Q(N9526), .DIN1(N8943), .DIN2(N8421) );
and2s1 U2590 ( .Q(N9531), .DIN1(N8943), .DIN2(N8421) );
nnd2s1 U2591 ( .Q(N9539), .DIN1(N9271), .DIN2(N8880) );
nnd2s1 U2592 ( .Q(N9540), .DIN1(N9273), .DIN2(N8884) );
hi1s1 U2593 ( .Q(N9541), .DIN(N9275) );
and2s1 U2594 ( .Q(N9543), .DIN1(N8857), .DIN2(N8254) );
and2s1 U2595 ( .Q(N9551), .DIN1(N8871), .DIN2(N8288) );
nnd2s1 U2596 ( .Q(N9555), .DIN1(N9272), .DIN2(N8882) );
nnd2s1 U2597 ( .Q(N9556), .DIN1(N9274), .DIN2(N8886) );
hi1s1 U2598 ( .Q(N9557), .DIN(N8898) );
and2s1 U2599 ( .Q(N9560), .DIN1(N8902), .DIN2(N8333) );
hi1s1 U2600 ( .Q(N9561), .DIN(N9099) );
nnd2s1 U2601 ( .Q(N9562), .DIN1(N9099), .DIN2(N9290) );
hi1s1 U2602 ( .Q(N9563), .DIN(N9103) );
nnd2s1 U2603 ( .Q(N9564), .DIN1(N9103), .DIN2(N9292) );
hi1s1 U2604 ( .Q(N9565), .DIN(N9107) );
nnd2s1 U2605 ( .Q(N9566), .DIN1(N9107), .DIN2(N9294) );
hi1s1 U2606 ( .Q(N9567), .DIN(N9111) );
nnd2s1 U2607 ( .Q(N9568), .DIN1(N9111), .DIN2(N9296) );
nnd2s1 U2608 ( .Q(N9569), .DIN1(N4844), .DIN2(N9298) );
nnd2s1 U2609 ( .Q(N9570), .DIN1(N6207), .DIN2(N9300) );
hi1s1 U2610 ( .Q(N9571), .DIN(N8920) );
hi1s1 U2611 ( .Q(N9575), .DIN(N8927) );
and2s1 U2612 ( .Q(N9579), .DIN1(N8365), .DIN2(N8927) );
hi1s1 U2613 ( .Q(N9581), .DIN(N8950) );
hi1s1 U2614 ( .Q(N9582), .DIN(N8956) );
and2s1 U2615 ( .Q(N9585), .DIN1(N8405), .DIN2(N8956) );
and2s1 U2616 ( .Q(N9591), .DIN1(N8966), .DIN2(N8430) );
hi1s1 U2617 ( .Q(N9592), .DIN(N9161) );
nnd2s1 U2618 ( .Q(N9593), .DIN1(N9161), .DIN2(N9352) );
hi1s1 U2619 ( .Q(N9594), .DIN(N9165) );
nnd2s1 U2620 ( .Q(N9595), .DIN1(N9165), .DIN2(N9354) );
hi1s1 U2621 ( .Q(N9596), .DIN(N9169) );
nnd2s1 U2622 ( .Q(N9597), .DIN1(N9169), .DIN2(N9356) );
hi1s1 U2623 ( .Q(N9598), .DIN(N9173) );
nnd2s1 U2624 ( .Q(N9599), .DIN1(N9173), .DIN2(N9358) );
nnd2s1 U2625 ( .Q(N9600), .DIN1(N4940), .DIN2(N9360) );
nnd2s1 U2626 ( .Q(N9601), .DIN1(N6220), .DIN2(N9362) );
and3s1 U2627 ( .Q(N9602), .DIN1(N8457), .DIN2(N7198), .DIN3(N9363) );
and3s1 U2628 ( .Q(N9603), .DIN1(N7194), .DIN2(N8460), .DIN3(N9364) );
and3s1 U2629 ( .Q(N9604), .DIN1(N8463), .DIN2(N7209), .DIN3(N9365) );
and3s1 U2630 ( .Q(N9605), .DIN1(N7205), .DIN2(N8466), .DIN3(N9366) );
hi1s1 U2631 ( .Q(N9608), .DIN(N9001) );
and2s1 U2632 ( .Q(N9611), .DIN1(N8485), .DIN2(N9001) );
and3s1 U2633 ( .Q(N9612), .DIN1(N8519), .DIN2(N7318), .DIN3(N9392) );
and3s1 U2634 ( .Q(N9613), .DIN1(N7314), .DIN2(N8522), .DIN3(N9393) );
and3s1 U2635 ( .Q(N9614), .DIN1(N7325), .DIN2(N6131), .DIN3(N9394) );
and3s1 U2636 ( .Q(N9615), .DIN1(N6127), .DIN2(N7328), .DIN3(N9395) );
hi1s1 U2637 ( .Q(N9616), .DIN(N9029) );
hi1s1 U2638 ( .Q(N9617), .DIN(N9035) );
and2s1 U2639 ( .Q(N9618), .DIN1(N8541), .DIN2(N9035) );
and3s1 U2640 ( .Q(N9621), .DIN1(N7384), .DIN2(N7387), .DIN3(N9413) );
and3s1 U2641 ( .Q(N9622), .DIN1(N6177), .DIN2(N8555), .DIN3(N9414) );
and3s1 U2642 ( .Q(N9623), .DIN1(N8558), .DIN2(N7398), .DIN3(N9415) );
and3s1 U2643 ( .Q(N9624), .DIN1(N7394), .DIN2(N8561), .DIN3(N9416) );
or5s1 U2644 ( .Q(N9626), .DIN1(N4563), .DIN2(N8352), .DIN3(N8353), .DIN4(N8354), .DIN5(N9285) );
or4s1 U2645 ( .Q(N9629), .DIN1(N4566), .DIN2(N8355), .DIN3(N8356), .DIN4(N9286) );
or3s1 U2646 ( .Q(N9632), .DIN1(N4570), .DIN2(N8357), .DIN3(N9287) );
or2s1 U2647 ( .Q(N9635), .DIN1(N5960), .DIN2(N9288) );
nnd2s1 U2648 ( .Q(N9642), .DIN1(N9067), .DIN2(N9432) );
hi1s1 U2649 ( .Q(N9645), .DIN(N9068) );
nnd2s1 U2650 ( .Q(N9646), .DIN1(N9073), .DIN2(N9435) );
hi1s1 U2651 ( .Q(N9649), .DIN(N9074) );
nnd2s1 U2652 ( .Q(N9650), .DIN1(N9257), .DIN2(N9256) );
nnd2s1 U2653 ( .Q(N9653), .DIN1(N9259), .DIN2(N9258) );
nnd2s1 U2654 ( .Q(N9656), .DIN1(N9261), .DIN2(N9260) );
hi1s1 U2655 ( .Q(N9659), .DIN(N9079) );
nnd2s1 U2656 ( .Q(N9660), .DIN1(N9079), .DIN2(N4809) );
hi1s1 U2657 ( .Q(N9661), .DIN(N9083) );
nnd2s1 U2658 ( .Q(N9662), .DIN1(N9083), .DIN2(N6202) );
nnd2s1 U2659 ( .Q(N9663), .DIN1(N9088), .DIN2(N9442) );
hi1s1 U2660 ( .Q(N9666), .DIN(N9089) );
nnd2s1 U2661 ( .Q(N9667), .DIN1(N9094), .DIN2(N9445) );
hi1s1 U2662 ( .Q(N9670), .DIN(N9095) );
or2s1 U2663 ( .Q(N9671), .DIN1(N8924), .DIN2(N8393) );
hi1s1 U2664 ( .Q(N9674), .DIN(N9117) );
hi1s1 U2665 ( .Q(N9675), .DIN(N8924) );
hi1s1 U2666 ( .Q(N9678), .DIN(N9127) );
or4s1 U2667 ( .Q(N9679), .DIN1(N4597), .DIN2(N8388), .DIN3(N8389), .DIN4(N9315) );
or2s1 U2668 ( .Q(N9682), .DIN1(N8931), .DIN2(N9318) );
or5s1 U2669 ( .Q(N9685), .DIN1(N4593), .DIN2(N8382), .DIN3(N8383), .DIN4(N8384), .DIN5(N9314) );
hi1s1 U2670 ( .Q(N9690), .DIN(N9146) );
nnd2s1 U2671 ( .Q(N9691), .DIN1(N9146), .DIN2(N8717) );
hi1s1 U2672 ( .Q(N9692), .DIN(N8931) );
hi1s1 U2673 ( .Q(N9695), .DIN(N9149) );
nnd2s1 U2674 ( .Q(N9698), .DIN1(N9401), .DIN2(N9400) );
nnd2s1 U2675 ( .Q(N9702), .DIN1(N9368), .DIN2(N9367) );
or2s1 U2676 ( .Q(N9707), .DIN1(N8996), .DIN2(N8517) );
hi1s1 U2677 ( .Q(N9710), .DIN(N9183) );
hi1s1 U2678 ( .Q(N9711), .DIN(N8996) );
hi1s1 U2679 ( .Q(N9714), .DIN(N9193) );
hi1s1 U2680 ( .Q(N9715), .DIN(N9203) );
nnd2s1 U2681 ( .Q(N9716), .DIN1(N9203), .DIN2(N6235) );
or2s1 U2682 ( .Q(N9717), .DIN1(N9005), .DIN2(N8518) );
hi1s1 U2683 ( .Q(N9720), .DIN(N9206) );
hi1s1 U2684 ( .Q(N9721), .DIN(N9220) );
nnd2s1 U2685 ( .Q(N9722), .DIN1(N9220), .DIN2(N7573) );
hi1s1 U2686 ( .Q(N9723), .DIN(N9005) );
hi1s1 U2687 ( .Q(N9726), .DIN(N9223) );
nnd2s1 U2688 ( .Q(N9727), .DIN1(N9418), .DIN2(N9417) );
and2s1 U2689 ( .Q(N9732), .DIN1(N9268), .DIN2(N8269) );
nnd2s1 U2690 ( .Q(N9733), .DIN1(N9581), .DIN2(N9326) );
and5s1 U2691 ( .Q(N9734), .DIN1(N89), .DIN2(N9408), .DIN3(N9332), .DIN4(N8394), .DIN5(N8421) );
and5s1 U2692 ( .Q(N9735), .DIN1(N89), .DIN2(N9408), .DIN3(N9332), .DIN4(N8394), .DIN5(N8421) );
and2s1 U2693 ( .Q(N9736), .DIN1(N9265), .DIN2(N8262) );
hi1s1 U2694 ( .Q(N9737), .DIN(N9555) );
hi1s1 U2695 ( .Q(N9738), .DIN(N9556) );
nnd2s1 U2696 ( .Q(N9739), .DIN1(N9361), .DIN2(N9601) );
nnd2s1 U2697 ( .Q(N9740), .DIN1(N9423), .DIN2(N1115) );
hi1s1 U2698 ( .Q(N9741), .DIN(N9423) );
nnd2s1 U2699 ( .Q(N9742), .DIN1(N9299), .DIN2(N9570) );
and2s1 U2700 ( .Q(N9754), .DIN1(N8333), .DIN2(N9280) );
or2s1 U2701 ( .Q(N9758), .DIN1(N8898), .DIN2(N9560) );
nnd2s1 U2702 ( .Q(N9762), .DIN1(N8660), .DIN2(N9561) );
nnd2s1 U2703 ( .Q(N9763), .DIN1(N8663), .DIN2(N9563) );
nnd2s1 U2704 ( .Q(N9764), .DIN1(N8666), .DIN2(N9565) );
nnd2s1 U2705 ( .Q(N9765), .DIN1(N8669), .DIN2(N9567) );
nnd2s1 U2706 ( .Q(N9766), .DIN1(N9297), .DIN2(N9569) );
and2s1 U2707 ( .Q(N9767), .DIN1(N9280), .DIN2(N367) );
nnd2s1 U2708 ( .Q(N9768), .DIN1(N9557), .DIN2(N9276) );
hi1s1 U2709 ( .Q(N9769), .DIN(N9307) );
nnd2s1 U2710 ( .Q(N9773), .DIN1(N9307), .DIN2(N367) );
nnd2s1 U2711 ( .Q(N9774), .DIN1(N9571), .DIN2(N9301) );
and2s1 U2712 ( .Q(N9775), .DIN1(N8365), .DIN2(N9307) );
or2s1 U2713 ( .Q(N9779), .DIN1(N8920), .DIN2(N9579) );
hi1s1 U2714 ( .Q(N9784), .DIN(N9478) );
nnd2s1 U2715 ( .Q(N9785), .DIN1(N9616), .DIN2(N9402) );
or2s1 U2716 ( .Q(N9786), .DIN1(N8950), .DIN2(N9585) );
and4s1 U2717 ( .Q(N9790), .DIN1(N89), .DIN2(N9408), .DIN3(N9332), .DIN4(N8394) );
or2s1 U2718 ( .Q(N9791), .DIN1(N8963), .DIN2(N9591) );
nnd2s1 U2719 ( .Q(N9795), .DIN1(N8735), .DIN2(N9592) );
nnd2s1 U2720 ( .Q(N9796), .DIN1(N8738), .DIN2(N9594) );
nnd2s1 U2721 ( .Q(N9797), .DIN1(N8741), .DIN2(N9596) );
nnd2s1 U2722 ( .Q(N9798), .DIN1(N8744), .DIN2(N9598) );
nnd2s1 U2723 ( .Q(N9799), .DIN1(N9359), .DIN2(N9600) );
nor2s1 U2724 ( .Q(N9800), .DIN1(N9602), .DIN2(N9369) );
nor2s1 U2725 ( .Q(N9801), .DIN1(N9603), .DIN2(N9370) );
nor2s1 U2726 ( .Q(N9802), .DIN1(N9604), .DIN2(N9371) );
nor2s1 U2727 ( .Q(N9803), .DIN1(N9605), .DIN2(N9372) );
hi1s1 U2728 ( .Q(N9805), .DIN(N9485) );
hi1s1 U2729 ( .Q(N9806), .DIN(N9488) );
or2s1 U2730 ( .Q(N9809), .DIN1(N8995), .DIN2(N9611) );
nor2s1 U2731 ( .Q(N9813), .DIN1(N9612), .DIN2(N9396) );
nor2s1 U2732 ( .Q(N9814), .DIN1(N9613), .DIN2(N9397) );
nor2s1 U2733 ( .Q(N9815), .DIN1(N9614), .DIN2(N9398) );
nor2s1 U2734 ( .Q(N9816), .DIN1(N9615), .DIN2(N9399) );
and2s1 U2735 ( .Q(N9817), .DIN1(N9617), .DIN2(N9407) );
or2s1 U2736 ( .Q(N9820), .DIN1(N9029), .DIN2(N9618) );
hi1s1 U2737 ( .Q(N9825), .DIN(N9517) );
hi1s1 U2738 ( .Q(N9826), .DIN(N9520) );
nor2s1 U2739 ( .Q(N9827), .DIN1(N9621), .DIN2(N9419) );
nor2s1 U2740 ( .Q(N9828), .DIN1(N9622), .DIN2(N9420) );
nor2s1 U2741 ( .Q(N9829), .DIN1(N9623), .DIN2(N9421) );
nor2s1 U2742 ( .Q(N9830), .DIN1(N9624), .DIN2(N9422) );
hi1s1 U2743 ( .Q(N9835), .DIN(N9426) );
nnd2s1 U2744 ( .Q(N9836), .DIN1(N9426), .DIN2(N4789) );
hi1s1 U2745 ( .Q(N9837), .DIN(N9429) );
nnd2s1 U2746 ( .Q(N9838), .DIN1(N9429), .DIN2(N4794) );
nnd2s1 U2747 ( .Q(N9846), .DIN1(N3625), .DIN2(N9659) );
nnd2s1 U2748 ( .Q(N9847), .DIN1(N4810), .DIN2(N9661) );
hi1s1 U2749 ( .Q(N9862), .DIN(N9462) );
nnd2s1 U2750 ( .Q(N9863), .DIN1(N7553), .DIN2(N9690) );
hi1s1 U2751 ( .Q(N9866), .DIN(N9473) );
nnd2s1 U2752 ( .Q(N9873), .DIN1(N5030), .DIN2(N9715) );
nnd2s1 U2753 ( .Q(N9876), .DIN1(N6236), .DIN2(N9721) );
nnd2s1 U2754 ( .Q(N9890), .DIN1(N9795), .DIN2(N9593) );
nnd2s1 U2755 ( .Q(N9891), .DIN1(N9797), .DIN2(N9597) );
hi1s1 U2756 ( .Q(N9892), .DIN(N9799) );
nnd2s1 U2757 ( .Q(N9893), .DIN1(N871), .DIN2(N9741) );
nnd2s1 U2758 ( .Q(N9894), .DIN1(N9762), .DIN2(N9562) );
nnd2s1 U2759 ( .Q(N9895), .DIN1(N9764), .DIN2(N9566) );
hi1s1 U2760 ( .Q(N9896), .DIN(N9766) );
hi1s1 U2761 ( .Q(N9897), .DIN(N9626) );
nnd2s1 U2762 ( .Q(N9898), .DIN1(N9626), .DIN2(N9249) );
hi1s1 U2763 ( .Q(N9899), .DIN(N9629) );
nnd2s1 U2764 ( .Q(N9900), .DIN1(N9629), .DIN2(N9250) );
hi1s1 U2765 ( .Q(N9901), .DIN(N9632) );
nnd2s1 U2766 ( .Q(N9902), .DIN1(N9632), .DIN2(N9251) );
hi1s1 U2767 ( .Q(N9903), .DIN(N9635) );
nnd2s1 U2768 ( .Q(N9904), .DIN1(N9635), .DIN2(N9252) );
hi1s1 U2769 ( .Q(N9905), .DIN(N9543) );
hi1s1 U2770 ( .Q(N9906), .DIN(N9650) );
nnd2s1 U2771 ( .Q(N9907), .DIN1(N9650), .DIN2(N5769) );
hi1s1 U2772 ( .Q(N9908), .DIN(N9653) );
nnd2s1 U2773 ( .Q(N9909), .DIN1(N9653), .DIN2(N5770) );
hi1s1 U2774 ( .Q(N9910), .DIN(N9656) );
nnd2s1 U2775 ( .Q(N9911), .DIN1(N9656), .DIN2(N9262) );
hi1s1 U2776 ( .Q(N9917), .DIN(N9551) );
nnd2s1 U2777 ( .Q(N9923), .DIN1(N9763), .DIN2(N9564) );
nnd2s1 U2778 ( .Q(N9924), .DIN1(N9765), .DIN2(N9568) );
or2s1 U2779 ( .Q(N9925), .DIN1(N8902), .DIN2(N9767) );
and2s1 U2780 ( .Q(N9932), .DIN1(N9575), .DIN2(N9773) );
and2s1 U2781 ( .Q(N9935), .DIN1(N9575), .DIN2(N9769) );
hi1s1 U2782 ( .Q(N9938), .DIN(N9698) );
nnd2s1 U2783 ( .Q(N9939), .DIN1(N9698), .DIN2(N9323) );
nnd2s1 U2784 ( .Q(N9945), .DIN1(N9796), .DIN2(N9595) );
nnd2s1 U2785 ( .Q(N9946), .DIN1(N9798), .DIN2(N9599) );
hi1s1 U2786 ( .Q(N9947), .DIN(N9702) );
nnd2s1 U2787 ( .Q(N9948), .DIN1(N9702), .DIN2(N6102) );
and2s1 U2788 ( .Q(N9949), .DIN1(N9608), .DIN2(N9375) );
hi1s1 U2789 ( .Q(N9953), .DIN(N9727) );
nnd2s1 U2790 ( .Q(N9954), .DIN1(N9727), .DIN2(N9412) );
nnd2s1 U2791 ( .Q(N9955), .DIN1(N3502), .DIN2(N9835) );
nnd2s1 U2792 ( .Q(N9956), .DIN1(N3510), .DIN2(N9837) );
hi1s1 U2793 ( .Q(N9957), .DIN(N9642) );
nnd2s1 U2794 ( .Q(N9958), .DIN1(N9642), .DIN2(N9645) );
hi1s1 U2795 ( .Q(N9959), .DIN(N9646) );
nnd2s1 U2796 ( .Q(N9960), .DIN1(N9646), .DIN2(N9649) );
nnd2s1 U2797 ( .Q(N9961), .DIN1(N9660), .DIN2(N9846) );
nnd2s1 U2798 ( .Q(N9964), .DIN1(N9662), .DIN2(N9847) );
hi1s1 U2799 ( .Q(N9967), .DIN(N9663) );
nnd2s1 U2800 ( .Q(N9968), .DIN1(N9663), .DIN2(N9666) );
hi1s1 U2801 ( .Q(N9969), .DIN(N9667) );
nnd2s1 U2802 ( .Q(N9970), .DIN1(N9667), .DIN2(N9670) );
hi1s1 U2803 ( .Q(N9971), .DIN(N9671) );
nnd2s1 U2804 ( .Q(N9972), .DIN1(N9671), .DIN2(N6213) );
hi1s1 U2805 ( .Q(N9973), .DIN(N9675) );
nnd2s1 U2806 ( .Q(N9974), .DIN1(N9675), .DIN2(N7551) );
hi1s1 U2807 ( .Q(N9975), .DIN(N9679) );
nnd2s1 U2808 ( .Q(N9976), .DIN1(N9679), .DIN2(N7552) );
hi1s1 U2809 ( .Q(N9977), .DIN(N9682) );
hi1s1 U2810 ( .Q(N9978), .DIN(N9685) );
nnd2s1 U2811 ( .Q(N9979), .DIN1(N9691), .DIN2(N9863) );
hi1s1 U2812 ( .Q(N9982), .DIN(N9692) );
nnd2s1 U2813 ( .Q(N9983), .DIN1(N9814), .DIN2(N9813) );
nnd2s1 U2814 ( .Q(N9986), .DIN1(N9816), .DIN2(N9815) );
nnd2s1 U2815 ( .Q(N9989), .DIN1(N9801), .DIN2(N9800) );
nnd2s1 U2816 ( .Q(N9992), .DIN1(N9803), .DIN2(N9802) );
hi1s1 U2817 ( .Q(N9995), .DIN(N9707) );
nnd2s1 U2818 ( .Q(N9996), .DIN1(N9707), .DIN2(N6231) );
hi1s1 U2819 ( .Q(N9997), .DIN(N9711) );
nnd2s1 U2820 ( .Q(N9998), .DIN1(N9711), .DIN2(N7572) );
nnd2s1 U2821 ( .Q(N9999), .DIN1(N9716), .DIN2(N9873) );
hi1s1 U2822 ( .Q(N10002), .DIN(N9717) );
nnd2s1 U2823 ( .Q(N10003), .DIN1(N9722), .DIN2(N9876) );
hi1s1 U2824 ( .Q(N10006), .DIN(N9723) );
nnd2s1 U2825 ( .Q(N10007), .DIN1(N9830), .DIN2(N9829) );
nnd2s1 U2826 ( .Q(N10010), .DIN1(N9828), .DIN2(N9827) );
and3s1 U2827 ( .Q(N10013), .DIN1(N9791), .DIN2(N8307), .DIN3(N8269) );
and4s1 U2828 ( .Q(N10014), .DIN1(N9758), .DIN2(N9344), .DIN3(N8307), .DIN4(N8269) );
and5s1 U2829 ( .Q(N10015), .DIN1(N367), .DIN2(N9754), .DIN3(N9344), .DIN4(N8307), .DIN5(N8269) );
and3s1 U2830 ( .Q(N10016), .DIN1(N9786), .DIN2(N8394), .DIN3(N8421) );
and4s1 U2831 ( .Q(N10017), .DIN1(N9820), .DIN2(N9332), .DIN3(N8394), .DIN4(N8421) );
and3s1 U2832 ( .Q(N10018), .DIN1(N9786), .DIN2(N8394), .DIN3(N8421) );
and4s1 U2833 ( .Q(N10019), .DIN1(N9820), .DIN2(N9332), .DIN3(N8394), .DIN4(N8421) );
and3s1 U2834 ( .Q(N10020), .DIN1(N9809), .DIN2(N8298), .DIN3(N8262) );
and4s1 U2835 ( .Q(N10021), .DIN1(N9779), .DIN2(N9385), .DIN3(N8298), .DIN4(N8262) );
and5s1 U2836 ( .Q(N10022), .DIN1(N367), .DIN2(N9775), .DIN3(N9385), .DIN4(N8298), .DIN5(N8262) );
hi1s1 U2837 ( .Q(N10023), .DIN(N9945) );
hi1s1 U2838 ( .Q(N10024), .DIN(N9946) );
nnd2s1 U2839 ( .Q(N10025), .DIN1(N9740), .DIN2(N9893) );
hi1s1 U2840 ( .Q(N10026), .DIN(N9923) );
hi1s1 U2841 ( .Q(N10028), .DIN(N9924) );
nnd2s1 U2842 ( .Q(N10032), .DIN1(N8595), .DIN2(N9897) );
nnd2s1 U2843 ( .Q(N10033), .DIN1(N8598), .DIN2(N9899) );
nnd2s1 U2844 ( .Q(N10034), .DIN1(N8601), .DIN2(N9901) );
nnd2s1 U2845 ( .Q(N10035), .DIN1(N8604), .DIN2(N9903) );
nnd2s1 U2846 ( .Q(N10036), .DIN1(N4803), .DIN2(N9906) );
nnd2s1 U2847 ( .Q(N10037), .DIN1(N4806), .DIN2(N9908) );
nnd2s1 U2848 ( .Q(N10038), .DIN1(N8627), .DIN2(N9910) );
and2s1 U2849 ( .Q(N10039), .DIN1(N9809), .DIN2(N8298) );
and3s1 U2850 ( .Q(N10040), .DIN1(N9779), .DIN2(N9385), .DIN3(N8298) );
and4s1 U2851 ( .Q(N10041), .DIN1(N367), .DIN2(N9775), .DIN3(N9385), .DIN4(N8298) );
and2s1 U2852 ( .Q(N10042), .DIN1(N9779), .DIN2(N9385) );
and3s1 U2853 ( .Q(N10043), .DIN1(N367), .DIN2(N9775), .DIN3(N9385) );
nnd2s1 U2854 ( .Q(N10050), .DIN1(N8727), .DIN2(N9938) );
hi1s1 U2855 ( .Q(N10053), .DIN(N9817) );
and2s1 U2856 ( .Q(N10054), .DIN1(N9817), .DIN2(N9029) );
and2s1 U2857 ( .Q(N10055), .DIN1(N9786), .DIN2(N8394) );
and3s1 U2858 ( .Q(N10056), .DIN1(N9820), .DIN2(N9332), .DIN3(N8394) );
and2s1 U2859 ( .Q(N10057), .DIN1(N9791), .DIN2(N8307) );
and3s1 U2860 ( .Q(N10058), .DIN1(N9758), .DIN2(N9344), .DIN3(N8307) );
and4s1 U2861 ( .Q(N10059), .DIN1(N367), .DIN2(N9754), .DIN3(N9344), .DIN4(N8307) );
and2s1 U2862 ( .Q(N10060), .DIN1(N9758), .DIN2(N9344) );
and3s1 U2863 ( .Q(N10061), .DIN1(N367), .DIN2(N9754), .DIN3(N9344) );
nnd2s1 U2864 ( .Q(N10062), .DIN1(N4997), .DIN2(N9947) );
nnd2s1 U2865 ( .Q(N10067), .DIN1(N8811), .DIN2(N9953) );
nnd2s1 U2866 ( .Q(N10070), .DIN1(N9955), .DIN2(N9836) );
nnd2s1 U2867 ( .Q(N10073), .DIN1(N9956), .DIN2(N9838) );
nnd2s1 U2868 ( .Q(N10076), .DIN1(N9068), .DIN2(N9957) );
nnd2s1 U2869 ( .Q(N10077), .DIN1(N9074), .DIN2(N9959) );
nnd2s1 U2870 ( .Q(N10082), .DIN1(N9089), .DIN2(N9967) );
nnd2s1 U2871 ( .Q(N10083), .DIN1(N9095), .DIN2(N9969) );
nnd2s1 U2872 ( .Q(N10084), .DIN1(N4871), .DIN2(N9971) );
nnd2s1 U2873 ( .Q(N10085), .DIN1(N6214), .DIN2(N9973) );
nnd2s1 U2874 ( .Q(N10086), .DIN1(N6217), .DIN2(N9975) );
nnd2s1 U2875 ( .Q(N10093), .DIN1(N5027), .DIN2(N9995) );
nnd2s1 U2876 ( .Q(N10094), .DIN1(N6232), .DIN2(N9997) );
or5s1 U2877 ( .Q(N10101), .DIN1(N9238), .DIN2(N9732), .DIN3(N10013), .DIN4(N10014), .DIN5(N10015) );
or5s1 U2878 ( .Q(N10102), .DIN1(N9339), .DIN2(N9526), .DIN3(N10016), .DIN4(N10017), .DIN5(N9734) );
or5s1 U2879 ( .Q(N10103), .DIN1(N9339), .DIN2(N9531), .DIN3(N10018), .DIN4(N10019), .DIN5(N9735) );
or5s1 U2880 ( .Q(N10104), .DIN1(N9242), .DIN2(N9736), .DIN3(N10020), .DIN4(N10021), .DIN5(N10022) );
and2s1 U2881 ( .Q(N10105), .DIN1(N9925), .DIN2(N9894) );
and2s1 U2882 ( .Q(N10106), .DIN1(N9925), .DIN2(N9895) );
and2s1 U2883 ( .Q(N10107), .DIN1(N9925), .DIN2(N9896) );
and2s1 U2884 ( .Q(N10108), .DIN1(N9925), .DIN2(N8253) );
nnd2s1 U2885 ( .Q(N10109), .DIN1(N10032), .DIN2(N9898) );
nnd2s1 U2886 ( .Q(N10110), .DIN1(N10033), .DIN2(N9900) );
nnd2s1 U2887 ( .Q(N10111), .DIN1(N10034), .DIN2(N9902) );
nnd2s1 U2888 ( .Q(N10112), .DIN1(N10035), .DIN2(N9904) );
nnd2s1 U2889 ( .Q(N10113), .DIN1(N10036), .DIN2(N9907) );
nnd2s1 U2890 ( .Q(N10114), .DIN1(N10037), .DIN2(N9909) );
nnd2s1 U2891 ( .Q(N10115), .DIN1(N10038), .DIN2(N9911) );
or4s1 U2892 ( .Q(N10116), .DIN1(N9265), .DIN2(N10039), .DIN3(N10040), .DIN4(N10041) );
or3s1 U2893 ( .Q(N10119), .DIN1(N9809), .DIN2(N10042), .DIN3(N10043) );
hi1s1 U2894 ( .Q(N10124), .DIN(N9925) );
and2s1 U2895 ( .Q(N10130), .DIN1(N9768), .DIN2(N9925) );
hi1s1 U2896 ( .Q(N10131), .DIN(N9932) );
hi1s1 U2897 ( .Q(N10132), .DIN(N9935) );
and2s1 U2898 ( .Q(N10133), .DIN1(N9932), .DIN2(N8920) );
nnd2s1 U2899 ( .Q(N10134), .DIN1(N10050), .DIN2(N9939) );
hi1s1 U2900 ( .Q(N10135), .DIN(N9983) );
nnd2s1 U2901 ( .Q(N10136), .DIN1(N9983), .DIN2(N9324) );
hi1s1 U2902 ( .Q(N10137), .DIN(N9986) );
nnd2s1 U2903 ( .Q(N10138), .DIN1(N9986), .DIN2(N9784) );
and2s1 U2904 ( .Q(N10139), .DIN1(N9785), .DIN2(N10053) );
or4s1 U2905 ( .Q(N10140), .DIN1(N8943), .DIN2(N10055), .DIN3(N10056), .DIN4(N9790) );
or4s1 U2906 ( .Q(N10141), .DIN1(N9268), .DIN2(N10057), .DIN3(N10058), .DIN4(N10059) );
or3s1 U2907 ( .Q(N10148), .DIN1(N9791), .DIN2(N10060), .DIN3(N10061) );
nnd2s1 U2908 ( .Q(N10155), .DIN1(N10062), .DIN2(N9948) );
hi1s1 U2909 ( .Q(N10156), .DIN(N9989) );
nnd2s1 U2910 ( .Q(N10157), .DIN1(N9989), .DIN2(N9805) );
hi1s1 U2911 ( .Q(N10158), .DIN(N9992) );
nnd2s1 U2912 ( .Q(N10159), .DIN1(N9992), .DIN2(N9806) );
hi1s1 U2913 ( .Q(N10160), .DIN(N9949) );
nnd2s1 U2914 ( .Q(N10161), .DIN1(N10067), .DIN2(N9954) );
hi1s1 U2915 ( .Q(N10162), .DIN(N10007) );
nnd2s1 U2916 ( .Q(N10163), .DIN1(N10007), .DIN2(N9825) );
hi1s1 U2917 ( .Q(N10164), .DIN(N10010) );
nnd2s1 U2918 ( .Q(N10165), .DIN1(N10010), .DIN2(N9826) );
nnd2s1 U2919 ( .Q(N10170), .DIN1(N10076), .DIN2(N9958) );
nnd2s1 U2920 ( .Q(N10173), .DIN1(N10077), .DIN2(N9960) );
hi1s1 U2921 ( .Q(N10176), .DIN(N9961) );
nnd2s1 U2922 ( .Q(N10177), .DIN1(N9961), .DIN2(N9082) );
hi1s1 U2923 ( .Q(N10178), .DIN(N9964) );
nnd2s1 U2924 ( .Q(N10179), .DIN1(N9964), .DIN2(N9086) );
nnd2s1 U2925 ( .Q(N10180), .DIN1(N10082), .DIN2(N9968) );
nnd2s1 U2926 ( .Q(N10183), .DIN1(N10083), .DIN2(N9970) );
nnd2s1 U2927 ( .Q(N10186), .DIN1(N9972), .DIN2(N10084) );
nnd2s1 U2928 ( .Q(N10189), .DIN1(N9974), .DIN2(N10085) );
nnd2s1 U2929 ( .Q(N10192), .DIN1(N9976), .DIN2(N10086) );
hi1s1 U2930 ( .Q(N10195), .DIN(N9979) );
nnd2s1 U2931 ( .Q(N10196), .DIN1(N9979), .DIN2(N9982) );
nnd2s1 U2932 ( .Q(N10197), .DIN1(N9996), .DIN2(N10093) );
nnd2s1 U2933 ( .Q(N10200), .DIN1(N9998), .DIN2(N10094) );
hi1s1 U2934 ( .Q(N10203), .DIN(N9999) );
nnd2s1 U2935 ( .Q(N10204), .DIN1(N9999), .DIN2(N10002) );
hi1s1 U2936 ( .Q(N10205), .DIN(N10003) );
nnd2s1 U2937 ( .Q(N10206), .DIN1(N10003), .DIN2(N10006) );
nnd2s1 U2938 ( .Q(N10212), .DIN1(N10070), .DIN2(N4308) );
nnd2s1 U2939 ( .Q(N10213), .DIN1(N10073), .DIN2(N4313) );
and2s1 U2940 ( .Q(N10230), .DIN1(N9774), .DIN2(N10131) );
nnd2s1 U2941 ( .Q(N10231), .DIN1(N8730), .DIN2(N10135) );
nnd2s1 U2942 ( .Q(N10232), .DIN1(N9478), .DIN2(N10137) );
or2s1 U2943 ( .Q(N10233), .DIN1(N10139), .DIN2(N10054) );
nnd2s1 U2944 ( .Q(N10234), .DIN1(N7100), .DIN2(N10140) );
nnd2s1 U2945 ( .Q(N10237), .DIN1(N9485), .DIN2(N10156) );
nnd2s1 U2946 ( .Q(N10238), .DIN1(N9488), .DIN2(N10158) );
nnd2s1 U2947 ( .Q(N10239), .DIN1(N9517), .DIN2(N10162) );
nnd2s1 U2948 ( .Q(N10240), .DIN1(N9520), .DIN2(N10164) );
hi1s1 U2949 ( .Q(N10241), .DIN(N10070) );
hi1s1 U2950 ( .Q(N10242), .DIN(N10073) );
nnd2s1 U2951 ( .Q(N10247), .DIN1(N8146), .DIN2(N10176) );
nnd2s1 U2952 ( .Q(N10248), .DIN1(N8156), .DIN2(N10178) );
nnd2s1 U2953 ( .Q(N10259), .DIN1(N9692), .DIN2(N10195) );
nnd2s1 U2954 ( .Q(N10264), .DIN1(N9717), .DIN2(N10203) );
nnd2s1 U2955 ( .Q(N10265), .DIN1(N9723), .DIN2(N10205) );
and2s1 U2956 ( .Q(N10266), .DIN1(N10026), .DIN2(N10124) );
and2s1 U2957 ( .Q(N10267), .DIN1(N10028), .DIN2(N10124) );
and2s1 U2958 ( .Q(N10268), .DIN1(N9742), .DIN2(N10124) );
and2s1 U2959 ( .Q(N10269), .DIN1(N6923), .DIN2(N10124) );
nnd2s1 U2960 ( .Q(N10270), .DIN1(N6762), .DIN2(N10116) );
nnd2s1 U2961 ( .Q(N10271), .DIN1(N3061), .DIN2(N10241) );
nnd2s1 U2962 ( .Q(N10272), .DIN1(N3064), .DIN2(N10242) );
nb1s1 U2963 ( .Q(N10273), .DIN(N10116) );
and5s1 U2964 ( .Q(N10278), .DIN1(N10141), .DIN2(N5728), .DIN3(N5707), .DIN4(N5718), .DIN5(N5697) );
and4s1 U2965 ( .Q(N10279), .DIN1(N10141), .DIN2(N5728), .DIN3(N5707), .DIN4(N5718) );
and3s1 U2966 ( .Q(N10280), .DIN1(N10141), .DIN2(N5728), .DIN3(N5718) );
and2s1 U2967 ( .Q(N10281), .DIN1(N10141), .DIN2(N5728) );
and2s1 U2968 ( .Q(N10282), .DIN1(N6784), .DIN2(N10141) );
hi1s1 U2969 ( .Q(N10283), .DIN(N10119) );
and5s1 U2970 ( .Q(N10287), .DIN1(N10148), .DIN2(N5936), .DIN3(N5915), .DIN4(N5926), .DIN5(N5905) );
and4s1 U2971 ( .Q(N10288), .DIN1(N10148), .DIN2(N5936), .DIN3(N5915), .DIN4(N5926) );
and3s1 U2972 ( .Q(N10289), .DIN1(N10148), .DIN2(N5936), .DIN3(N5926) );
and2s1 U2973 ( .Q(N10290), .DIN1(N10148), .DIN2(N5936) );
and2s1 U2974 ( .Q(N10291), .DIN1(N6881), .DIN2(N10148) );
and2s1 U2975 ( .Q(N10292), .DIN1(N8898), .DIN2(N10124) );
nnd2s1 U2976 ( .Q(N10293), .DIN1(N10231), .DIN2(N10136) );
nnd2s1 U2977 ( .Q(N10294), .DIN1(N10232), .DIN2(N10138) );
nnd2s1 U2978 ( .Q(N10295), .DIN1(N8412), .DIN2(N10233) );
and2s1 U2979 ( .Q(N10296), .DIN1(N8959), .DIN2(N10234) );
nnd2s1 U2980 ( .Q(N10299), .DIN1(N10237), .DIN2(N10157) );
nnd2s1 U2981 ( .Q(N10300), .DIN1(N10238), .DIN2(N10159) );
or2s1 U2982 ( .Q(N10301), .DIN1(N10230), .DIN2(N10133) );
nnd2s1 U2983 ( .Q(N10306), .DIN1(N10239), .DIN2(N10163) );
nnd2s1 U2984 ( .Q(N10307), .DIN1(N10240), .DIN2(N10165) );
nb1s1 U2985 ( .Q(N10308), .DIN(N10148) );
nb1s1 U2986 ( .Q(N10311), .DIN(N10141) );
hi1s1 U2987 ( .Q(N10314), .DIN(N10170) );
nnd2s1 U2988 ( .Q(N10315), .DIN1(N10170), .DIN2(N9071) );
hi1s1 U2989 ( .Q(N10316), .DIN(N10173) );
nnd2s1 U2990 ( .Q(N10317), .DIN1(N10173), .DIN2(N9077) );
nnd2s1 U2991 ( .Q(N10318), .DIN1(N10247), .DIN2(N10177) );
nnd2s1 U2992 ( .Q(N10321), .DIN1(N10248), .DIN2(N10179) );
hi1s1 U2993 ( .Q(N10324), .DIN(N10180) );
nnd2s1 U2994 ( .Q(N10325), .DIN1(N10180), .DIN2(N9092) );
hi1s1 U2995 ( .Q(N10326), .DIN(N10183) );
nnd2s1 U2996 ( .Q(N10327), .DIN1(N10183), .DIN2(N9098) );
hi1s1 U2997 ( .Q(N10328), .DIN(N10186) );
nnd2s1 U2998 ( .Q(N10329), .DIN1(N10186), .DIN2(N9674) );
hi1s1 U2999 ( .Q(N10330), .DIN(N10189) );
nnd2s1 U3000 ( .Q(N10331), .DIN1(N10189), .DIN2(N9678) );
hi1s1 U3001 ( .Q(N10332), .DIN(N10192) );
nnd2s1 U3002 ( .Q(N10333), .DIN1(N10192), .DIN2(N9977) );
nnd2s1 U3003 ( .Q(N10334), .DIN1(N10259), .DIN2(N10196) );
hi1s1 U3004 ( .Q(N10337), .DIN(N10197) );
nnd2s1 U3005 ( .Q(N10338), .DIN1(N10197), .DIN2(N9710) );
hi1s1 U3006 ( .Q(N10339), .DIN(N10200) );
nnd2s1 U3007 ( .Q(N10340), .DIN1(N10200), .DIN2(N9714) );
nnd2s1 U3008 ( .Q(N10341), .DIN1(N10264), .DIN2(N10204) );
nnd2s1 U3009 ( .Q(N10344), .DIN1(N10265), .DIN2(N10206) );
or2s1 U3010 ( .Q(N10350), .DIN1(N10266), .DIN2(N10105) );
or2s1 U3011 ( .Q(N10351), .DIN1(N10267), .DIN2(N10106) );
or2s1 U3012 ( .Q(N10352), .DIN1(N10268), .DIN2(N10107) );
or2s1 U3013 ( .Q(N10353), .DIN1(N10269), .DIN2(N10108) );
and2s1 U3014 ( .Q(N10354), .DIN1(N8857), .DIN2(N10270) );
nnd2s1 U3015 ( .Q(N10357), .DIN1(N10271), .DIN2(N10212) );
nnd2s1 U3016 ( .Q(N10360), .DIN1(N10272), .DIN2(N10213) );
or2s1 U3017 ( .Q(N10367), .DIN1(N7620), .DIN2(N10282) );
or2s1 U3018 ( .Q(N10375), .DIN1(N7671), .DIN2(N10291) );
or2s1 U3019 ( .Q(N10381), .DIN1(N10292), .DIN2(N10130) );
and4s1 U3020 ( .Q(N10388), .DIN1(N10114), .DIN2(N10134), .DIN3(N10293), .DIN4(N10294) );
and2s1 U3021 ( .Q(N10391), .DIN1(N9582), .DIN2(N10295) );
and4s1 U3022 ( .Q(N10399), .DIN1(N10113), .DIN2(N10115), .DIN3(N10299), .DIN4(N10300) );
and4s1 U3023 ( .Q(N10402), .DIN1(N10155), .DIN2(N10161), .DIN3(N10306), .DIN4(N10307) );
or5s1 U3024 ( .Q(N10406), .DIN1(N3229), .DIN2(N6888), .DIN3(N6889), .DIN4(N6890), .DIN5(N10287) );
or4s1 U3025 ( .Q(N10409), .DIN1(N3232), .DIN2(N6891), .DIN3(N6892), .DIN4(N10288) );
or3s1 U3026 ( .Q(N10412), .DIN1(N3236), .DIN2(N6893), .DIN3(N10289) );
or2s1 U3027 ( .Q(N10415), .DIN1(N3241), .DIN2(N10290) );
or5s1 U3028 ( .Q(N10419), .DIN1(N3137), .DIN2(N6791), .DIN3(N6792), .DIN4(N6793), .DIN5(N10278) );
or4s1 U3029 ( .Q(N10422), .DIN1(N3140), .DIN2(N6794), .DIN3(N6795), .DIN4(N10279) );
or3s1 U3030 ( .Q(N10425), .DIN1(N3144), .DIN2(N6796), .DIN3(N10280) );
or2s1 U3031 ( .Q(N10428), .DIN1(N3149), .DIN2(N10281) );
nnd2s1 U3032 ( .Q(N10431), .DIN1(N8117), .DIN2(N10314) );
nnd2s1 U3033 ( .Q(N10432), .DIN1(N8134), .DIN2(N10316) );
nnd2s1 U3034 ( .Q(N10437), .DIN1(N8169), .DIN2(N10324) );
nnd2s1 U3035 ( .Q(N10438), .DIN1(N8186), .DIN2(N10326) );
nnd2s1 U3036 ( .Q(N10439), .DIN1(N9117), .DIN2(N10328) );
nnd2s1 U3037 ( .Q(N10440), .DIN1(N9127), .DIN2(N10330) );
nnd2s1 U3038 ( .Q(N10441), .DIN1(N9682), .DIN2(N10332) );
nnd2s1 U3039 ( .Q(N10444), .DIN1(N9183), .DIN2(N10337) );
nnd2s1 U3040 ( .Q(N10445), .DIN1(N9193), .DIN2(N10339) );
hi1s1 U3041 ( .Q(N10450), .DIN(N10296) );
and2s1 U3042 ( .Q(N10451), .DIN1(N10296), .DIN2(N4193) );
hi1s1 U3043 ( .Q(N10455), .DIN(N10308) );
nnd2s1 U3044 ( .Q(N10456), .DIN1(N10308), .DIN2(N8242) );
hi1s1 U3045 ( .Q(N10465), .DIN(N10311) );
nnd2s1 U3046 ( .Q(N10466), .DIN1(N10311), .DIN2(N8247) );
hi1s1 U3047 ( .Q(N10479), .DIN(N10273) );
hi1s1 U3048 ( .Q(N10497), .DIN(N10301) );
nnd2s1 U3049 ( .Q(N10509), .DIN1(N10431), .DIN2(N10315) );
nnd2s1 U3050 ( .Q(N10512), .DIN1(N10432), .DIN2(N10317) );
hi1s1 U3051 ( .Q(N10515), .DIN(N10318) );
nnd2s1 U3052 ( .Q(N10516), .DIN1(N10318), .DIN2(N8632) );
hi1s1 U3053 ( .Q(N10517), .DIN(N10321) );
nnd2s1 U3054 ( .Q(N10518), .DIN1(N10321), .DIN2(N8637) );
nnd2s1 U3055 ( .Q(N10519), .DIN1(N10437), .DIN2(N10325) );
nnd2s1 U3056 ( .Q(N10522), .DIN1(N10438), .DIN2(N10327) );
nnd2s1 U3057 ( .Q(N10525), .DIN1(N10439), .DIN2(N10329) );
nnd2s1 U3058 ( .Q(N10528), .DIN1(N10440), .DIN2(N10331) );
nnd2s1 U3059 ( .Q(N10531), .DIN1(N10441), .DIN2(N10333) );
hi1s1 U3060 ( .Q(N10534), .DIN(N10334) );
nnd2s1 U3061 ( .Q(N10535), .DIN1(N10334), .DIN2(N9695) );
nnd2s1 U3062 ( .Q(N10536), .DIN1(N10444), .DIN2(N10338) );
nnd2s1 U3063 ( .Q(N10539), .DIN1(N10445), .DIN2(N10340) );
hi1s1 U3064 ( .Q(N10542), .DIN(N10341) );
nnd2s1 U3065 ( .Q(N10543), .DIN1(N10341), .DIN2(N9720) );
hi1s1 U3066 ( .Q(N10544), .DIN(N10344) );
nnd2s1 U3067 ( .Q(N10545), .DIN1(N10344), .DIN2(N9726) );
and2s1 U3068 ( .Q(N10546), .DIN1(N5631), .DIN2(N10450) );
hi1s1 U3069 ( .Q(N10547), .DIN(N10391) );
and2s1 U3070 ( .Q(N10548), .DIN1(N10391), .DIN2(N8950) );
and2s1 U3071 ( .Q(N10549), .DIN1(N5165), .DIN2(N10367) );
hi1s1 U3072 ( .Q(N10550), .DIN(N10354) );
and2s1 U3073 ( .Q(N10551), .DIN1(N10354), .DIN2(N3126) );
nnd2s1 U3074 ( .Q(N10552), .DIN1(N7411), .DIN2(N10455) );
and2s1 U3075 ( .Q(N10553), .DIN1(N10375), .DIN2(N9539) );
and2s1 U3076 ( .Q(N10554), .DIN1(N10375), .DIN2(N9540) );
and2s1 U3077 ( .Q(N10555), .DIN1(N10375), .DIN2(N9541) );
and2s1 U3078 ( .Q(N10556), .DIN1(N10375), .DIN2(N6761) );
hi1s1 U3079 ( .Q(N10557), .DIN(N10406) );
nnd2s1 U3080 ( .Q(N10558), .DIN1(N10406), .DIN2(N8243) );
hi1s1 U3081 ( .Q(N10559), .DIN(N10409) );
nnd2s1 U3082 ( .Q(N10560), .DIN1(N10409), .DIN2(N8244) );
hi1s1 U3083 ( .Q(N10561), .DIN(N10412) );
nnd2s1 U3084 ( .Q(N10562), .DIN1(N10412), .DIN2(N8245) );
hi1s1 U3085 ( .Q(N10563), .DIN(N10415) );
nnd2s1 U3086 ( .Q(N10564), .DIN1(N10415), .DIN2(N8246) );
nnd2s1 U3087 ( .Q(N10565), .DIN1(N7426), .DIN2(N10465) );
hi1s1 U3088 ( .Q(N10566), .DIN(N10419) );
nnd2s1 U3089 ( .Q(N10567), .DIN1(N10419), .DIN2(N8248) );
hi1s1 U3090 ( .Q(N10568), .DIN(N10422) );
nnd2s1 U3091 ( .Q(N10569), .DIN1(N10422), .DIN2(N8249) );
hi1s1 U3092 ( .Q(N10570), .DIN(N10425) );
nnd2s1 U3093 ( .Q(N10571), .DIN1(N10425), .DIN2(N8250) );
hi1s1 U3094 ( .Q(N10572), .DIN(N10428) );
nnd2s1 U3095 ( .Q(N10573), .DIN1(N10428), .DIN2(N8251) );
hi1s1 U3096 ( .Q(N10574), .DIN(N10399) );
hi1s1 U3097 ( .Q(N10575), .DIN(N10402) );
hi1s1 U3098 ( .Q(N10576), .DIN(N10388) );
and3s1 U3099 ( .Q(N10577), .DIN1(N10399), .DIN2(N10402), .DIN3(N10388) );
and3s1 U3100 ( .Q(N10581), .DIN1(N10360), .DIN2(N9543), .DIN3(N10273) );
and3s1 U3101 ( .Q(N10582), .DIN1(N10357), .DIN2(N9905), .DIN3(N10273) );
hi1s1 U3102 ( .Q(N10583), .DIN(N10367) );
and2s1 U3103 ( .Q(N10587), .DIN1(N10367), .DIN2(N5735) );
and2s1 U3104 ( .Q(N10588), .DIN1(N10367), .DIN2(N3135) );
hi1s1 U3105 ( .Q(N10589), .DIN(N10375) );
and5s1 U3106 ( .Q(N10594), .DIN1(N10381), .DIN2(N7180), .DIN3(N7159), .DIN4(N7170), .DIN5(N7149) );
and4s1 U3107 ( .Q(N10595), .DIN1(N10381), .DIN2(N7180), .DIN3(N7159), .DIN4(N7170) );
and3s1 U3108 ( .Q(N10596), .DIN1(N10381), .DIN2(N7180), .DIN3(N7170) );
and2s1 U3109 ( .Q(N10597), .DIN1(N10381), .DIN2(N7180) );
and2s1 U3110 ( .Q(N10598), .DIN1(N8444), .DIN2(N10381) );
nb1s1 U3111 ( .Q(N10602), .DIN(N10381) );
nnd2s1 U3112 ( .Q(N10609), .DIN1(N7479), .DIN2(N10515) );
nnd2s1 U3113 ( .Q(N10610), .DIN1(N7491), .DIN2(N10517) );
nnd2s1 U3114 ( .Q(N10621), .DIN1(N9149), .DIN2(N10534) );
nnd2s1 U3115 ( .Q(N10626), .DIN1(N9206), .DIN2(N10542) );
nnd2s1 U3116 ( .Q(N10627), .DIN1(N9223), .DIN2(N10544) );
or2s1 U3117 ( .Q(N10628), .DIN1(N10546), .DIN2(N10451) );
and2s1 U3118 ( .Q(N10629), .DIN1(N9733), .DIN2(N10547) );
and2s1 U3119 ( .Q(N10631), .DIN1(N5166), .DIN2(N10550) );
nnd2s1 U3120 ( .Q(N10632), .DIN1(N10552), .DIN2(N10456) );
nnd2s1 U3121 ( .Q(N10637), .DIN1(N7414), .DIN2(N10557) );
nnd2s1 U3122 ( .Q(N10638), .DIN1(N7417), .DIN2(N10559) );
nnd2s1 U3123 ( .Q(N10639), .DIN1(N7420), .DIN2(N10561) );
nnd2s1 U3124 ( .Q(N10640), .DIN1(N7423), .DIN2(N10563) );
nnd2s1 U3125 ( .Q(N10641), .DIN1(N10565), .DIN2(N10466) );
nnd2s1 U3126 ( .Q(N10642), .DIN1(N7429), .DIN2(N10566) );
nnd2s1 U3127 ( .Q(N10643), .DIN1(N7432), .DIN2(N10568) );
nnd2s1 U3128 ( .Q(N10644), .DIN1(N7435), .DIN2(N10570) );
nnd2s1 U3129 ( .Q(N10645), .DIN1(N7438), .DIN2(N10572) );
and3s1 U3130 ( .Q(N10647), .DIN1(N886), .DIN2(N887), .DIN3(N10577) );
and3s1 U3131 ( .Q(N10648), .DIN1(N10360), .DIN2(N8857), .DIN3(N10479) );
and3s1 U3132 ( .Q(N10649), .DIN1(N10357), .DIN2(N7609), .DIN3(N10479) );
or2s1 U3133 ( .Q(N10652), .DIN1(N8966), .DIN2(N10598) );
or5s1 U3134 ( .Q(N10659), .DIN1(N4675), .DIN2(N8451), .DIN3(N8452), .DIN4(N8453), .DIN5(N10594) );
or4s1 U3135 ( .Q(N10662), .DIN1(N4678), .DIN2(N8454), .DIN3(N8455), .DIN4(N10595) );
or3s1 U3136 ( .Q(N10665), .DIN1(N4682), .DIN2(N8456), .DIN3(N10596) );
or2s1 U3137 ( .Q(N10668), .DIN1(N4687), .DIN2(N10597) );
hi1s1 U3138 ( .Q(N10671), .DIN(N10509) );
nnd2s1 U3139 ( .Q(N10672), .DIN1(N10509), .DIN2(N8615) );
hi1s1 U3140 ( .Q(N10673), .DIN(N10512) );
nnd2s1 U3141 ( .Q(N10674), .DIN1(N10512), .DIN2(N8624) );
nnd2s1 U3142 ( .Q(N10675), .DIN1(N10609), .DIN2(N10516) );
nnd2s1 U3143 ( .Q(N10678), .DIN1(N10610), .DIN2(N10518) );
hi1s1 U3144 ( .Q(N10681), .DIN(N10519) );
nnd2s1 U3145 ( .Q(N10682), .DIN1(N10519), .DIN2(N8644) );
hi1s1 U3146 ( .Q(N10683), .DIN(N10522) );
nnd2s1 U3147 ( .Q(N10684), .DIN1(N10522), .DIN2(N8653) );
hi1s1 U3148 ( .Q(N10685), .DIN(N10525) );
nnd2s1 U3149 ( .Q(N10686), .DIN1(N10525), .DIN2(N9454) );
hi1s1 U3150 ( .Q(N10687), .DIN(N10528) );
nnd2s1 U3151 ( .Q(N10688), .DIN1(N10528), .DIN2(N9459) );
hi1s1 U3152 ( .Q(N10689), .DIN(N10531) );
nnd2s1 U3153 ( .Q(N10690), .DIN1(N10531), .DIN2(N9978) );
nnd2s1 U3154 ( .Q(N10691), .DIN1(N10621), .DIN2(N10535) );
hi1s1 U3155 ( .Q(N10694), .DIN(N10536) );
nnd2s1 U3156 ( .Q(N10695), .DIN1(N10536), .DIN2(N9493) );
hi1s1 U3157 ( .Q(N10696), .DIN(N10539) );
nnd2s1 U3158 ( .Q(N10697), .DIN1(N10539), .DIN2(N9498) );
nnd2s1 U3159 ( .Q(N10698), .DIN1(N10626), .DIN2(N10543) );
nnd2s1 U3160 ( .Q(N10701), .DIN1(N10627), .DIN2(N10545) );
or2s1 U3161 ( .Q(N10704), .DIN1(N10629), .DIN2(N10548) );
and2s1 U3162 ( .Q(N10705), .DIN1(N3159), .DIN2(N10583) );
or2s1 U3163 ( .Q(N10706), .DIN1(N10631), .DIN2(N10551) );
and2s1 U3164 ( .Q(N10707), .DIN1(N9737), .DIN2(N10589) );
and2s1 U3165 ( .Q(N10708), .DIN1(N9738), .DIN2(N10589) );
and2s1 U3166 ( .Q(N10709), .DIN1(N9243), .DIN2(N10589) );
and2s1 U3167 ( .Q(N10710), .DIN1(N5892), .DIN2(N10589) );
nnd2s1 U3168 ( .Q(N10711), .DIN1(N10637), .DIN2(N10558) );
nnd2s1 U3169 ( .Q(N10712), .DIN1(N10638), .DIN2(N10560) );
nnd2s1 U3170 ( .Q(N10713), .DIN1(N10639), .DIN2(N10562) );
nnd2s1 U3171 ( .Q(N10714), .DIN1(N10640), .DIN2(N10564) );
nnd2s1 U3172 ( .Q(N10715), .DIN1(N10642), .DIN2(N10567) );
nnd2s1 U3173 ( .Q(N10716), .DIN1(N10643), .DIN2(N10569) );
nnd2s1 U3174 ( .Q(N10717), .DIN1(N10644), .DIN2(N10571) );
nnd2s1 U3175 ( .Q(N10718), .DIN1(N10645), .DIN2(N10573) );
hi1s1 U3176 ( .Q(N10719), .DIN(N10602) );
nnd2s1 U3177 ( .Q(N10720), .DIN1(N10602), .DIN2(N9244) );
hi1s1 U3178 ( .Q(N10729), .DIN(N10647) );
and2s1 U3179 ( .Q(N10730), .DIN1(N5178), .DIN2(N10583) );
and2s1 U3180 ( .Q(N10731), .DIN1(N2533), .DIN2(N10583) );
nnd2s1 U3181 ( .Q(N10737), .DIN1(N7447), .DIN2(N10671) );
nnd2s1 U3182 ( .Q(N10738), .DIN1(N7465), .DIN2(N10673) );
or4s1 U3183 ( .Q(N10739), .DIN1(N10648), .DIN2(N10649), .DIN3(N10581), .DIN4(N10582) );
nnd2s1 U3184 ( .Q(N10746), .DIN1(N7503), .DIN2(N10681) );
nnd2s1 U3185 ( .Q(N10747), .DIN1(N7521), .DIN2(N10683) );
nnd2s1 U3186 ( .Q(N10748), .DIN1(N8678), .DIN2(N10685) );
nnd2s1 U3187 ( .Q(N10749), .DIN1(N8690), .DIN2(N10687) );
nnd2s1 U3188 ( .Q(N10750), .DIN1(N9685), .DIN2(N10689) );
nnd2s1 U3189 ( .Q(N10753), .DIN1(N8757), .DIN2(N10694) );
nnd2s1 U3190 ( .Q(N10754), .DIN1(N8769), .DIN2(N10696) );
or2s1 U3191 ( .Q(N10759), .DIN1(N10705), .DIN2(N10549) );
or2s1 U3192 ( .Q(N10760), .DIN1(N10707), .DIN2(N10553) );
or2s1 U3193 ( .Q(N10761), .DIN1(N10708), .DIN2(N10554) );
or2s1 U3194 ( .Q(N10762), .DIN1(N10709), .DIN2(N10555) );
or2s1 U3195 ( .Q(N10763), .DIN1(N10710), .DIN2(N10556) );
nnd2s1 U3196 ( .Q(N10764), .DIN1(N8580), .DIN2(N10719) );
and2s1 U3197 ( .Q(N10765), .DIN1(N10652), .DIN2(N9890) );
and2s1 U3198 ( .Q(N10766), .DIN1(N10652), .DIN2(N9891) );
and2s1 U3199 ( .Q(N10767), .DIN1(N10652), .DIN2(N9892) );
and2s1 U3200 ( .Q(N10768), .DIN1(N10652), .DIN2(N8252) );
hi1s1 U3201 ( .Q(N10769), .DIN(N10659) );
nnd2s1 U3202 ( .Q(N10770), .DIN1(N10659), .DIN2(N9245) );
hi1s1 U3203 ( .Q(N10771), .DIN(N10662) );
nnd2s1 U3204 ( .Q(N10772), .DIN1(N10662), .DIN2(N9246) );
hi1s1 U3205 ( .Q(N10773), .DIN(N10665) );
nnd2s1 U3206 ( .Q(N10774), .DIN1(N10665), .DIN2(N9247) );
hi1s1 U3207 ( .Q(N10775), .DIN(N10668) );
nnd2s1 U3208 ( .Q(N10776), .DIN1(N10668), .DIN2(N9248) );
or2s1 U3209 ( .Q(N10778), .DIN1(N10730), .DIN2(N10587) );
or2s1 U3210 ( .Q(N10781), .DIN1(N10731), .DIN2(N10588) );
hi1s1 U3211 ( .Q(N10784), .DIN(N10652) );
nnd2s1 U3212 ( .Q(N10789), .DIN1(N10737), .DIN2(N10672) );
nnd2s1 U3213 ( .Q(N10792), .DIN1(N10738), .DIN2(N10674) );
hi1s1 U3214 ( .Q(N10796), .DIN(N10675) );
nnd2s1 U3215 ( .Q(N10797), .DIN1(N10675), .DIN2(N8633) );
hi1s1 U3216 ( .Q(N10798), .DIN(N10678) );
nnd2s1 U3217 ( .Q(N10799), .DIN1(N10678), .DIN2(N8638) );
nnd2s1 U3218 ( .Q(N10800), .DIN1(N10746), .DIN2(N10682) );
nnd2s1 U3219 ( .Q(N10803), .DIN1(N10747), .DIN2(N10684) );
nnd2s1 U3220 ( .Q(N10806), .DIN1(N10748), .DIN2(N10686) );
nnd2s1 U3221 ( .Q(N10809), .DIN1(N10749), .DIN2(N10688) );
nnd2s1 U3222 ( .Q(N10812), .DIN1(N10750), .DIN2(N10690) );
hi1s1 U3223 ( .Q(N10815), .DIN(N10691) );
nnd2s1 U3224 ( .Q(N10816), .DIN1(N10691), .DIN2(N9866) );
nnd2s1 U3225 ( .Q(N10817), .DIN1(N10753), .DIN2(N10695) );
nnd2s1 U3226 ( .Q(N10820), .DIN1(N10754), .DIN2(N10697) );
hi1s1 U3227 ( .Q(N10823), .DIN(N10698) );
nnd2s1 U3228 ( .Q(N10824), .DIN1(N10698), .DIN2(N9505) );
hi1s1 U3229 ( .Q(N10825), .DIN(N10701) );
nnd2s1 U3230 ( .Q(N10826), .DIN1(N10701), .DIN2(N9514) );
nnd2s1 U3231 ( .Q(N10827), .DIN1(N10764), .DIN2(N10720) );
nnd2s1 U3232 ( .Q(N10832), .DIN1(N8583), .DIN2(N10769) );
nnd2s1 U3233 ( .Q(N10833), .DIN1(N8586), .DIN2(N10771) );
nnd2s1 U3234 ( .Q(N10834), .DIN1(N8589), .DIN2(N10773) );
nnd2s1 U3235 ( .Q(N10835), .DIN1(N8592), .DIN2(N10775) );
hi1s1 U3236 ( .Q(N10836), .DIN(N10739) );
nb1s1 U3237 ( .Q(N10837), .DIN(N10778) );
nb1s1 U3238 ( .Q(N10838), .DIN(N10778) );
nb1s1 U3239 ( .Q(N10839), .DIN(N10781) );
nb1s1 U3240 ( .Q(N10840), .DIN(N10781) );
nnd2s1 U3241 ( .Q(N10845), .DIN1(N7482), .DIN2(N10796) );
nnd2s1 U3242 ( .Q(N10846), .DIN1(N7494), .DIN2(N10798) );
nnd2s1 U3243 ( .Q(N10857), .DIN1(N9473), .DIN2(N10815) );
nnd2s1 U3244 ( .Q(N10862), .DIN1(N8781), .DIN2(N10823) );
nnd2s1 U3245 ( .Q(N10863), .DIN1(N8799), .DIN2(N10825) );
and2s1 U3246 ( .Q(N10864), .DIN1(N10023), .DIN2(N10784) );
and2s1 U3247 ( .Q(N10865), .DIN1(N10024), .DIN2(N10784) );
and2s1 U3248 ( .Q(N10866), .DIN1(N9739), .DIN2(N10784) );
and2s1 U3249 ( .Q(N10867), .DIN1(N7136), .DIN2(N10784) );
nnd2s1 U3250 ( .Q(N10868), .DIN1(N10832), .DIN2(N10770) );
nnd2s1 U3251 ( .Q(N10869), .DIN1(N10833), .DIN2(N10772) );
nnd2s1 U3252 ( .Q(N10870), .DIN1(N10834), .DIN2(N10774) );
nnd2s1 U3253 ( .Q(N10871), .DIN1(N10835), .DIN2(N10776) );
hi1s1 U3254 ( .Q(N10872), .DIN(N10789) );
nnd2s1 U3255 ( .Q(N10873), .DIN1(N10789), .DIN2(N8616) );
hi1s1 U3256 ( .Q(N10874), .DIN(N10792) );
nnd2s1 U3257 ( .Q(N10875), .DIN1(N10792), .DIN2(N8625) );
nnd2s1 U3258 ( .Q(N10876), .DIN1(N10845), .DIN2(N10797) );
nnd2s1 U3259 ( .Q(N10879), .DIN1(N10846), .DIN2(N10799) );
hi1s1 U3260 ( .Q(N10882), .DIN(N10800) );
nnd2s1 U3261 ( .Q(N10883), .DIN1(N10800), .DIN2(N8645) );
hi1s1 U3262 ( .Q(N10884), .DIN(N10803) );
nnd2s1 U3263 ( .Q(N10885), .DIN1(N10803), .DIN2(N8654) );
hi1s1 U3264 ( .Q(N10886), .DIN(N10806) );
nnd2s1 U3265 ( .Q(N10887), .DIN1(N10806), .DIN2(N9455) );
hi1s1 U3266 ( .Q(N10888), .DIN(N10809) );
nnd2s1 U3267 ( .Q(N10889), .DIN1(N10809), .DIN2(N9460) );
hi1s1 U3268 ( .Q(N10890), .DIN(N10812) );
nnd2s1 U3269 ( .Q(N10891), .DIN1(N10812), .DIN2(N9862) );
nnd2s1 U3270 ( .Q(N10892), .DIN1(N10857), .DIN2(N10816) );
hi1s1 U3271 ( .Q(N10895), .DIN(N10817) );
nnd2s1 U3272 ( .Q(N10896), .DIN1(N10817), .DIN2(N9494) );
hi1s1 U3273 ( .Q(N10897), .DIN(N10820) );
nnd2s1 U3274 ( .Q(N10898), .DIN1(N10820), .DIN2(N9499) );
nnd2s1 U3275 ( .Q(N10899), .DIN1(N10862), .DIN2(N10824) );
nnd2s1 U3276 ( .Q(N10902), .DIN1(N10863), .DIN2(N10826) );
or2s1 U3277 ( .Q(N10905), .DIN1(N10864), .DIN2(N10765) );
or2s1 U3278 ( .Q(N10906), .DIN1(N10865), .DIN2(N10766) );
or2s1 U3279 ( .Q(N10907), .DIN1(N10866), .DIN2(N10767) );
or2s1 U3280 ( .Q(N10908), .DIN1(N10867), .DIN2(N10768) );
nnd2s1 U3281 ( .Q(N10909), .DIN1(N7450), .DIN2(N10872) );
nnd2s1 U3282 ( .Q(N10910), .DIN1(N7468), .DIN2(N10874) );
nnd2s1 U3283 ( .Q(N10915), .DIN1(N7506), .DIN2(N10882) );
nnd2s1 U3284 ( .Q(N10916), .DIN1(N7524), .DIN2(N10884) );
nnd2s1 U3285 ( .Q(N10917), .DIN1(N8681), .DIN2(N10886) );
nnd2s1 U3286 ( .Q(N10918), .DIN1(N8693), .DIN2(N10888) );
nnd2s1 U3287 ( .Q(N10919), .DIN1(N9462), .DIN2(N10890) );
nnd2s1 U3288 ( .Q(N10922), .DIN1(N8760), .DIN2(N10895) );
nnd2s1 U3289 ( .Q(N10923), .DIN1(N8772), .DIN2(N10897) );
nnd2s1 U3290 ( .Q(N10928), .DIN1(N10909), .DIN2(N10873) );
nnd2s1 U3291 ( .Q(N10931), .DIN1(N10910), .DIN2(N10875) );
hi1s1 U3292 ( .Q(N10934), .DIN(N10876) );
nnd2s1 U3293 ( .Q(N10935), .DIN1(N10876), .DIN2(N8634) );
hi1s1 U3294 ( .Q(N10936), .DIN(N10879) );
nnd2s1 U3295 ( .Q(N10937), .DIN1(N10879), .DIN2(N8639) );
nnd2s1 U3296 ( .Q(N10938), .DIN1(N10915), .DIN2(N10883) );
nnd2s1 U3297 ( .Q(N10941), .DIN1(N10916), .DIN2(N10885) );
nnd2s1 U3298 ( .Q(N10944), .DIN1(N10917), .DIN2(N10887) );
nnd2s1 U3299 ( .Q(N10947), .DIN1(N10918), .DIN2(N10889) );
nnd2s1 U3300 ( .Q(N10950), .DIN1(N10919), .DIN2(N10891) );
hi1s1 U3301 ( .Q(N10953), .DIN(N10892) );
nnd2s1 U3302 ( .Q(N10954), .DIN1(N10892), .DIN2(N9476) );
nnd2s1 U3303 ( .Q(N10955), .DIN1(N10922), .DIN2(N10896) );
nnd2s1 U3304 ( .Q(N10958), .DIN1(N10923), .DIN2(N10898) );
hi1s1 U3305 ( .Q(N10961), .DIN(N10899) );
nnd2s1 U3306 ( .Q(N10962), .DIN1(N10899), .DIN2(N9506) );
hi1s1 U3307 ( .Q(N10963), .DIN(N10902) );
nnd2s1 U3308 ( .Q(N10964), .DIN1(N10902), .DIN2(N9515) );
nnd2s1 U3309 ( .Q(N10969), .DIN1(N7485), .DIN2(N10934) );
nnd2s1 U3310 ( .Q(N10970), .DIN1(N7497), .DIN2(N10936) );
nnd2s1 U3311 ( .Q(N10981), .DIN1(N8718), .DIN2(N10953) );
nnd2s1 U3312 ( .Q(N10986), .DIN1(N8784), .DIN2(N10961) );
nnd2s1 U3313 ( .Q(N10987), .DIN1(N8802), .DIN2(N10963) );
hi1s1 U3314 ( .Q(N10988), .DIN(N10928) );
nnd2s1 U3315 ( .Q(N10989), .DIN1(N10928), .DIN2(N8617) );
hi1s1 U3316 ( .Q(N10990), .DIN(N10931) );
nnd2s1 U3317 ( .Q(N10991), .DIN1(N10931), .DIN2(N8626) );
nnd2s1 U3318 ( .Q(N10992), .DIN1(N10969), .DIN2(N10935) );
nnd2s1 U3319 ( .Q(N10995), .DIN1(N10970), .DIN2(N10937) );
hi1s1 U3320 ( .Q(N10998), .DIN(N10938) );
nnd2s1 U3321 ( .Q(N10999), .DIN1(N10938), .DIN2(N8646) );
hi1s1 U3322 ( .Q(N11000), .DIN(N10941) );
nnd2s1 U3323 ( .Q(N11001), .DIN1(N10941), .DIN2(N8655) );
hi1s1 U3324 ( .Q(N11002), .DIN(N10944) );
nnd2s1 U3325 ( .Q(N11003), .DIN1(N10944), .DIN2(N9456) );
hi1s1 U3326 ( .Q(N11004), .DIN(N10947) );
nnd2s1 U3327 ( .Q(N11005), .DIN1(N10947), .DIN2(N9461) );
hi1s1 U3328 ( .Q(N11006), .DIN(N10950) );
nnd2s1 U3329 ( .Q(N11007), .DIN1(N10950), .DIN2(N9465) );
nnd2s1 U3330 ( .Q(N11008), .DIN1(N10981), .DIN2(N10954) );
hi1s1 U3331 ( .Q(N11011), .DIN(N10955) );
nnd2s1 U3332 ( .Q(N11012), .DIN1(N10955), .DIN2(N9495) );
hi1s1 U3333 ( .Q(N11013), .DIN(N10958) );
nnd2s1 U3334 ( .Q(N11014), .DIN1(N10958), .DIN2(N9500) );
nnd2s1 U3335 ( .Q(N11015), .DIN1(N10986), .DIN2(N10962) );
nnd2s1 U3336 ( .Q(N11018), .DIN1(N10987), .DIN2(N10964) );
nnd2s1 U3337 ( .Q(N11023), .DIN1(N7453), .DIN2(N10988) );
nnd2s1 U3338 ( .Q(N11024), .DIN1(N7471), .DIN2(N10990) );
nnd2s1 U3339 ( .Q(N11027), .DIN1(N7509), .DIN2(N10998) );
nnd2s1 U3340 ( .Q(N11028), .DIN1(N7527), .DIN2(N11000) );
nnd2s1 U3341 ( .Q(N11029), .DIN1(N8684), .DIN2(N11002) );
nnd2s1 U3342 ( .Q(N11030), .DIN1(N8696), .DIN2(N11004) );
nnd2s1 U3343 ( .Q(N11031), .DIN1(N8702), .DIN2(N11006) );
nnd2s1 U3344 ( .Q(N11034), .DIN1(N8763), .DIN2(N11011) );
nnd2s1 U3345 ( .Q(N11035), .DIN1(N8775), .DIN2(N11013) );
hi1s1 U3346 ( .Q(N11040), .DIN(N10992) );
nnd2s1 U3347 ( .Q(N11041), .DIN1(N10992), .DIN2(N8294) );
hi1s1 U3348 ( .Q(N11042), .DIN(N10995) );
nnd2s1 U3349 ( .Q(N11043), .DIN1(N10995), .DIN2(N8295) );
nnd2s1 U3350 ( .Q(N11044), .DIN1(N11023), .DIN2(N10989) );
nnd2s1 U3351 ( .Q(N11047), .DIN1(N11024), .DIN2(N10991) );
nnd2s1 U3352 ( .Q(N11050), .DIN1(N11027), .DIN2(N10999) );
nnd2s1 U3353 ( .Q(N11053), .DIN1(N11028), .DIN2(N11001) );
nnd2s1 U3354 ( .Q(N11056), .DIN1(N11029), .DIN2(N11003) );
nnd2s1 U3355 ( .Q(N11059), .DIN1(N11030), .DIN2(N11005) );
nnd2s1 U3356 ( .Q(N11062), .DIN1(N11031), .DIN2(N11007) );
hi1s1 U3357 ( .Q(N11065), .DIN(N11008) );
nnd2s1 U3358 ( .Q(N11066), .DIN1(N11008), .DIN2(N9477) );
nnd2s1 U3359 ( .Q(N11067), .DIN1(N11034), .DIN2(N11012) );
nnd2s1 U3360 ( .Q(N11070), .DIN1(N11035), .DIN2(N11014) );
hi1s1 U3361 ( .Q(N11073), .DIN(N11015) );
nnd2s1 U3362 ( .Q(N11074), .DIN1(N11015), .DIN2(N9507) );
hi1s1 U3363 ( .Q(N11075), .DIN(N11018) );
nnd2s1 U3364 ( .Q(N11076), .DIN1(N11018), .DIN2(N9516) );
nnd2s1 U3365 ( .Q(N11077), .DIN1(N7488), .DIN2(N11040) );
nnd2s1 U3366 ( .Q(N11078), .DIN1(N7500), .DIN2(N11042) );
nnd2s1 U3367 ( .Q(N11095), .DIN1(N8721), .DIN2(N11065) );
nnd2s1 U3368 ( .Q(N11098), .DIN1(N8787), .DIN2(N11073) );
nnd2s1 U3369 ( .Q(N11099), .DIN1(N8805), .DIN2(N11075) );
nnd2s1 U3370 ( .Q(N11100), .DIN1(N11077), .DIN2(N11041) );
nnd2s1 U3371 ( .Q(N11103), .DIN1(N11078), .DIN2(N11043) );
hi1s1 U3372 ( .Q(N11106), .DIN(N11056) );
nnd2s1 U3373 ( .Q(N11107), .DIN1(N11056), .DIN2(N9319) );
hi1s1 U3374 ( .Q(N11108), .DIN(N11059) );
nnd2s1 U3375 ( .Q(N11109), .DIN1(N11059), .DIN2(N9320) );
hi1s1 U3376 ( .Q(N11110), .DIN(N11067) );
nnd2s1 U3377 ( .Q(N11111), .DIN1(N11067), .DIN2(N9381) );
hi1s1 U3378 ( .Q(N11112), .DIN(N11070) );
nnd2s1 U3379 ( .Q(N11113), .DIN1(N11070), .DIN2(N9382) );
hi1s1 U3380 ( .Q(N11114), .DIN(N11044) );
nnd2s1 U3381 ( .Q(N11115), .DIN1(N11044), .DIN2(N8618) );
hi1s1 U3382 ( .Q(N11116), .DIN(N11047) );
nnd2s1 U3383 ( .Q(N11117), .DIN1(N11047), .DIN2(N8619) );
hi1s1 U3384 ( .Q(N11118), .DIN(N11050) );
nnd2s1 U3385 ( .Q(N11119), .DIN1(N11050), .DIN2(N8647) );
hi1s1 U3386 ( .Q(N11120), .DIN(N11053) );
nnd2s1 U3387 ( .Q(N11121), .DIN1(N11053), .DIN2(N8648) );
hi1s1 U3388 ( .Q(N11122), .DIN(N11062) );
nnd2s1 U3389 ( .Q(N11123), .DIN1(N11062), .DIN2(N9466) );
nnd2s1 U3390 ( .Q(N11124), .DIN1(N11095), .DIN2(N11066) );
nnd2s1 U3391 ( .Q(N11127), .DIN1(N11098), .DIN2(N11074) );
nnd2s1 U3392 ( .Q(N11130), .DIN1(N11099), .DIN2(N11076) );
nnd2s1 U3393 ( .Q(N11137), .DIN1(N8687), .DIN2(N11106) );
nnd2s1 U3394 ( .Q(N11138), .DIN1(N8699), .DIN2(N11108) );
nnd2s1 U3395 ( .Q(N11139), .DIN1(N8766), .DIN2(N11110) );
nnd2s1 U3396 ( .Q(N11140), .DIN1(N8778), .DIN2(N11112) );
nnd2s1 U3397 ( .Q(N11141), .DIN1(N7456), .DIN2(N11114) );
nnd2s1 U3398 ( .Q(N11142), .DIN1(N7474), .DIN2(N11116) );
nnd2s1 U3399 ( .Q(N11143), .DIN1(N7512), .DIN2(N11118) );
nnd2s1 U3400 ( .Q(N11144), .DIN1(N7530), .DIN2(N11120) );
nnd2s1 U3401 ( .Q(N11145), .DIN1(N8705), .DIN2(N11122) );
and3s1 U3402 ( .Q(N11152), .DIN1(N11103), .DIN2(N8871), .DIN3(N10283) );
and3s1 U3403 ( .Q(N11153), .DIN1(N11100), .DIN2(N7655), .DIN3(N10283) );
and3s1 U3404 ( .Q(N11154), .DIN1(N11103), .DIN2(N9551), .DIN3(N10119) );
and3s1 U3405 ( .Q(N11155), .DIN1(N11100), .DIN2(N9917), .DIN3(N10119) );
nnd2s1 U3406 ( .Q(N11156), .DIN1(N11137), .DIN2(N11107) );
nnd2s1 U3407 ( .Q(N11159), .DIN1(N11138), .DIN2(N11109) );
nnd2s1 U3408 ( .Q(N11162), .DIN1(N11139), .DIN2(N11111) );
nnd2s1 U3409 ( .Q(N11165), .DIN1(N11140), .DIN2(N11113) );
nnd2s1 U3410 ( .Q(N11168), .DIN1(N11141), .DIN2(N11115) );
nnd2s1 U3411 ( .Q(N11171), .DIN1(N11142), .DIN2(N11117) );
nnd2s1 U3412 ( .Q(N11174), .DIN1(N11143), .DIN2(N11119) );
nnd2s1 U3413 ( .Q(N11177), .DIN1(N11144), .DIN2(N11121) );
nnd2s1 U3414 ( .Q(N11180), .DIN1(N11145), .DIN2(N11123) );
hi1s1 U3415 ( .Q(N11183), .DIN(N11124) );
nnd2s1 U3416 ( .Q(N11184), .DIN1(N11124), .DIN2(N9468) );
hi1s1 U3417 ( .Q(N11185), .DIN(N11127) );
nnd2s1 U3418 ( .Q(N11186), .DIN1(N11127), .DIN2(N9508) );
hi1s1 U3419 ( .Q(N11187), .DIN(N11130) );
nnd2s1 U3420 ( .Q(N11188), .DIN1(N11130), .DIN2(N9509) );
or4s1 U3421 ( .Q(N11205), .DIN1(N11152), .DIN2(N11153), .DIN3(N11154), .DIN4(N11155) );
nnd2s1 U3422 ( .Q(N11210), .DIN1(N8724), .DIN2(N11183) );
nnd2s1 U3423 ( .Q(N11211), .DIN1(N8790), .DIN2(N11185) );
nnd2s1 U3424 ( .Q(N11212), .DIN1(N8808), .DIN2(N11187) );
hi1s1 U3425 ( .Q(N11213), .DIN(N11168) );
nnd2s1 U3426 ( .Q(N11214), .DIN1(N11168), .DIN2(N8260) );
hi1s1 U3427 ( .Q(N11215), .DIN(N11171) );
nnd2s1 U3428 ( .Q(N11216), .DIN1(N11171), .DIN2(N8261) );
hi1s1 U3429 ( .Q(N11217), .DIN(N11174) );
nnd2s1 U3430 ( .Q(N11218), .DIN1(N11174), .DIN2(N8296) );
hi1s1 U3431 ( .Q(N11219), .DIN(N11177) );
nnd2s1 U3432 ( .Q(N11220), .DIN1(N11177), .DIN2(N8297) );
and3s1 U3433 ( .Q(N11222), .DIN1(N11159), .DIN2(N9575), .DIN3(N1218) );
and3s1 U3434 ( .Q(N11223), .DIN1(N11156), .DIN2(N8927), .DIN3(N1218) );
and3s1 U3435 ( .Q(N11224), .DIN1(N11159), .DIN2(N9935), .DIN3(N750) );
and3s1 U3436 ( .Q(N11225), .DIN1(N11156), .DIN2(N10132), .DIN3(N750) );
and3s1 U3437 ( .Q(N11226), .DIN1(N11165), .DIN2(N9608), .DIN3(N10497) );
and3s1 U3438 ( .Q(N11227), .DIN1(N11162), .DIN2(N9001), .DIN3(N10497) );
and3s1 U3439 ( .Q(N11228), .DIN1(N11165), .DIN2(N9949), .DIN3(N10301) );
and3s1 U3440 ( .Q(N11229), .DIN1(N11162), .DIN2(N10160), .DIN3(N10301) );
hi1s1 U3441 ( .Q(N11231), .DIN(N11180) );
nnd2s1 U3442 ( .Q(N11232), .DIN1(N11180), .DIN2(N9467) );
nnd2s1 U3443 ( .Q(N11233), .DIN1(N11210), .DIN2(N11184) );
nnd2s1 U3444 ( .Q(N11236), .DIN1(N11211), .DIN2(N11186) );
nnd2s1 U3445 ( .Q(N11239), .DIN1(N11212), .DIN2(N11188) );
nnd2s1 U3446 ( .Q(N11242), .DIN1(N7459), .DIN2(N11213) );
nnd2s1 U3447 ( .Q(N11243), .DIN1(N7462), .DIN2(N11215) );
nnd2s1 U3448 ( .Q(N11244), .DIN1(N7515), .DIN2(N11217) );
nnd2s1 U3449 ( .Q(N11245), .DIN1(N7518), .DIN2(N11219) );
hi1s1 U3450 ( .Q(N11246), .DIN(N11205) );
nnd2s1 U3451 ( .Q(N11250), .DIN1(N8708), .DIN2(N11231) );
or4s1 U3452 ( .Q(N11252), .DIN1(N11222), .DIN2(N11223), .DIN3(N11224), .DIN4(N11225) );
or4s1 U3453 ( .Q(N11257), .DIN1(N11226), .DIN2(N11227), .DIN3(N11228), .DIN4(N11229) );
nnd2s1 U3454 ( .Q(N11260), .DIN1(N11242), .DIN2(N11214) );
nnd2s1 U3455 ( .Q(N11261), .DIN1(N11243), .DIN2(N11216) );
nnd2s1 U3456 ( .Q(N11262), .DIN1(N11244), .DIN2(N11218) );
nnd2s1 U3457 ( .Q(N11263), .DIN1(N11245), .DIN2(N11220) );
hi1s1 U3458 ( .Q(N11264), .DIN(N11233) );
nnd2s1 U3459 ( .Q(N11265), .DIN1(N11233), .DIN2(N9322) );
hi1s1 U3460 ( .Q(N11267), .DIN(N11236) );
nnd2s1 U3461 ( .Q(N11268), .DIN1(N11236), .DIN2(N9383) );
hi1s1 U3462 ( .Q(N11269), .DIN(N11239) );
nnd2s1 U3463 ( .Q(N11270), .DIN1(N11239), .DIN2(N9384) );
nnd2s1 U3464 ( .Q(N11272), .DIN1(N11250), .DIN2(N11232) );
hi1s1 U3465 ( .Q(N11277), .DIN(N11261) );
and2s1 U3466 ( .Q(N11278), .DIN1(N10273), .DIN2(N11260) );
hi1s1 U3467 ( .Q(N11279), .DIN(N11263) );
and2s1 U3468 ( .Q(N11280), .DIN1(N10119), .DIN2(N11262) );
nnd2s1 U3469 ( .Q(N11282), .DIN1(N8714), .DIN2(N11264) );
hi1s1 U3470 ( .Q(N11283), .DIN(N11252) );
nnd2s1 U3471 ( .Q(N11284), .DIN1(N8793), .DIN2(N11267) );
nnd2s1 U3472 ( .Q(N11285), .DIN1(N8796), .DIN2(N11269) );
hi1s1 U3473 ( .Q(N11286), .DIN(N11257) );
and2s1 U3474 ( .Q(N11288), .DIN1(N11277), .DIN2(N10479) );
and2s1 U3475 ( .Q(N11289), .DIN1(N11279), .DIN2(N10283) );
hi1s1 U3476 ( .Q(N11290), .DIN(N11272) );
nnd2s1 U3477 ( .Q(N11291), .DIN1(N11272), .DIN2(N9321) );
nnd2s1 U3478 ( .Q(N11292), .DIN1(N11282), .DIN2(N11265) );
nnd2s1 U3479 ( .Q(N11293), .DIN1(N11284), .DIN2(N11268) );
nnd2s1 U3480 ( .Q(N11294), .DIN1(N11285), .DIN2(N11270) );
nnd2s1 U3481 ( .Q(N11295), .DIN1(N8711), .DIN2(N11290) );
hi1s1 U3482 ( .Q(N11296), .DIN(N11292) );
hi1s1 U3483 ( .Q(N11297), .DIN(N11294) );
and2s1 U3484 ( .Q(N11298), .DIN1(N10301), .DIN2(N11293) );
or2s1 U3485 ( .Q(N11299), .DIN1(N11288), .DIN2(N11278) );
or2s1 U3486 ( .Q(N11302), .DIN1(N11289), .DIN2(N11280) );
nnd2s1 U3487 ( .Q(N11307), .DIN1(N11295), .DIN2(N11291) );
and2s1 U3488 ( .Q(N11308), .DIN1(N11296), .DIN2(N1218) );
and2s1 U3489 ( .Q(N11309), .DIN1(N11297), .DIN2(N10497) );
nnd2s1 U3490 ( .Q(N11312), .DIN1(N11302), .DIN2(N11246) );
nnd2s1 U3491 ( .Q(N11313), .DIN1(N11299), .DIN2(N10836) );
hi1s1 U3492 ( .Q(N11314), .DIN(N11299) );
hi1s1 U3493 ( .Q(N11315), .DIN(N11302) );
and2s1 U3494 ( .Q(N11316), .DIN1(N750), .DIN2(N11307) );
or2s1 U3495 ( .Q(N11317), .DIN1(N11309), .DIN2(N11298) );
nnd2s1 U3496 ( .Q(N11320), .DIN1(N11205), .DIN2(N11315) );
nnd2s1 U3497 ( .Q(N11321), .DIN1(N10739), .DIN2(N11314) );
or2s1 U3498 ( .Q(N11323), .DIN1(N11308), .DIN2(N11316) );
nnd2s1 U3499 ( .Q(N11327), .DIN1(N11312), .DIN2(N11320) );
nnd2s1 U3500 ( .Q(N11328), .DIN1(N11313), .DIN2(N11321) );
nnd2s1 U3501 ( .Q(N11329), .DIN1(N11317), .DIN2(N11286) );
hi1s1 U3502 ( .Q(N11331), .DIN(N11317) );
hi1s1 U3503 ( .Q(N11333), .DIN(N11327) );
hi1s1 U3504 ( .Q(N11334), .DIN(N11328) );
nnd2s1 U3505 ( .Q(N11335), .DIN1(N11257), .DIN2(N11331) );
nnd2s1 U3506 ( .Q(N11336), .DIN1(N11323), .DIN2(N11283) );
hi1s1 U3507 ( .Q(N11337), .DIN(N11323) );
nnd2s1 U3508 ( .Q(N11338), .DIN1(N11329), .DIN2(N11335) );
nnd2s1 U3509 ( .Q(N11339), .DIN1(N11252), .DIN2(N11337) );
hi1s1 U3510 ( .Q(N11340), .DIN(N11338) );
nnd2s1 U3511 ( .Q(N11341), .DIN1(N11336), .DIN2(N11339) );
hi1s1 U3512 ( .Q(N11342), .DIN(N11341) );
nb1s1 U3513 ( .Q(B241), .DIN(N241) );
endmodule
