module mips_16_core_top_syn_copy_renamed ( clk, rst, pc_7_, pc_6_, pc_5_, pc_4_, pc_3_, pc_2_, pc_1_, pc_0_ , MEM_stage_inst_N6, EX_stage_inst_N4, MEM_stage_inst_N4, EX_stage_inst_N5, MEM_stage_inst_N5, EX_stage_inst_N6, EX_stage_inst_N3, EX_stage_inst_N7, EX_stage_inst_N24, MEM_stage_inst_N7, EX_stage_inst_N40, MEM_stage_inst_N39, EX_stage_inst_N23, EX_stage_inst_N25, MEM_stage_inst_N24, EX_stage_inst_N8, EX_stage_inst_N33, MEM_stage_inst_N32, EX_stage_inst_N16, EX_stage_inst_N35, MEM_stage_inst_N34, EX_stage_inst_N18, EX_stage_inst_N37, MEM_stage_inst_N36, EX_stage_inst_N20, EX_stage_inst_N39, MEM_stage_inst_N38, EX_stage_inst_N22, EX_stage_inst_N29, MEM_stage_inst_N28, EX_stage_inst_N12, EX_stage_inst_N31, MEM_stage_inst_N30, EX_stage_inst_N14, EX_stage_inst_N36, MEM_stage_inst_N35, EX_stage_inst_N19, EX_stage_inst_N38, MEM_stage_inst_N37, EX_stage_inst_N21, EX_stage_inst_N27, MEM_stage_inst_N26, EX_stage_inst_N10, EX_stage_inst_N28, MEM_stage_inst_N27, EX_stage_inst_N11, EX_stage_inst_N26, MEM_stage_inst_N25, EX_stage_inst_N9, EX_stage_inst_N30, MEM_stage_inst_N29, EX_stage_inst_N13, EX_stage_inst_N34, MEM_stage_inst_N33, EX_stage_inst_N17, EX_stage_inst_N32, MEM_stage_inst_N31, EX_stage_inst_N15, MEM_stage_inst_N8, MEM_stage_inst_N9, MEM_stage_inst_N10, MEM_stage_inst_N11, MEM_stage_inst_N12, MEM_stage_inst_N13, MEM_stage_inst_N14, MEM_stage_inst_N15, MEM_stage_inst_N16, MEM_stage_inst_N17, MEM_stage_inst_N18, MEM_stage_inst_N19, MEM_stage_inst_N20, MEM_stage_inst_N21, MEM_stage_inst_N22, MEM_stage_inst_N23, n1734, n3520, n1731, n3517, n1730, n1741, n1729, n1739, n1728, n1727, n1724, n3521, n1722, n3518, n1725, n1723, n1713, n1714, n1726, n1721, n1720, n1719, n1718, ID_stage_inst_ir_dest_with_bubble_0, n1717, ID_stage_inst_ir_dest_with_bubble_1, n1716, ID_stage_inst_ir_dest_with_bubble_2, n1715, n1712, ID_stage_inst_ex_alu_cmd_1, ID_stage_inst_ex_alu_cmd_0, ID_stage_inst_ex_alu_cmd_2, ID_stage_inst_write_back_result_mux, ID_stage_inst_write_back_en, n1738, n1735, reg_read_data_1_15, n1606, n1605, n3519, n1604, n1603, n1602, n1601, reg_read_data_2_15, ID_stage_inst_ex_alu_src2_15, n1711, n1710, n1709, n1708, n1707, n1706, n1705, reg_read_data_2_0, reg_read_data_1_0, n1655, n1654, n1653, n1652, n1651, n1650, n1649, reg_read_data_2_8, ID_stage_inst_ex_alu_src2_8, reg_read_data_1_8, n1641, n1640, n1639, n1638, n1637, n1636, n1635, reg_read_data_2_10, ID_stage_inst_ex_alu_src2_10, reg_read_data_1_10, n1627, n1626, n1625, n1624, n1623, n1622, n1621, reg_read_data_2_12, ID_stage_inst_ex_alu_src2_12, reg_read_data_1_12, n1613, n1612, n1611, n1610, n1609, n1608, n1607, reg_read_data_2_14, ID_stage_inst_ex_alu_src2_14, reg_read_data_1_14, n1683, n1682, n1681, n1680, n1679, n1678, n1677, reg_read_data_2_4, ID_stage_inst_ex_alu_src2_4, reg_read_data_1_4, n1669, n1668, n1667, n1666, n1665, n1664, n1663, reg_read_data_2_6, ID_stage_inst_ex_alu_src2_6, reg_read_data_1_6, n1634, n1633, n1632, n1631, n1630, n1629, n1628, reg_read_data_2_11, ID_stage_inst_ex_alu_src2_11, reg_read_data_1_11, n1620, n1619, n1618, n1617, n1616, n1615, n1614, reg_read_data_2_13, ID_stage_inst_ex_alu_src2_13, reg_read_data_1_13, n1697, n1696, n1695, n1694, n1693, n1692, n1691, reg_read_data_2_2, reg_read_data_1_2, n1690, n1689, n1688, n1687, n1686, n1685, n1684, reg_read_data_2_3, reg_read_data_1_3, n1704, n1703, n1702, n1701, n1700, n1699, n1698, reg_read_data_2_1, reg_read_data_1_1, n1676, n1675, n1674, n1673, n1672, n1671, n1670, reg_read_data_2_5, ID_stage_inst_ex_alu_src2_5, reg_read_data_1_5, n1648, n1647, n1646, n1645, n1644, n1643, n1642, reg_read_data_2_9, ID_stage_inst_ex_alu_src2_9, reg_read_data_1_9, n1662, n1661, n1660, n1659, n1658, n1657, n1656, reg_read_data_2_7, ID_stage_inst_ex_alu_src2_7, reg_read_data_1_7, n1732, ID_stage_inst_ex_alu_src2_1, MEM_stage_inst_N3, ID_stage_inst_ex_alu_src2_2, ID_stage_inst_ex_alu_src2_0, ID_stage_inst_ex_alu_src2_3, n1733, MEM_stage_inst_dmem_n8763, MEM_stage_inst_dmem_n21529, MEM_stage_inst_dmem_n8764, MEM_stage_inst_dmem_n21573, MEM_stage_inst_dmem_n8765, MEM_stage_inst_dmem_n21564, MEM_stage_inst_dmem_n8766, MEM_stage_inst_dmem_n21580, MEM_stage_inst_dmem_n8767, MEM_stage_inst_dmem_n21538, MEM_stage_inst_dmem_n8768, MEM_stage_inst_dmem_n21540, MEM_stage_inst_dmem_n8769, MEM_stage_inst_dmem_n21605, MEM_stage_inst_dmem_n8770, MEM_stage_inst_dmem_n21579, MEM_stage_inst_dmem_n8771, MEM_stage_inst_dmem_n21575, MEM_stage_inst_dmem_n8772, MEM_stage_inst_dmem_n21584, MEM_stage_inst_dmem_n8773, MEM_stage_inst_dmem_n21597, MEM_stage_inst_dmem_n8774, MEM_stage_inst_dmem_n21542, MEM_stage_inst_dmem_n8775, MEM_stage_inst_dmem_n21586, MEM_stage_inst_dmem_n8776, MEM_stage_inst_dmem_n21570, MEM_stage_inst_dmem_n8777, MEM_stage_inst_dmem_n21546, MEM_stage_inst_dmem_n8778, MEM_stage_inst_dmem_n21532, MEM_stage_inst_dmem_n8779, MEM_stage_inst_dmem_n21549, MEM_stage_inst_dmem_n8780, MEM_stage_inst_dmem_n21553, MEM_stage_inst_dmem_n8781, MEM_stage_inst_dmem_n21629, MEM_stage_inst_dmem_n8782, MEM_stage_inst_dmem_n21547, MEM_stage_inst_dmem_n8783, MEM_stage_inst_dmem_n21572, MEM_stage_inst_dmem_n8784, MEM_stage_inst_dmem_n21559, MEM_stage_inst_dmem_n8785, MEM_stage_inst_dmem_n21600, MEM_stage_inst_dmem_n8786, MEM_stage_inst_dmem_n21554, MEM_stage_inst_dmem_n8787, MEM_stage_inst_dmem_n8788, MEM_stage_inst_dmem_n8789, MEM_stage_inst_dmem_n8790, MEM_stage_inst_dmem_n21591, MEM_stage_inst_dmem_n8791, MEM_stage_inst_dmem_n21527, MEM_stage_inst_dmem_n8792, MEM_stage_inst_dmem_n21622, MEM_stage_inst_dmem_n8793, MEM_stage_inst_dmem_n8794, MEM_stage_inst_dmem_n21590, MEM_stage_inst_dmem_n8795, MEM_stage_inst_dmem_n21610, MEM_stage_inst_dmem_n8796, MEM_stage_inst_dmem_n21612, MEM_stage_inst_dmem_n8797, MEM_stage_inst_dmem_n21616, MEM_stage_inst_dmem_n8798, MEM_stage_inst_dmem_n21582, MEM_stage_inst_dmem_n8799, MEM_stage_inst_dmem_n21537, MEM_stage_inst_dmem_n8800, MEM_stage_inst_dmem_n21602, MEM_stage_inst_dmem_n8801, MEM_stage_inst_dmem_n21574, MEM_stage_inst_dmem_n8802, MEM_stage_inst_dmem_n21566, MEM_stage_inst_dmem_n8803, MEM_stage_inst_dmem_n8804, MEM_stage_inst_dmem_n21543, MEM_stage_inst_dmem_n8805, MEM_stage_inst_dmem_n8806, MEM_stage_inst_dmem_n8807, MEM_stage_inst_dmem_n8808, MEM_stage_inst_dmem_n8809, MEM_stage_inst_dmem_n8810, MEM_stage_inst_dmem_n8811, MEM_stage_inst_dmem_n21619, MEM_stage_inst_dmem_n8812, MEM_stage_inst_dmem_n21525, MEM_stage_inst_dmem_n8813, MEM_stage_inst_dmem_n21593, MEM_stage_inst_dmem_n8814, MEM_stage_inst_dmem_n8815, MEM_stage_inst_dmem_n21524, MEM_stage_inst_dmem_n8816, MEM_stage_inst_dmem_n21511, MEM_stage_inst_dmem_n8817, MEM_stage_inst_dmem_n21556, MEM_stage_inst_dmem_n8818, MEM_stage_inst_dmem_n8819, MEM_stage_inst_dmem_n21576, MEM_stage_inst_dmem_n8820, MEM_stage_inst_dmem_n8821, MEM_stage_inst_dmem_n8822, MEM_stage_inst_dmem_n21544, MEM_stage_inst_dmem_n8823, MEM_stage_inst_dmem_n8824, MEM_stage_inst_dmem_n21519, MEM_stage_inst_dmem_n8825, MEM_stage_inst_dmem_n21510, MEM_stage_inst_dmem_n8826, MEM_stage_inst_dmem_n8827, MEM_stage_inst_dmem_n21569, MEM_stage_inst_dmem_n8828, MEM_stage_inst_dmem_n21625, MEM_stage_inst_dmem_n8829, MEM_stage_inst_dmem_n21608, MEM_stage_inst_dmem_n8830, MEM_stage_inst_dmem_n21563, MEM_stage_inst_dmem_n8831, MEM_stage_inst_dmem_n21526, MEM_stage_inst_dmem_n8832, MEM_stage_inst_dmem_n21588, MEM_stage_inst_dmem_n8833, MEM_stage_inst_dmem_n21618, MEM_stage_inst_dmem_n8834, MEM_stage_inst_dmem_n21624, MEM_stage_inst_dmem_n8835, MEM_stage_inst_dmem_n21522, MEM_stage_inst_dmem_n8836, MEM_stage_inst_dmem_n21615, MEM_stage_inst_dmem_n8837, MEM_stage_inst_dmem_n21617, MEM_stage_inst_dmem_n8838, MEM_stage_inst_dmem_n8839, MEM_stage_inst_dmem_n21555, MEM_stage_inst_dmem_n8840, MEM_stage_inst_dmem_n21606, MEM_stage_inst_dmem_n8841, MEM_stage_inst_dmem_n21539, MEM_stage_inst_dmem_n8842, MEM_stage_inst_dmem_n21568, MEM_stage_inst_dmem_n8843, MEM_stage_inst_dmem_n8844, MEM_stage_inst_dmem_n8845, MEM_stage_inst_dmem_n8846, MEM_stage_inst_dmem_n21594, MEM_stage_inst_dmem_n8847, MEM_stage_inst_dmem_n21548, MEM_stage_inst_dmem_n8848, MEM_stage_inst_dmem_n21565, MEM_stage_inst_dmem_n8849, MEM_stage_inst_dmem_n8850, MEM_stage_inst_dmem_n8851, MEM_stage_inst_dmem_n21534, MEM_stage_inst_dmem_n8852, MEM_stage_inst_dmem_n8853, MEM_stage_inst_dmem_n21609, MEM_stage_inst_dmem_n8854, MEM_stage_inst_dmem_n8855, MEM_stage_inst_dmem_n21621, MEM_stage_inst_dmem_n8856, MEM_stage_inst_dmem_n8857, MEM_stage_inst_dmem_n21633, MEM_stage_inst_dmem_n8858, MEM_stage_inst_dmem_n21604, MEM_stage_inst_dmem_n8859, MEM_stage_inst_dmem_n21518, MEM_stage_inst_dmem_n8860, MEM_stage_inst_dmem_n8861, MEM_stage_inst_dmem_n8862, MEM_stage_inst_dmem_n8863, MEM_stage_inst_dmem_n21636, MEM_stage_inst_dmem_n8864, MEM_stage_inst_dmem_n8865, MEM_stage_inst_dmem_n8866, MEM_stage_inst_dmem_n8867, MEM_stage_inst_dmem_n21589, MEM_stage_inst_dmem_n8868, MEM_stage_inst_dmem_n8869, MEM_stage_inst_dmem_n8870, MEM_stage_inst_dmem_n8871, MEM_stage_inst_dmem_n8872, MEM_stage_inst_dmem_n8873, MEM_stage_inst_dmem_n8874, MEM_stage_inst_dmem_n21514, MEM_stage_inst_dmem_n8875, MEM_stage_inst_dmem_n21592, MEM_stage_inst_dmem_n8876, MEM_stage_inst_dmem_n21628, MEM_stage_inst_dmem_n8877, MEM_stage_inst_dmem_n21513, MEM_stage_inst_dmem_n8878, MEM_stage_inst_dmem_n8879, MEM_stage_inst_dmem_n21623, MEM_stage_inst_dmem_n8880, MEM_stage_inst_dmem_n21583, MEM_stage_inst_dmem_n8881, MEM_stage_inst_dmem_n21613, MEM_stage_inst_dmem_n8882, MEM_stage_inst_dmem_n8883, MEM_stage_inst_dmem_n21516, MEM_stage_inst_dmem_n8884, MEM_stage_inst_dmem_n8885, MEM_stage_inst_dmem_n21509, MEM_stage_inst_dmem_n8886, MEM_stage_inst_dmem_n8887, MEM_stage_inst_dmem_n21558, MEM_stage_inst_dmem_n8888, MEM_stage_inst_dmem_n8889, MEM_stage_inst_dmem_n8890, MEM_stage_inst_dmem_n8891, MEM_stage_inst_dmem_n8892, MEM_stage_inst_dmem_n8893, MEM_stage_inst_dmem_n8894, MEM_stage_inst_dmem_n8895, MEM_stage_inst_dmem_n8896, MEM_stage_inst_dmem_n21587, MEM_stage_inst_dmem_n8897, MEM_stage_inst_dmem_n8898, MEM_stage_inst_dmem_n21626, MEM_stage_inst_dmem_n8899, MEM_stage_inst_dmem_n21599, MEM_stage_inst_dmem_n8900, MEM_stage_inst_dmem_n8901, MEM_stage_inst_dmem_n21598, MEM_stage_inst_dmem_n8902, MEM_stage_inst_dmem_n21552, MEM_stage_inst_dmem_n8903, MEM_stage_inst_dmem_n8904, MEM_stage_inst_dmem_n8905, MEM_stage_inst_dmem_n21523, MEM_stage_inst_dmem_n8906, MEM_stage_inst_dmem_n21517, MEM_stage_inst_dmem_n8907, MEM_stage_inst_dmem_n21601, MEM_stage_inst_dmem_n8908, MEM_stage_inst_dmem_n21603, MEM_stage_inst_dmem_n8909, MEM_stage_inst_dmem_n8910, MEM_stage_inst_dmem_n8911, MEM_stage_inst_dmem_n8912, MEM_stage_inst_dmem_n21515, MEM_stage_inst_dmem_n8913, MEM_stage_inst_dmem_n8914, MEM_stage_inst_dmem_n21578, MEM_stage_inst_dmem_n8915, MEM_stage_inst_dmem_n8916, MEM_stage_inst_dmem_n8917, MEM_stage_inst_dmem_n8918, MEM_stage_inst_dmem_n8919, MEM_stage_inst_dmem_n8920, MEM_stage_inst_dmem_n8921, MEM_stage_inst_dmem_n8922, MEM_stage_inst_dmem_n21551, MEM_stage_inst_dmem_n8923, MEM_stage_inst_dmem_n8924, MEM_stage_inst_dmem_n21620, MEM_stage_inst_dmem_n8925, MEM_stage_inst_dmem_n8926, MEM_stage_inst_dmem_n8927, MEM_stage_inst_dmem_n8928, MEM_stage_inst_dmem_n8929, MEM_stage_inst_dmem_n8930, MEM_stage_inst_dmem_n8931, MEM_stage_inst_dmem_n8932, MEM_stage_inst_dmem_n21596, MEM_stage_inst_dmem_n8933, MEM_stage_inst_dmem_n8934, MEM_stage_inst_dmem_n8935, MEM_stage_inst_dmem_n8936, MEM_stage_inst_dmem_n8937, MEM_stage_inst_dmem_n21550, MEM_stage_inst_dmem_n8938, MEM_stage_inst_dmem_n8939, MEM_stage_inst_dmem_n8940, MEM_stage_inst_dmem_n21632, MEM_stage_inst_dmem_n8941, MEM_stage_inst_dmem_n21635, MEM_stage_inst_dmem_n8942, MEM_stage_inst_dmem_n8943, MEM_stage_inst_dmem_n8944, MEM_stage_inst_dmem_n8945, MEM_stage_inst_dmem_n8946, MEM_stage_inst_dmem_n8947, MEM_stage_inst_dmem_n8948, MEM_stage_inst_dmem_n8949, MEM_stage_inst_dmem_n8950, MEM_stage_inst_dmem_n8951, MEM_stage_inst_dmem_n21611, MEM_stage_inst_dmem_n8952, MEM_stage_inst_dmem_n8953, MEM_stage_inst_dmem_n8954, MEM_stage_inst_dmem_n21512, MEM_stage_inst_dmem_n8955, MEM_stage_inst_dmem_n8956, MEM_stage_inst_dmem_n21607, MEM_stage_inst_dmem_n8957, MEM_stage_inst_dmem_n21545, MEM_stage_inst_dmem_n8958, MEM_stage_inst_dmem_n8959, MEM_stage_inst_dmem_n8960, MEM_stage_inst_dmem_n8961, MEM_stage_inst_dmem_n8962, MEM_stage_inst_dmem_n8963, MEM_stage_inst_dmem_n8964, MEM_stage_inst_dmem_n8965, MEM_stage_inst_dmem_n21581, MEM_stage_inst_dmem_n8966, MEM_stage_inst_dmem_n8967, MEM_stage_inst_dmem_n8968, MEM_stage_inst_dmem_n8969, MEM_stage_inst_dmem_n8970, MEM_stage_inst_dmem_n8971, MEM_stage_inst_dmem_n8972, MEM_stage_inst_dmem_n8973, MEM_stage_inst_dmem_n21520, MEM_stage_inst_dmem_n8974, MEM_stage_inst_dmem_n8975, MEM_stage_inst_dmem_n21560, MEM_stage_inst_dmem_n8976, MEM_stage_inst_dmem_n8977, MEM_stage_inst_dmem_n8978, MEM_stage_inst_dmem_n8979, MEM_stage_inst_dmem_n8980, MEM_stage_inst_dmem_n8981, MEM_stage_inst_dmem_n8982, MEM_stage_inst_dmem_n8983, MEM_stage_inst_dmem_n8984, MEM_stage_inst_dmem_n8985, MEM_stage_inst_dmem_n8986, MEM_stage_inst_dmem_n8987, MEM_stage_inst_dmem_n8988, MEM_stage_inst_dmem_n21585, MEM_stage_inst_dmem_n8989, MEM_stage_inst_dmem_n8990, MEM_stage_inst_dmem_n8991, MEM_stage_inst_dmem_n8992, MEM_stage_inst_dmem_n8993, MEM_stage_inst_dmem_n8994, MEM_stage_inst_dmem_n8995, MEM_stage_inst_dmem_n8996, MEM_stage_inst_dmem_n8997, MEM_stage_inst_dmem_n21530, MEM_stage_inst_dmem_n8998, MEM_stage_inst_dmem_n8999, MEM_stage_inst_dmem_n21535, MEM_stage_inst_dmem_n9000, MEM_stage_inst_dmem_n9001, MEM_stage_inst_dmem_n9002, MEM_stage_inst_dmem_n9003, MEM_stage_inst_dmem_n9004, MEM_stage_inst_dmem_n9005, MEM_stage_inst_dmem_n9006, MEM_stage_inst_dmem_n9007, MEM_stage_inst_dmem_n9008, MEM_stage_inst_dmem_n9009, MEM_stage_inst_dmem_n9010, MEM_stage_inst_dmem_n9011, MEM_stage_inst_dmem_n21614, MEM_stage_inst_dmem_n9012, MEM_stage_inst_dmem_n9013, MEM_stage_inst_dmem_n9014, MEM_stage_inst_dmem_n9015, MEM_stage_inst_dmem_n9016, MEM_stage_inst_dmem_n9017, MEM_stage_inst_dmem_n21577, MEM_stage_inst_dmem_n9018, MEM_stage_inst_dmem_n9019, MEM_stage_inst_dmem_n9020, MEM_stage_inst_dmem_n9021, MEM_stage_inst_dmem_n9022, MEM_stage_inst_dmem_n9023, MEM_stage_inst_dmem_n9024, MEM_stage_inst_dmem_n9025, MEM_stage_inst_dmem_n9026, MEM_stage_inst_dmem_n9027, MEM_stage_inst_dmem_n9028, MEM_stage_inst_dmem_n9029, MEM_stage_inst_dmem_n9030, MEM_stage_inst_dmem_n9031, MEM_stage_inst_dmem_n21595, MEM_stage_inst_dmem_n9032, MEM_stage_inst_dmem_n9033, MEM_stage_inst_dmem_n9034, MEM_stage_inst_dmem_n9035, MEM_stage_inst_dmem_n21531, MEM_stage_inst_dmem_n9036, MEM_stage_inst_dmem_n9037, MEM_stage_inst_dmem_n9038, MEM_stage_inst_dmem_n9039, MEM_stage_inst_dmem_n9040, MEM_stage_inst_dmem_n9041, MEM_stage_inst_dmem_n9042, MEM_stage_inst_dmem_n9043, MEM_stage_inst_dmem_n9044, MEM_stage_inst_dmem_n9045, MEM_stage_inst_dmem_n9046, MEM_stage_inst_dmem_n9047, MEM_stage_inst_dmem_n9048, MEM_stage_inst_dmem_n9049, MEM_stage_inst_dmem_n9050, MEM_stage_inst_dmem_n9051, MEM_stage_inst_dmem_n21528, MEM_stage_inst_dmem_n9052, MEM_stage_inst_dmem_n9053, MEM_stage_inst_dmem_n9054, MEM_stage_inst_dmem_n9055, MEM_stage_inst_dmem_n9056, MEM_stage_inst_dmem_n9057, MEM_stage_inst_dmem_n9058, MEM_stage_inst_dmem_n9059, MEM_stage_inst_dmem_n9060, MEM_stage_inst_dmem_n9061, MEM_stage_inst_dmem_n9062, MEM_stage_inst_dmem_n9063, MEM_stage_inst_dmem_n9064, MEM_stage_inst_dmem_n21631, MEM_stage_inst_dmem_n9065, MEM_stage_inst_dmem_n9066, MEM_stage_inst_dmem_n21634, MEM_stage_inst_dmem_n9067, MEM_stage_inst_dmem_n9068, MEM_stage_inst_dmem_n9069, MEM_stage_inst_dmem_n9070, MEM_stage_inst_dmem_n21627, MEM_stage_inst_dmem_n9071, MEM_stage_inst_dmem_n9072, MEM_stage_inst_dmem_n9073, MEM_stage_inst_dmem_n9074, MEM_stage_inst_dmem_n9075, MEM_stage_inst_dmem_n9076, MEM_stage_inst_dmem_n9077, MEM_stage_inst_dmem_n9078, MEM_stage_inst_dmem_n9079, MEM_stage_inst_dmem_n21562, MEM_stage_inst_dmem_n9080, MEM_stage_inst_dmem_n9081, MEM_stage_inst_dmem_n21557, MEM_stage_inst_dmem_n9082, MEM_stage_inst_dmem_n9083, MEM_stage_inst_dmem_n9084, MEM_stage_inst_dmem_n9085, MEM_stage_inst_dmem_n9086, MEM_stage_inst_dmem_n9087, MEM_stage_inst_dmem_n9088, MEM_stage_inst_dmem_n9089, MEM_stage_inst_dmem_n9090, MEM_stage_inst_dmem_n9091, MEM_stage_inst_dmem_n9092, MEM_stage_inst_dmem_n9093, MEM_stage_inst_dmem_n9094, MEM_stage_inst_dmem_n9095, MEM_stage_inst_dmem_n21571, MEM_stage_inst_dmem_n9096, MEM_stage_inst_dmem_n9097, MEM_stage_inst_dmem_n9098, MEM_stage_inst_dmem_n9099, MEM_stage_inst_dmem_n9100, MEM_stage_inst_dmem_n9101, MEM_stage_inst_dmem_n9102, MEM_stage_inst_dmem_n9103, MEM_stage_inst_dmem_n9104, MEM_stage_inst_dmem_n9105, MEM_stage_inst_dmem_n9106, MEM_stage_inst_dmem_n9107, MEM_stage_inst_dmem_n9108, MEM_stage_inst_dmem_n9109, MEM_stage_inst_dmem_n9110, MEM_stage_inst_dmem_n9111, MEM_stage_inst_dmem_n9112, MEM_stage_inst_dmem_n9113, MEM_stage_inst_dmem_n21561, MEM_stage_inst_dmem_n9114, MEM_stage_inst_dmem_n9115, MEM_stage_inst_dmem_n9116, MEM_stage_inst_dmem_n9117, MEM_stage_inst_dmem_n9118, MEM_stage_inst_dmem_n9119, MEM_stage_inst_dmem_n9120, MEM_stage_inst_dmem_n9121, MEM_stage_inst_dmem_n9122, MEM_stage_inst_dmem_n9123, MEM_stage_inst_dmem_n9124, MEM_stage_inst_dmem_n9125, MEM_stage_inst_dmem_n9126, MEM_stage_inst_dmem_n9127, MEM_stage_inst_dmem_n9128, MEM_stage_inst_dmem_n9129, MEM_stage_inst_dmem_n9130, MEM_stage_inst_dmem_n9131, MEM_stage_inst_dmem_n21541, MEM_stage_inst_dmem_n9132, MEM_stage_inst_dmem_n9133, MEM_stage_inst_dmem_n9134, MEM_stage_inst_dmem_n9135, MEM_stage_inst_dmem_n21567, MEM_stage_inst_dmem_n9136, MEM_stage_inst_dmem_n9137, MEM_stage_inst_dmem_n9138, MEM_stage_inst_dmem_n9139, MEM_stage_inst_dmem_n9140, MEM_stage_inst_dmem_n9141, MEM_stage_inst_dmem_n9142, MEM_stage_inst_dmem_n9143, MEM_stage_inst_dmem_n9144, MEM_stage_inst_dmem_n9145, MEM_stage_inst_dmem_n9146, MEM_stage_inst_dmem_n9147, MEM_stage_inst_dmem_n9148, MEM_stage_inst_dmem_n9149, MEM_stage_inst_dmem_n9150, MEM_stage_inst_dmem_n9151, MEM_stage_inst_dmem_n9152, MEM_stage_inst_dmem_n9153, MEM_stage_inst_dmem_n9154, MEM_stage_inst_dmem_n9155, MEM_stage_inst_dmem_n9156, MEM_stage_inst_dmem_n9157, MEM_stage_inst_dmem_n9158, MEM_stage_inst_dmem_n9159, MEM_stage_inst_dmem_n9160, MEM_stage_inst_dmem_n9161, MEM_stage_inst_dmem_n9162, MEM_stage_inst_dmem_n9163, MEM_stage_inst_dmem_n9164, MEM_stage_inst_dmem_n9165, MEM_stage_inst_dmem_n9166, MEM_stage_inst_dmem_n9167, MEM_stage_inst_dmem_n9168, MEM_stage_inst_dmem_n9169, MEM_stage_inst_dmem_n9170, MEM_stage_inst_dmem_n9171, MEM_stage_inst_dmem_n9172, MEM_stage_inst_dmem_n9173, MEM_stage_inst_dmem_n9174, MEM_stage_inst_dmem_n9175, MEM_stage_inst_dmem_n9176, MEM_stage_inst_dmem_n9177, MEM_stage_inst_dmem_n9178, MEM_stage_inst_dmem_n9179, MEM_stage_inst_dmem_n9180, MEM_stage_inst_dmem_n9181, MEM_stage_inst_dmem_n9182, MEM_stage_inst_dmem_n9183, MEM_stage_inst_dmem_n9184, MEM_stage_inst_dmem_n9185, MEM_stage_inst_dmem_n9186, MEM_stage_inst_dmem_n9187, MEM_stage_inst_dmem_n9188, MEM_stage_inst_dmem_n9189, MEM_stage_inst_dmem_n9190, MEM_stage_inst_dmem_n9191, MEM_stage_inst_dmem_n9192, MEM_stage_inst_dmem_n9193, MEM_stage_inst_dmem_n9194, MEM_stage_inst_dmem_n9195, MEM_stage_inst_dmem_n21630, MEM_stage_inst_dmem_n9196, MEM_stage_inst_dmem_n9197, MEM_stage_inst_dmem_n9198, MEM_stage_inst_dmem_n9199, MEM_stage_inst_dmem_n9200, MEM_stage_inst_dmem_n9201, MEM_stage_inst_dmem_n9202, MEM_stage_inst_dmem_n9203, MEM_stage_inst_dmem_n9204, MEM_stage_inst_dmem_n9205, MEM_stage_inst_dmem_n9206, MEM_stage_inst_dmem_n9207, MEM_stage_inst_dmem_n9208, MEM_stage_inst_dmem_n9209, MEM_stage_inst_dmem_n9210, MEM_stage_inst_dmem_n9211, MEM_stage_inst_dmem_n9212, MEM_stage_inst_dmem_n9213, MEM_stage_inst_dmem_n9214, MEM_stage_inst_dmem_n9215, MEM_stage_inst_dmem_n9216, MEM_stage_inst_dmem_n9217, MEM_stage_inst_dmem_n9218, MEM_stage_inst_dmem_n9219, MEM_stage_inst_dmem_n9220, MEM_stage_inst_dmem_n9221, MEM_stage_inst_dmem_n9222, MEM_stage_inst_dmem_n9223, MEM_stage_inst_dmem_n9224, MEM_stage_inst_dmem_n9225, MEM_stage_inst_dmem_n9226, MEM_stage_inst_dmem_n9227, MEM_stage_inst_dmem_n9228, MEM_stage_inst_dmem_n9229, MEM_stage_inst_dmem_n9230, MEM_stage_inst_dmem_n9231, MEM_stage_inst_dmem_n9232, MEM_stage_inst_dmem_n9233, MEM_stage_inst_dmem_n9234, MEM_stage_inst_dmem_n9235, MEM_stage_inst_dmem_n9236, MEM_stage_inst_dmem_n9237, MEM_stage_inst_dmem_n9238, MEM_stage_inst_dmem_n9239, MEM_stage_inst_dmem_n9240, MEM_stage_inst_dmem_n9241, MEM_stage_inst_dmem_n21521, MEM_stage_inst_dmem_n9242, MEM_stage_inst_dmem_n9243, MEM_stage_inst_dmem_n9244, MEM_stage_inst_dmem_n9245, MEM_stage_inst_dmem_n9246, MEM_stage_inst_dmem_n9247, MEM_stage_inst_dmem_n9248, MEM_stage_inst_dmem_n9249, MEM_stage_inst_dmem_n9250, MEM_stage_inst_dmem_n9251, MEM_stage_inst_dmem_n9252, MEM_stage_inst_dmem_n9253, MEM_stage_inst_dmem_n9254, MEM_stage_inst_dmem_n9255, MEM_stage_inst_dmem_n9256, MEM_stage_inst_dmem_n9257, MEM_stage_inst_dmem_n9258, MEM_stage_inst_dmem_n9259, MEM_stage_inst_dmem_n9260, MEM_stage_inst_dmem_n9261, MEM_stage_inst_dmem_n9262, MEM_stage_inst_dmem_n9263, MEM_stage_inst_dmem_n9264, MEM_stage_inst_dmem_n9265, MEM_stage_inst_dmem_n9266, MEM_stage_inst_dmem_n9267, MEM_stage_inst_dmem_n9268, MEM_stage_inst_dmem_n9269, MEM_stage_inst_dmem_n9270, MEM_stage_inst_dmem_n9271, MEM_stage_inst_dmem_n9272, MEM_stage_inst_dmem_n9273, MEM_stage_inst_dmem_n9274, MEM_stage_inst_dmem_n9275, MEM_stage_inst_dmem_n9276, MEM_stage_inst_dmem_n9277, MEM_stage_inst_dmem_n9278, MEM_stage_inst_dmem_n9279, MEM_stage_inst_dmem_n9280, MEM_stage_inst_dmem_n9281, MEM_stage_inst_dmem_n9282, MEM_stage_inst_dmem_n9283, MEM_stage_inst_dmem_n9284, MEM_stage_inst_dmem_n9285, MEM_stage_inst_dmem_n9286, MEM_stage_inst_dmem_n9287, MEM_stage_inst_dmem_n9288, MEM_stage_inst_dmem_n9289, MEM_stage_inst_dmem_n9290, MEM_stage_inst_dmem_n9291, MEM_stage_inst_dmem_n9292, MEM_stage_inst_dmem_n9293, MEM_stage_inst_dmem_n9294, MEM_stage_inst_dmem_n9295, MEM_stage_inst_dmem_n9296, MEM_stage_inst_dmem_n9297, MEM_stage_inst_dmem_n9298, MEM_stage_inst_dmem_n9299, MEM_stage_inst_dmem_n9300, MEM_stage_inst_dmem_n9301, MEM_stage_inst_dmem_n9302, MEM_stage_inst_dmem_n9303, MEM_stage_inst_dmem_n9304, MEM_stage_inst_dmem_n9305, MEM_stage_inst_dmem_n9306, MEM_stage_inst_dmem_n9307, MEM_stage_inst_dmem_n9308, MEM_stage_inst_dmem_n9309, MEM_stage_inst_dmem_n9310, MEM_stage_inst_dmem_n9311, MEM_stage_inst_dmem_n9312, MEM_stage_inst_dmem_n9313, MEM_stage_inst_dmem_n9314, MEM_stage_inst_dmem_n9315, MEM_stage_inst_dmem_n9316, MEM_stage_inst_dmem_n9317, MEM_stage_inst_dmem_n9318, MEM_stage_inst_dmem_n9319, MEM_stage_inst_dmem_n9320, MEM_stage_inst_dmem_n9321, MEM_stage_inst_dmem_n9322, MEM_stage_inst_dmem_n9323, MEM_stage_inst_dmem_n9324, MEM_stage_inst_dmem_n9325, MEM_stage_inst_dmem_n9326, MEM_stage_inst_dmem_n9327, MEM_stage_inst_dmem_n9328, MEM_stage_inst_dmem_n9329, MEM_stage_inst_dmem_n9330, MEM_stage_inst_dmem_n9331, MEM_stage_inst_dmem_n9332, MEM_stage_inst_dmem_n9333, MEM_stage_inst_dmem_n9334, MEM_stage_inst_dmem_n9335, MEM_stage_inst_dmem_n9336, MEM_stage_inst_dmem_n9337, MEM_stage_inst_dmem_n9338, MEM_stage_inst_dmem_n9339, MEM_stage_inst_dmem_n9340, MEM_stage_inst_dmem_n9341, MEM_stage_inst_dmem_n9342, MEM_stage_inst_dmem_n9343, MEM_stage_inst_dmem_n9344, MEM_stage_inst_dmem_n9345, MEM_stage_inst_dmem_n9346, MEM_stage_inst_dmem_n9347, MEM_stage_inst_dmem_n9348, MEM_stage_inst_dmem_n9349, MEM_stage_inst_dmem_n9350, MEM_stage_inst_dmem_n9351, MEM_stage_inst_dmem_n9352, MEM_stage_inst_dmem_n9353, MEM_stage_inst_dmem_n9354, MEM_stage_inst_dmem_n9355, MEM_stage_inst_dmem_n9356, MEM_stage_inst_dmem_n9357, MEM_stage_inst_dmem_n9358, MEM_stage_inst_dmem_n9359, MEM_stage_inst_dmem_n9360, MEM_stage_inst_dmem_n9361, MEM_stage_inst_dmem_n9362, MEM_stage_inst_dmem_n9363, MEM_stage_inst_dmem_n9364, MEM_stage_inst_dmem_n9365, MEM_stage_inst_dmem_n9366, MEM_stage_inst_dmem_n9367, MEM_stage_inst_dmem_n9368, MEM_stage_inst_dmem_n9369, MEM_stage_inst_dmem_n9370, MEM_stage_inst_dmem_n9371, MEM_stage_inst_dmem_n9372, MEM_stage_inst_dmem_n9373, MEM_stage_inst_dmem_n9374, MEM_stage_inst_dmem_n9375, MEM_stage_inst_dmem_n9376, MEM_stage_inst_dmem_n9377, MEM_stage_inst_dmem_n9378, MEM_stage_inst_dmem_n9379, MEM_stage_inst_dmem_n9380, MEM_stage_inst_dmem_n9381, MEM_stage_inst_dmem_n9382, MEM_stage_inst_dmem_n9383, MEM_stage_inst_dmem_n9384, MEM_stage_inst_dmem_n9385, MEM_stage_inst_dmem_n9386, MEM_stage_inst_dmem_n9387, MEM_stage_inst_dmem_n9388, MEM_stage_inst_dmem_n9389, MEM_stage_inst_dmem_n9390, MEM_stage_inst_dmem_n9391, MEM_stage_inst_dmem_n9392, MEM_stage_inst_dmem_n9393, MEM_stage_inst_dmem_n9394, MEM_stage_inst_dmem_n9395, MEM_stage_inst_dmem_n9396, MEM_stage_inst_dmem_n21533, MEM_stage_inst_dmem_n9397, MEM_stage_inst_dmem_n9398, MEM_stage_inst_dmem_n9399, MEM_stage_inst_dmem_n9400, MEM_stage_inst_dmem_n9401, MEM_stage_inst_dmem_n9402, MEM_stage_inst_dmem_n21637, MEM_stage_inst_dmem_n9403, MEM_stage_inst_dmem_n9404, MEM_stage_inst_dmem_n9405, MEM_stage_inst_dmem_n9406, MEM_stage_inst_dmem_n9407, MEM_stage_inst_dmem_n9408, MEM_stage_inst_dmem_n9409, MEM_stage_inst_dmem_n9410, MEM_stage_inst_dmem_n9411, MEM_stage_inst_dmem_n9412, MEM_stage_inst_dmem_n9413, MEM_stage_inst_dmem_n9414, MEM_stage_inst_dmem_n9415, MEM_stage_inst_dmem_n9416, MEM_stage_inst_dmem_n9417, MEM_stage_inst_dmem_n9418, MEM_stage_inst_dmem_n9419, MEM_stage_inst_dmem_n9420, MEM_stage_inst_dmem_n9421, MEM_stage_inst_dmem_n9422, MEM_stage_inst_dmem_n9423, MEM_stage_inst_dmem_n9424, MEM_stage_inst_dmem_n9425, MEM_stage_inst_dmem_n9426, MEM_stage_inst_dmem_n9427, MEM_stage_inst_dmem_n9428, MEM_stage_inst_dmem_n9429, MEM_stage_inst_dmem_n9430, MEM_stage_inst_dmem_n9431, MEM_stage_inst_dmem_n9432, MEM_stage_inst_dmem_n9433, MEM_stage_inst_dmem_n9434, MEM_stage_inst_dmem_n9435, MEM_stage_inst_dmem_n9436, MEM_stage_inst_dmem_n9437, MEM_stage_inst_dmem_n9438, MEM_stage_inst_dmem_n9439, MEM_stage_inst_dmem_n9440, MEM_stage_inst_dmem_n9441, MEM_stage_inst_dmem_n9442, MEM_stage_inst_dmem_n9443, MEM_stage_inst_dmem_n9444, MEM_stage_inst_dmem_n9445, MEM_stage_inst_dmem_n9446, MEM_stage_inst_dmem_n9447, MEM_stage_inst_dmem_n9448, MEM_stage_inst_dmem_n9449, MEM_stage_inst_dmem_n9450, MEM_stage_inst_dmem_n9451, MEM_stage_inst_dmem_n9452, MEM_stage_inst_dmem_n9453, MEM_stage_inst_dmem_n9454, MEM_stage_inst_dmem_n9455, MEM_stage_inst_dmem_n9456, MEM_stage_inst_dmem_n9457, MEM_stage_inst_dmem_n9458, MEM_stage_inst_dmem_n9459, MEM_stage_inst_dmem_n9460, MEM_stage_inst_dmem_n9461, MEM_stage_inst_dmem_n9462, MEM_stage_inst_dmem_n9463, MEM_stage_inst_dmem_n9464, MEM_stage_inst_dmem_n9465, MEM_stage_inst_dmem_n9466, MEM_stage_inst_dmem_n9467, MEM_stage_inst_dmem_n9468, MEM_stage_inst_dmem_n9469, MEM_stage_inst_dmem_n9470, MEM_stage_inst_dmem_n9471, MEM_stage_inst_dmem_n9472, MEM_stage_inst_dmem_n9473, MEM_stage_inst_dmem_n9474, MEM_stage_inst_dmem_n9475, MEM_stage_inst_dmem_n9476, MEM_stage_inst_dmem_n9477, MEM_stage_inst_dmem_n9478, MEM_stage_inst_dmem_n9479, MEM_stage_inst_dmem_n9480, MEM_stage_inst_dmem_n9481, MEM_stage_inst_dmem_n9482, MEM_stage_inst_dmem_n9483, MEM_stage_inst_dmem_n9484, MEM_stage_inst_dmem_n9485, MEM_stage_inst_dmem_n9486, MEM_stage_inst_dmem_n9487, MEM_stage_inst_dmem_n9488, MEM_stage_inst_dmem_n9489, MEM_stage_inst_dmem_n9490, MEM_stage_inst_dmem_n9491, MEM_stage_inst_dmem_n9492, MEM_stage_inst_dmem_n9493, MEM_stage_inst_dmem_n9494, MEM_stage_inst_dmem_n9495, MEM_stage_inst_dmem_n9496, MEM_stage_inst_dmem_n9497, MEM_stage_inst_dmem_n21536, MEM_stage_inst_dmem_n9498, MEM_stage_inst_dmem_n9499, MEM_stage_inst_dmem_n9500, MEM_stage_inst_dmem_n9501, MEM_stage_inst_dmem_n9502, MEM_stage_inst_dmem_n9503, MEM_stage_inst_dmem_n9504, MEM_stage_inst_dmem_n9505, MEM_stage_inst_dmem_n9506, MEM_stage_inst_dmem_n9507, MEM_stage_inst_dmem_n9508, MEM_stage_inst_dmem_n9509, MEM_stage_inst_dmem_n9510, MEM_stage_inst_dmem_n9511, MEM_stage_inst_dmem_n9512, MEM_stage_inst_dmem_n9513, MEM_stage_inst_dmem_n9514, MEM_stage_inst_dmem_n9515, MEM_stage_inst_dmem_n9516, MEM_stage_inst_dmem_n9517, MEM_stage_inst_dmem_n9518, MEM_stage_inst_dmem_n9519, MEM_stage_inst_dmem_n9520, MEM_stage_inst_dmem_n9521, MEM_stage_inst_dmem_n9522, MEM_stage_inst_dmem_n9523, MEM_stage_inst_dmem_n9524, MEM_stage_inst_dmem_n9525, MEM_stage_inst_dmem_n9526, MEM_stage_inst_dmem_n9527, MEM_stage_inst_dmem_n9528, MEM_stage_inst_dmem_n9529, MEM_stage_inst_dmem_n9530, MEM_stage_inst_dmem_n9531, MEM_stage_inst_dmem_n9532, MEM_stage_inst_dmem_n9533, MEM_stage_inst_dmem_n9534, MEM_stage_inst_dmem_n9535, MEM_stage_inst_dmem_n9536, MEM_stage_inst_dmem_n9537, MEM_stage_inst_dmem_n9538, MEM_stage_inst_dmem_n9539, MEM_stage_inst_dmem_n9540, MEM_stage_inst_dmem_n9541, MEM_stage_inst_dmem_n9542, MEM_stage_inst_dmem_n9543, MEM_stage_inst_dmem_n9544, MEM_stage_inst_dmem_n9545, MEM_stage_inst_dmem_n9546, MEM_stage_inst_dmem_n9547, MEM_stage_inst_dmem_n9548, MEM_stage_inst_dmem_n9549, MEM_stage_inst_dmem_n9550, MEM_stage_inst_dmem_n9551, MEM_stage_inst_dmem_n9552, MEM_stage_inst_dmem_n9553, MEM_stage_inst_dmem_n9554, MEM_stage_inst_dmem_n9555, MEM_stage_inst_dmem_n9556, MEM_stage_inst_dmem_n9557, MEM_stage_inst_dmem_n9558, MEM_stage_inst_dmem_n9559, MEM_stage_inst_dmem_n9560, MEM_stage_inst_dmem_n9561, MEM_stage_inst_dmem_n9562, MEM_stage_inst_dmem_n9563, MEM_stage_inst_dmem_n9564, MEM_stage_inst_dmem_n9565, MEM_stage_inst_dmem_n9566, MEM_stage_inst_dmem_n9567, MEM_stage_inst_dmem_n9568, MEM_stage_inst_dmem_n9569, MEM_stage_inst_dmem_n9570, MEM_stage_inst_dmem_n9571, MEM_stage_inst_dmem_n9572, MEM_stage_inst_dmem_n9573, MEM_stage_inst_dmem_n9574, MEM_stage_inst_dmem_n9575, MEM_stage_inst_dmem_n9576, MEM_stage_inst_dmem_n9577, MEM_stage_inst_dmem_n9578, MEM_stage_inst_dmem_n9579, MEM_stage_inst_dmem_n9580, MEM_stage_inst_dmem_n9581, MEM_stage_inst_dmem_n9582, MEM_stage_inst_dmem_n9583, MEM_stage_inst_dmem_n9584, MEM_stage_inst_dmem_n9585, MEM_stage_inst_dmem_n9586, MEM_stage_inst_dmem_n9587, MEM_stage_inst_dmem_n9588, MEM_stage_inst_dmem_n9589, MEM_stage_inst_dmem_n9590, MEM_stage_inst_dmem_n9591, MEM_stage_inst_dmem_n9592, MEM_stage_inst_dmem_n9593, MEM_stage_inst_dmem_n9594, MEM_stage_inst_dmem_n9595, MEM_stage_inst_dmem_n9596, MEM_stage_inst_dmem_n9597, MEM_stage_inst_dmem_n9598, MEM_stage_inst_dmem_n9599, MEM_stage_inst_dmem_n9600, MEM_stage_inst_dmem_n9601, MEM_stage_inst_dmem_n9602, MEM_stage_inst_dmem_n9603, MEM_stage_inst_dmem_n9604, MEM_stage_inst_dmem_n9605, MEM_stage_inst_dmem_n9606, MEM_stage_inst_dmem_n9607, MEM_stage_inst_dmem_n9608, MEM_stage_inst_dmem_n9609, MEM_stage_inst_dmem_n9610, MEM_stage_inst_dmem_n9611, MEM_stage_inst_dmem_n9612, MEM_stage_inst_dmem_n9613, MEM_stage_inst_dmem_n9614, MEM_stage_inst_dmem_n9615, MEM_stage_inst_dmem_n9616, MEM_stage_inst_dmem_n9617, MEM_stage_inst_dmem_n9618, MEM_stage_inst_dmem_n9619, MEM_stage_inst_dmem_n9620, MEM_stage_inst_dmem_n9621, MEM_stage_inst_dmem_n9622, MEM_stage_inst_dmem_n9623, MEM_stage_inst_dmem_n9624, MEM_stage_inst_dmem_n9625, MEM_stage_inst_dmem_n9626, MEM_stage_inst_dmem_n9627, MEM_stage_inst_dmem_n9628, MEM_stage_inst_dmem_n9629, MEM_stage_inst_dmem_n9630, MEM_stage_inst_dmem_n9631, MEM_stage_inst_dmem_n9632, MEM_stage_inst_dmem_n9633, MEM_stage_inst_dmem_n9634, MEM_stage_inst_dmem_n9635, MEM_stage_inst_dmem_n9636, MEM_stage_inst_dmem_n9637, MEM_stage_inst_dmem_n9638, MEM_stage_inst_dmem_n9639, MEM_stage_inst_dmem_n9640, MEM_stage_inst_dmem_n9641, MEM_stage_inst_dmem_n9642, MEM_stage_inst_dmem_n9643, MEM_stage_inst_dmem_n9644, MEM_stage_inst_dmem_n9645, MEM_stage_inst_dmem_n9646, MEM_stage_inst_dmem_n9647, MEM_stage_inst_dmem_n9648, MEM_stage_inst_dmem_n9649, MEM_stage_inst_dmem_n9650, MEM_stage_inst_dmem_n9651, MEM_stage_inst_dmem_n9652, MEM_stage_inst_dmem_n9653, MEM_stage_inst_dmem_n9654, MEM_stage_inst_dmem_n9655, MEM_stage_inst_dmem_n9656, MEM_stage_inst_dmem_n9657, MEM_stage_inst_dmem_n9658, MEM_stage_inst_dmem_n9659, MEM_stage_inst_dmem_n9660, MEM_stage_inst_dmem_n9661, MEM_stage_inst_dmem_n9662, MEM_stage_inst_dmem_n9663, MEM_stage_inst_dmem_n9664, MEM_stage_inst_dmem_n9665, MEM_stage_inst_dmem_n9666, MEM_stage_inst_dmem_n9667, MEM_stage_inst_dmem_n9668, MEM_stage_inst_dmem_n9669, MEM_stage_inst_dmem_n9670, MEM_stage_inst_dmem_n9671, MEM_stage_inst_dmem_n9672, MEM_stage_inst_dmem_n9673, MEM_stage_inst_dmem_n9674, MEM_stage_inst_dmem_n9675, MEM_stage_inst_dmem_n9676, MEM_stage_inst_dmem_n9677, MEM_stage_inst_dmem_n9678, MEM_stage_inst_dmem_n9679, MEM_stage_inst_dmem_n9680, MEM_stage_inst_dmem_n9681, MEM_stage_inst_dmem_n9682, MEM_stage_inst_dmem_n9683, MEM_stage_inst_dmem_n9684, MEM_stage_inst_dmem_n9685, MEM_stage_inst_dmem_n9686, MEM_stage_inst_dmem_n9687, MEM_stage_inst_dmem_n9688, MEM_stage_inst_dmem_n9689, MEM_stage_inst_dmem_n9690, MEM_stage_inst_dmem_n9691, MEM_stage_inst_dmem_n9692, MEM_stage_inst_dmem_n9693, MEM_stage_inst_dmem_n9694, MEM_stage_inst_dmem_n9695, MEM_stage_inst_dmem_n9696, MEM_stage_inst_dmem_n9697, MEM_stage_inst_dmem_n9698, MEM_stage_inst_dmem_n9699, MEM_stage_inst_dmem_n9700, MEM_stage_inst_dmem_n9701, MEM_stage_inst_dmem_n9702, MEM_stage_inst_dmem_n9703, MEM_stage_inst_dmem_n9704, MEM_stage_inst_dmem_n9705, MEM_stage_inst_dmem_n9706, MEM_stage_inst_dmem_n9707, MEM_stage_inst_dmem_n9708, MEM_stage_inst_dmem_n9709, MEM_stage_inst_dmem_n9710, MEM_stage_inst_dmem_n9711, MEM_stage_inst_dmem_n9712, MEM_stage_inst_dmem_n9713, MEM_stage_inst_dmem_n9714, MEM_stage_inst_dmem_n9715, MEM_stage_inst_dmem_n9716, MEM_stage_inst_dmem_n9717, MEM_stage_inst_dmem_n9718, MEM_stage_inst_dmem_n9719, MEM_stage_inst_dmem_n9720, MEM_stage_inst_dmem_n9721, MEM_stage_inst_dmem_n9722, MEM_stage_inst_dmem_n9723, MEM_stage_inst_dmem_n9724, MEM_stage_inst_dmem_n9725, MEM_stage_inst_dmem_n9726, MEM_stage_inst_dmem_n9727, MEM_stage_inst_dmem_n9728, MEM_stage_inst_dmem_n9729, MEM_stage_inst_dmem_n9730, MEM_stage_inst_dmem_n9731, MEM_stage_inst_dmem_n9732, MEM_stage_inst_dmem_n9733, MEM_stage_inst_dmem_n9734, MEM_stage_inst_dmem_n9735, MEM_stage_inst_dmem_n9736, MEM_stage_inst_dmem_n9737, MEM_stage_inst_dmem_n9738, MEM_stage_inst_dmem_n9739, MEM_stage_inst_dmem_n9740, MEM_stage_inst_dmem_n9741, MEM_stage_inst_dmem_n9742, MEM_stage_inst_dmem_n9743, MEM_stage_inst_dmem_n9744, MEM_stage_inst_dmem_n9745, MEM_stage_inst_dmem_n9746, MEM_stage_inst_dmem_n9747, MEM_stage_inst_dmem_n9748, MEM_stage_inst_dmem_n9749, MEM_stage_inst_dmem_n9750, MEM_stage_inst_dmem_n9751, MEM_stage_inst_dmem_n9752, MEM_stage_inst_dmem_n9753, MEM_stage_inst_dmem_n9754, MEM_stage_inst_dmem_n9755, MEM_stage_inst_dmem_n9756, MEM_stage_inst_dmem_n9757, MEM_stage_inst_dmem_n9758, MEM_stage_inst_dmem_n9759, MEM_stage_inst_dmem_n9760, MEM_stage_inst_dmem_n9761, MEM_stage_inst_dmem_n9762, MEM_stage_inst_dmem_n9763, MEM_stage_inst_dmem_n9764, MEM_stage_inst_dmem_n9765, MEM_stage_inst_dmem_n9766, MEM_stage_inst_dmem_n9767, MEM_stage_inst_dmem_n9768, MEM_stage_inst_dmem_n9769, MEM_stage_inst_dmem_n9770, MEM_stage_inst_dmem_n9771, MEM_stage_inst_dmem_n9772, MEM_stage_inst_dmem_n9773, MEM_stage_inst_dmem_n9774, MEM_stage_inst_dmem_n9775, MEM_stage_inst_dmem_n9776, MEM_stage_inst_dmem_n9777, MEM_stage_inst_dmem_n9778, MEM_stage_inst_dmem_n9779, MEM_stage_inst_dmem_n9780, MEM_stage_inst_dmem_n9781, MEM_stage_inst_dmem_n9782, MEM_stage_inst_dmem_n9783, MEM_stage_inst_dmem_n9784, MEM_stage_inst_dmem_n9785, MEM_stage_inst_dmem_n9786, MEM_stage_inst_dmem_n9787, MEM_stage_inst_dmem_n9788, MEM_stage_inst_dmem_n9789, MEM_stage_inst_dmem_n9790, MEM_stage_inst_dmem_n9791, MEM_stage_inst_dmem_n9792, MEM_stage_inst_dmem_n9793, MEM_stage_inst_dmem_n9794, MEM_stage_inst_dmem_n9795, MEM_stage_inst_dmem_n9796, MEM_stage_inst_dmem_n9797, MEM_stage_inst_dmem_n9798, MEM_stage_inst_dmem_n9799, MEM_stage_inst_dmem_n9800, MEM_stage_inst_dmem_n9801, MEM_stage_inst_dmem_n9802, MEM_stage_inst_dmem_n9803, MEM_stage_inst_dmem_n9804, MEM_stage_inst_dmem_n9805, MEM_stage_inst_dmem_n9806, MEM_stage_inst_dmem_n9807, MEM_stage_inst_dmem_n9808, MEM_stage_inst_dmem_n9809, MEM_stage_inst_dmem_n9810, MEM_stage_inst_dmem_n9811, MEM_stage_inst_dmem_n9812, MEM_stage_inst_dmem_n9813, MEM_stage_inst_dmem_n9814, MEM_stage_inst_dmem_n9815, MEM_stage_inst_dmem_n9816, MEM_stage_inst_dmem_n9817, MEM_stage_inst_dmem_n9818, MEM_stage_inst_dmem_n9819, MEM_stage_inst_dmem_n9820, MEM_stage_inst_dmem_n9821, MEM_stage_inst_dmem_n9822, MEM_stage_inst_dmem_n9823, MEM_stage_inst_dmem_n9824, MEM_stage_inst_dmem_n9825, MEM_stage_inst_dmem_n9826, MEM_stage_inst_dmem_n9827, MEM_stage_inst_dmem_n9828, MEM_stage_inst_dmem_n9829, MEM_stage_inst_dmem_n9830, MEM_stage_inst_dmem_n9831, MEM_stage_inst_dmem_n9832, MEM_stage_inst_dmem_n9833, MEM_stage_inst_dmem_n9834, MEM_stage_inst_dmem_n9835, MEM_stage_inst_dmem_n9836, MEM_stage_inst_dmem_n9837, MEM_stage_inst_dmem_n9838, MEM_stage_inst_dmem_n9839, MEM_stage_inst_dmem_n9840, MEM_stage_inst_dmem_n9841, MEM_stage_inst_dmem_n9842, MEM_stage_inst_dmem_n9843, MEM_stage_inst_dmem_n9844, MEM_stage_inst_dmem_n9845, MEM_stage_inst_dmem_n9846, MEM_stage_inst_dmem_n9847, MEM_stage_inst_dmem_n9848, MEM_stage_inst_dmem_n9849, MEM_stage_inst_dmem_n9850, MEM_stage_inst_dmem_n9851, MEM_stage_inst_dmem_n9852, MEM_stage_inst_dmem_n9853, MEM_stage_inst_dmem_n9854, MEM_stage_inst_dmem_n9855, MEM_stage_inst_dmem_n9856, MEM_stage_inst_dmem_n9857, MEM_stage_inst_dmem_n9858, MEM_stage_inst_dmem_n9859, MEM_stage_inst_dmem_n9860, MEM_stage_inst_dmem_n9861, MEM_stage_inst_dmem_n9862, MEM_stage_inst_dmem_n9863, MEM_stage_inst_dmem_n9864, MEM_stage_inst_dmem_n9865, MEM_stage_inst_dmem_n9866, MEM_stage_inst_dmem_n9867, MEM_stage_inst_dmem_n9868, MEM_stage_inst_dmem_n9869, MEM_stage_inst_dmem_n9870, MEM_stage_inst_dmem_n9871, MEM_stage_inst_dmem_n9872, MEM_stage_inst_dmem_n9873, MEM_stage_inst_dmem_n9874, MEM_stage_inst_dmem_n9875, MEM_stage_inst_dmem_n9876, MEM_stage_inst_dmem_n9877, MEM_stage_inst_dmem_n9878, MEM_stage_inst_dmem_n9879, MEM_stage_inst_dmem_n9880, MEM_stage_inst_dmem_n9881, MEM_stage_inst_dmem_n9882, MEM_stage_inst_dmem_n9883, MEM_stage_inst_dmem_n9884, MEM_stage_inst_dmem_n9885, MEM_stage_inst_dmem_n9886, MEM_stage_inst_dmem_n9887, MEM_stage_inst_dmem_n9888, MEM_stage_inst_dmem_n9889, MEM_stage_inst_dmem_n9890, MEM_stage_inst_dmem_n9891, MEM_stage_inst_dmem_n9892, MEM_stage_inst_dmem_n9893, MEM_stage_inst_dmem_n9894, MEM_stage_inst_dmem_n9895, MEM_stage_inst_dmem_n9896, MEM_stage_inst_dmem_n9897, MEM_stage_inst_dmem_n9898, MEM_stage_inst_dmem_n9899, MEM_stage_inst_dmem_n9900, MEM_stage_inst_dmem_n9901, MEM_stage_inst_dmem_n9902, MEM_stage_inst_dmem_n9903, MEM_stage_inst_dmem_n9904, MEM_stage_inst_dmem_n9905, MEM_stage_inst_dmem_n9906, MEM_stage_inst_dmem_n9907, MEM_stage_inst_dmem_n9908, MEM_stage_inst_dmem_n9909, MEM_stage_inst_dmem_n9910, MEM_stage_inst_dmem_n9911, MEM_stage_inst_dmem_n9912, MEM_stage_inst_dmem_n9913, MEM_stage_inst_dmem_n9914, MEM_stage_inst_dmem_n9915, MEM_stage_inst_dmem_n9916, MEM_stage_inst_dmem_n9917, MEM_stage_inst_dmem_n9918, MEM_stage_inst_dmem_n9919, MEM_stage_inst_dmem_n9920, MEM_stage_inst_dmem_n9921, MEM_stage_inst_dmem_n9922, MEM_stage_inst_dmem_n9923, MEM_stage_inst_dmem_n9924, MEM_stage_inst_dmem_n9925, MEM_stage_inst_dmem_n9926, MEM_stage_inst_dmem_n9927, MEM_stage_inst_dmem_n9928, MEM_stage_inst_dmem_n9929, MEM_stage_inst_dmem_n9930, MEM_stage_inst_dmem_n9931, MEM_stage_inst_dmem_n9932, MEM_stage_inst_dmem_n9933, MEM_stage_inst_dmem_n9934, MEM_stage_inst_dmem_n9935, MEM_stage_inst_dmem_n9936, MEM_stage_inst_dmem_n9937, MEM_stage_inst_dmem_n9938, MEM_stage_inst_dmem_n9939, MEM_stage_inst_dmem_n9940, MEM_stage_inst_dmem_n9941, MEM_stage_inst_dmem_n9942, MEM_stage_inst_dmem_n9943, MEM_stage_inst_dmem_n9944, MEM_stage_inst_dmem_n9945, MEM_stage_inst_dmem_n9946, MEM_stage_inst_dmem_n9947, MEM_stage_inst_dmem_n9948, MEM_stage_inst_dmem_n9949, MEM_stage_inst_dmem_n9950, MEM_stage_inst_dmem_n9951, MEM_stage_inst_dmem_n9952, MEM_stage_inst_dmem_n9953, MEM_stage_inst_dmem_n9954, MEM_stage_inst_dmem_n9955, MEM_stage_inst_dmem_n9956, MEM_stage_inst_dmem_n9957, MEM_stage_inst_dmem_n9958, MEM_stage_inst_dmem_n9959, MEM_stage_inst_dmem_n9960, MEM_stage_inst_dmem_n9961, MEM_stage_inst_dmem_n9962, MEM_stage_inst_dmem_n9963, MEM_stage_inst_dmem_n9964, MEM_stage_inst_dmem_n9965, MEM_stage_inst_dmem_n9966, MEM_stage_inst_dmem_n9967, MEM_stage_inst_dmem_n9968, MEM_stage_inst_dmem_n9969, MEM_stage_inst_dmem_n9970, MEM_stage_inst_dmem_n9971, MEM_stage_inst_dmem_n9972, MEM_stage_inst_dmem_n9973, MEM_stage_inst_dmem_n9974, MEM_stage_inst_dmem_n9975, MEM_stage_inst_dmem_n9976, MEM_stage_inst_dmem_n9977, MEM_stage_inst_dmem_n9978, MEM_stage_inst_dmem_n9979, MEM_stage_inst_dmem_n9980, MEM_stage_inst_dmem_n9981, MEM_stage_inst_dmem_n9982, MEM_stage_inst_dmem_n9983, MEM_stage_inst_dmem_n9984, MEM_stage_inst_dmem_n9985, MEM_stage_inst_dmem_n9986, MEM_stage_inst_dmem_n9987, MEM_stage_inst_dmem_n9988, MEM_stage_inst_dmem_n9989, MEM_stage_inst_dmem_n9990, MEM_stage_inst_dmem_n9991, MEM_stage_inst_dmem_n9992, MEM_stage_inst_dmem_n9993, MEM_stage_inst_dmem_n9994, MEM_stage_inst_dmem_n9995, MEM_stage_inst_dmem_n9996, MEM_stage_inst_dmem_n9997, MEM_stage_inst_dmem_n9998, MEM_stage_inst_dmem_n9999, MEM_stage_inst_dmem_n10000, MEM_stage_inst_dmem_n10001, MEM_stage_inst_dmem_n10002, MEM_stage_inst_dmem_n10003, MEM_stage_inst_dmem_n10004, MEM_stage_inst_dmem_n10005, MEM_stage_inst_dmem_n10006, MEM_stage_inst_dmem_n10007, MEM_stage_inst_dmem_n10008, MEM_stage_inst_dmem_n10009, MEM_stage_inst_dmem_n10010, MEM_stage_inst_dmem_n10011, MEM_stage_inst_dmem_n10012, MEM_stage_inst_dmem_n10013, MEM_stage_inst_dmem_n10014, MEM_stage_inst_dmem_n10015, MEM_stage_inst_dmem_n10016, MEM_stage_inst_dmem_n10017, MEM_stage_inst_dmem_n10018, MEM_stage_inst_dmem_n10019, MEM_stage_inst_dmem_n10020, MEM_stage_inst_dmem_n10021, MEM_stage_inst_dmem_n10022, MEM_stage_inst_dmem_n10023, MEM_stage_inst_dmem_n10024, MEM_stage_inst_dmem_n10025, MEM_stage_inst_dmem_n10026, MEM_stage_inst_dmem_n10027, MEM_stage_inst_dmem_n10028, MEM_stage_inst_dmem_n10029, MEM_stage_inst_dmem_n10030, MEM_stage_inst_dmem_n10031, MEM_stage_inst_dmem_n10032, MEM_stage_inst_dmem_n10033, MEM_stage_inst_dmem_n10034, MEM_stage_inst_dmem_n10035, MEM_stage_inst_dmem_n10036, MEM_stage_inst_dmem_n10037, MEM_stage_inst_dmem_n10038, MEM_stage_inst_dmem_n10039, MEM_stage_inst_dmem_n10040, MEM_stage_inst_dmem_n10041, MEM_stage_inst_dmem_n10042, MEM_stage_inst_dmem_n10043, MEM_stage_inst_dmem_n10044, MEM_stage_inst_dmem_n10045, MEM_stage_inst_dmem_n10046, MEM_stage_inst_dmem_n10047, MEM_stage_inst_dmem_n10048, MEM_stage_inst_dmem_n10049, MEM_stage_inst_dmem_n10050, MEM_stage_inst_dmem_n10051, MEM_stage_inst_dmem_n10052, MEM_stage_inst_dmem_n10053, MEM_stage_inst_dmem_n10054, MEM_stage_inst_dmem_n10055, MEM_stage_inst_dmem_n10056, MEM_stage_inst_dmem_n10057, MEM_stage_inst_dmem_n10058, MEM_stage_inst_dmem_n10059, MEM_stage_inst_dmem_n10060, MEM_stage_inst_dmem_n10061, MEM_stage_inst_dmem_n10062, MEM_stage_inst_dmem_n10063, MEM_stage_inst_dmem_n10064, MEM_stage_inst_dmem_n10065, MEM_stage_inst_dmem_n10066, MEM_stage_inst_dmem_n10067, MEM_stage_inst_dmem_n10068, MEM_stage_inst_dmem_n10069, MEM_stage_inst_dmem_n10070, MEM_stage_inst_dmem_n10071, MEM_stage_inst_dmem_n10072, MEM_stage_inst_dmem_n10073, MEM_stage_inst_dmem_n10074, MEM_stage_inst_dmem_n10075, MEM_stage_inst_dmem_n10076, MEM_stage_inst_dmem_n10077, MEM_stage_inst_dmem_n10078, MEM_stage_inst_dmem_n10079, MEM_stage_inst_dmem_n10080, MEM_stage_inst_dmem_n10081, MEM_stage_inst_dmem_n10082, MEM_stage_inst_dmem_n10083, MEM_stage_inst_dmem_n10084, MEM_stage_inst_dmem_n10085, MEM_stage_inst_dmem_n10086, MEM_stage_inst_dmem_n10087, MEM_stage_inst_dmem_n10088, MEM_stage_inst_dmem_n10089, MEM_stage_inst_dmem_n10090, MEM_stage_inst_dmem_n10091, MEM_stage_inst_dmem_n10092, MEM_stage_inst_dmem_n10093, MEM_stage_inst_dmem_n10094, MEM_stage_inst_dmem_n10095, MEM_stage_inst_dmem_n10096, MEM_stage_inst_dmem_n10097, MEM_stage_inst_dmem_n10098, MEM_stage_inst_dmem_n10099, MEM_stage_inst_dmem_n10100, MEM_stage_inst_dmem_n10101, MEM_stage_inst_dmem_n10102, MEM_stage_inst_dmem_n10103, MEM_stage_inst_dmem_n10104, MEM_stage_inst_dmem_n10105, MEM_stage_inst_dmem_n10106, MEM_stage_inst_dmem_n10107, MEM_stage_inst_dmem_n10108, MEM_stage_inst_dmem_n10109, MEM_stage_inst_dmem_n10110, MEM_stage_inst_dmem_n10111, MEM_stage_inst_dmem_n10112, MEM_stage_inst_dmem_n10113, MEM_stage_inst_dmem_n10114, MEM_stage_inst_dmem_n10115, MEM_stage_inst_dmem_n10116, MEM_stage_inst_dmem_n10117, MEM_stage_inst_dmem_n10118, MEM_stage_inst_dmem_n10119, MEM_stage_inst_dmem_n10120, MEM_stage_inst_dmem_n10121, MEM_stage_inst_dmem_n10122, MEM_stage_inst_dmem_n10123, MEM_stage_inst_dmem_n10124, MEM_stage_inst_dmem_n10125, MEM_stage_inst_dmem_n10126, MEM_stage_inst_dmem_n10127, MEM_stage_inst_dmem_n10128, MEM_stage_inst_dmem_n10129, MEM_stage_inst_dmem_n10130, MEM_stage_inst_dmem_n10131, MEM_stage_inst_dmem_n10132, MEM_stage_inst_dmem_n10133, MEM_stage_inst_dmem_n10134, MEM_stage_inst_dmem_n10135, MEM_stage_inst_dmem_n10136, MEM_stage_inst_dmem_n10137, MEM_stage_inst_dmem_n10138, MEM_stage_inst_dmem_n10139, MEM_stage_inst_dmem_n10140, MEM_stage_inst_dmem_n10141, MEM_stage_inst_dmem_n10142, MEM_stage_inst_dmem_n10143, MEM_stage_inst_dmem_n10144, MEM_stage_inst_dmem_n10145, MEM_stage_inst_dmem_n10146, MEM_stage_inst_dmem_n10147, MEM_stage_inst_dmem_n10148, MEM_stage_inst_dmem_n10149, MEM_stage_inst_dmem_n10150, MEM_stage_inst_dmem_n10151, MEM_stage_inst_dmem_n10152, MEM_stage_inst_dmem_n10153, MEM_stage_inst_dmem_n10154, MEM_stage_inst_dmem_n10155, MEM_stage_inst_dmem_n10156, MEM_stage_inst_dmem_n10157, MEM_stage_inst_dmem_n10158, MEM_stage_inst_dmem_n10159, MEM_stage_inst_dmem_n10160, MEM_stage_inst_dmem_n10161, MEM_stage_inst_dmem_n10162, MEM_stage_inst_dmem_n10163, MEM_stage_inst_dmem_n10164, MEM_stage_inst_dmem_n10165, MEM_stage_inst_dmem_n10166, MEM_stage_inst_dmem_n10167, MEM_stage_inst_dmem_n10168, MEM_stage_inst_dmem_n10169, MEM_stage_inst_dmem_n10170, MEM_stage_inst_dmem_n10171, MEM_stage_inst_dmem_n10172, MEM_stage_inst_dmem_n10173, MEM_stage_inst_dmem_n10174, MEM_stage_inst_dmem_n10175, MEM_stage_inst_dmem_n10176, MEM_stage_inst_dmem_n10177, MEM_stage_inst_dmem_n10178, MEM_stage_inst_dmem_n10179, MEM_stage_inst_dmem_n10180, MEM_stage_inst_dmem_n10181, MEM_stage_inst_dmem_n10182, MEM_stage_inst_dmem_n10183, MEM_stage_inst_dmem_n10184, MEM_stage_inst_dmem_n10185, MEM_stage_inst_dmem_n10186, MEM_stage_inst_dmem_n10187, MEM_stage_inst_dmem_n10188, MEM_stage_inst_dmem_n10189, MEM_stage_inst_dmem_n10190, MEM_stage_inst_dmem_n10191, MEM_stage_inst_dmem_n10192, MEM_stage_inst_dmem_n10193, MEM_stage_inst_dmem_n10194, MEM_stage_inst_dmem_n10195, MEM_stage_inst_dmem_n10196, MEM_stage_inst_dmem_n10197, MEM_stage_inst_dmem_n10198, MEM_stage_inst_dmem_n10199, MEM_stage_inst_dmem_n10200, MEM_stage_inst_dmem_n10201, MEM_stage_inst_dmem_n10202, MEM_stage_inst_dmem_n10203, MEM_stage_inst_dmem_n10204, MEM_stage_inst_dmem_n10205, MEM_stage_inst_dmem_n10206, MEM_stage_inst_dmem_n10207, MEM_stage_inst_dmem_n10208, MEM_stage_inst_dmem_n10209, MEM_stage_inst_dmem_n10210, MEM_stage_inst_dmem_n10211, MEM_stage_inst_dmem_n10212, MEM_stage_inst_dmem_n10213, MEM_stage_inst_dmem_n10214, MEM_stage_inst_dmem_n10215, MEM_stage_inst_dmem_n10216, MEM_stage_inst_dmem_n10217, MEM_stage_inst_dmem_n10218, MEM_stage_inst_dmem_n10219, MEM_stage_inst_dmem_n10220, MEM_stage_inst_dmem_n10221, MEM_stage_inst_dmem_n10222, MEM_stage_inst_dmem_n10223, MEM_stage_inst_dmem_n10224, MEM_stage_inst_dmem_n10225, MEM_stage_inst_dmem_n10226, MEM_stage_inst_dmem_n10227, MEM_stage_inst_dmem_n10228, MEM_stage_inst_dmem_n10229, MEM_stage_inst_dmem_n10230, MEM_stage_inst_dmem_n10231, MEM_stage_inst_dmem_n10232, MEM_stage_inst_dmem_n10233, MEM_stage_inst_dmem_n10234, MEM_stage_inst_dmem_n10235, MEM_stage_inst_dmem_n10236, MEM_stage_inst_dmem_n10237, MEM_stage_inst_dmem_n10238, MEM_stage_inst_dmem_n10239, MEM_stage_inst_dmem_n10240, MEM_stage_inst_dmem_n10241, MEM_stage_inst_dmem_n10242, MEM_stage_inst_dmem_n10243, MEM_stage_inst_dmem_n10244, MEM_stage_inst_dmem_n10245, MEM_stage_inst_dmem_n10246, MEM_stage_inst_dmem_n10247, MEM_stage_inst_dmem_n10248, MEM_stage_inst_dmem_n10249, MEM_stage_inst_dmem_n10250, MEM_stage_inst_dmem_n10251, MEM_stage_inst_dmem_n10252, MEM_stage_inst_dmem_n10253, MEM_stage_inst_dmem_n10254, MEM_stage_inst_dmem_n10255, MEM_stage_inst_dmem_n10256, MEM_stage_inst_dmem_n10257, MEM_stage_inst_dmem_n10258, MEM_stage_inst_dmem_n10259, MEM_stage_inst_dmem_n10260, MEM_stage_inst_dmem_n10261, MEM_stage_inst_dmem_n10262, MEM_stage_inst_dmem_n10263, MEM_stage_inst_dmem_n10264, MEM_stage_inst_dmem_n10265, MEM_stage_inst_dmem_n10266, MEM_stage_inst_dmem_n10267, MEM_stage_inst_dmem_n10268, MEM_stage_inst_dmem_n10269, MEM_stage_inst_dmem_n10270, MEM_stage_inst_dmem_n10271, MEM_stage_inst_dmem_n10272, MEM_stage_inst_dmem_n10273, MEM_stage_inst_dmem_n10274, MEM_stage_inst_dmem_n10275, MEM_stage_inst_dmem_n10276, MEM_stage_inst_dmem_n10277, MEM_stage_inst_dmem_n10278, MEM_stage_inst_dmem_n10279, MEM_stage_inst_dmem_n10280, MEM_stage_inst_dmem_n10281, MEM_stage_inst_dmem_n10282, MEM_stage_inst_dmem_n10283, MEM_stage_inst_dmem_n10284, MEM_stage_inst_dmem_n10285, MEM_stage_inst_dmem_n10286, MEM_stage_inst_dmem_n10287, MEM_stage_inst_dmem_n10288, MEM_stage_inst_dmem_n10289, MEM_stage_inst_dmem_n10290, MEM_stage_inst_dmem_n10291, MEM_stage_inst_dmem_n10292, MEM_stage_inst_dmem_n10293, MEM_stage_inst_dmem_n10294, MEM_stage_inst_dmem_n10295, MEM_stage_inst_dmem_n10296, MEM_stage_inst_dmem_n10297, MEM_stage_inst_dmem_n10298, MEM_stage_inst_dmem_n10299, MEM_stage_inst_dmem_n10300, MEM_stage_inst_dmem_n10301, MEM_stage_inst_dmem_n10302, MEM_stage_inst_dmem_n10303, MEM_stage_inst_dmem_n10304, MEM_stage_inst_dmem_n10305, MEM_stage_inst_dmem_n10306, MEM_stage_inst_dmem_n10307, MEM_stage_inst_dmem_n10308, MEM_stage_inst_dmem_n10309, MEM_stage_inst_dmem_n10310, MEM_stage_inst_dmem_n10311, MEM_stage_inst_dmem_n10312, MEM_stage_inst_dmem_n10313, MEM_stage_inst_dmem_n10314, MEM_stage_inst_dmem_n10315, MEM_stage_inst_dmem_n10316, MEM_stage_inst_dmem_n10317, MEM_stage_inst_dmem_n10318, MEM_stage_inst_dmem_n10319, MEM_stage_inst_dmem_n10320, MEM_stage_inst_dmem_n10321, MEM_stage_inst_dmem_n10322, MEM_stage_inst_dmem_n10323, MEM_stage_inst_dmem_n10324, MEM_stage_inst_dmem_n10325, MEM_stage_inst_dmem_n10326, MEM_stage_inst_dmem_n10327, MEM_stage_inst_dmem_n10328, MEM_stage_inst_dmem_n10329, MEM_stage_inst_dmem_n10330, MEM_stage_inst_dmem_n10331, MEM_stage_inst_dmem_n10332, MEM_stage_inst_dmem_n10333, MEM_stage_inst_dmem_n10334, MEM_stage_inst_dmem_n10335, MEM_stage_inst_dmem_n10336, MEM_stage_inst_dmem_n10337, MEM_stage_inst_dmem_n10338, MEM_stage_inst_dmem_n10339, MEM_stage_inst_dmem_n10340, MEM_stage_inst_dmem_n10341, MEM_stage_inst_dmem_n10342, MEM_stage_inst_dmem_n10343, MEM_stage_inst_dmem_n10344, MEM_stage_inst_dmem_n10345, MEM_stage_inst_dmem_n10346, MEM_stage_inst_dmem_n10347, MEM_stage_inst_dmem_n10348, MEM_stage_inst_dmem_n10349, MEM_stage_inst_dmem_n10350, MEM_stage_inst_dmem_n10351, MEM_stage_inst_dmem_n10352, MEM_stage_inst_dmem_n10353, MEM_stage_inst_dmem_n10354, MEM_stage_inst_dmem_n10355, MEM_stage_inst_dmem_n10356, MEM_stage_inst_dmem_n10357, MEM_stage_inst_dmem_n10358, MEM_stage_inst_dmem_n10359, MEM_stage_inst_dmem_n10360, MEM_stage_inst_dmem_n10361, MEM_stage_inst_dmem_n10362, MEM_stage_inst_dmem_n10363, MEM_stage_inst_dmem_n10364, MEM_stage_inst_dmem_n10365, MEM_stage_inst_dmem_n10366, MEM_stage_inst_dmem_n10367, MEM_stage_inst_dmem_n10368, MEM_stage_inst_dmem_n10369, MEM_stage_inst_dmem_n10370, MEM_stage_inst_dmem_n10371, MEM_stage_inst_dmem_n10372, MEM_stage_inst_dmem_n10373, MEM_stage_inst_dmem_n10374, MEM_stage_inst_dmem_n10375, MEM_stage_inst_dmem_n10376, MEM_stage_inst_dmem_n10377, MEM_stage_inst_dmem_n10378, MEM_stage_inst_dmem_n10379, MEM_stage_inst_dmem_n10380, MEM_stage_inst_dmem_n10381, MEM_stage_inst_dmem_n10382, MEM_stage_inst_dmem_n10383, MEM_stage_inst_dmem_n10384, MEM_stage_inst_dmem_n10385, MEM_stage_inst_dmem_n10386, MEM_stage_inst_dmem_n10387, MEM_stage_inst_dmem_n10388, MEM_stage_inst_dmem_n10389, MEM_stage_inst_dmem_n10390, MEM_stage_inst_dmem_n10391, MEM_stage_inst_dmem_n10392, MEM_stage_inst_dmem_n10393, MEM_stage_inst_dmem_n10394, MEM_stage_inst_dmem_n10395, MEM_stage_inst_dmem_n10396, MEM_stage_inst_dmem_n10397, MEM_stage_inst_dmem_n10398, MEM_stage_inst_dmem_n10399, MEM_stage_inst_dmem_n10400, MEM_stage_inst_dmem_n10401, MEM_stage_inst_dmem_n10402, MEM_stage_inst_dmem_n10403, MEM_stage_inst_dmem_n10404, MEM_stage_inst_dmem_n10405, MEM_stage_inst_dmem_n10406, MEM_stage_inst_dmem_n10407, MEM_stage_inst_dmem_n10408, MEM_stage_inst_dmem_n10409, MEM_stage_inst_dmem_n10410, MEM_stage_inst_dmem_n10411, MEM_stage_inst_dmem_n10412, MEM_stage_inst_dmem_n10413, MEM_stage_inst_dmem_n10414, MEM_stage_inst_dmem_n10415, MEM_stage_inst_dmem_n10416, MEM_stage_inst_dmem_n10417, MEM_stage_inst_dmem_n10418, MEM_stage_inst_dmem_n10419, MEM_stage_inst_dmem_n10420, MEM_stage_inst_dmem_n10421, MEM_stage_inst_dmem_n10422, MEM_stage_inst_dmem_n10423, MEM_stage_inst_dmem_n10424, MEM_stage_inst_dmem_n10425, MEM_stage_inst_dmem_n10426, MEM_stage_inst_dmem_n10427, MEM_stage_inst_dmem_n10428, MEM_stage_inst_dmem_n10429, MEM_stage_inst_dmem_n10430, MEM_stage_inst_dmem_n10431, MEM_stage_inst_dmem_n10432, MEM_stage_inst_dmem_n10433, MEM_stage_inst_dmem_n10434, MEM_stage_inst_dmem_n10435, MEM_stage_inst_dmem_n10436, MEM_stage_inst_dmem_n10437, MEM_stage_inst_dmem_n10438, MEM_stage_inst_dmem_n10439, MEM_stage_inst_dmem_n10440, MEM_stage_inst_dmem_n10441, MEM_stage_inst_dmem_n10442, MEM_stage_inst_dmem_n10443, MEM_stage_inst_dmem_n10444, MEM_stage_inst_dmem_n10445, MEM_stage_inst_dmem_n10446, MEM_stage_inst_dmem_n10447, MEM_stage_inst_dmem_n10448, MEM_stage_inst_dmem_n10449, MEM_stage_inst_dmem_n10450, MEM_stage_inst_dmem_n10451, MEM_stage_inst_dmem_n10452, MEM_stage_inst_dmem_n10453, MEM_stage_inst_dmem_n10454, MEM_stage_inst_dmem_n10455, MEM_stage_inst_dmem_n10456, MEM_stage_inst_dmem_n10457, MEM_stage_inst_dmem_n10458, MEM_stage_inst_dmem_n10459, MEM_stage_inst_dmem_n10460, MEM_stage_inst_dmem_n10461, MEM_stage_inst_dmem_n10462, MEM_stage_inst_dmem_n10463, MEM_stage_inst_dmem_n10464, MEM_stage_inst_dmem_n10465, MEM_stage_inst_dmem_n10466, MEM_stage_inst_dmem_n10467, MEM_stage_inst_dmem_n10468, MEM_stage_inst_dmem_n10469, MEM_stage_inst_dmem_n10470, MEM_stage_inst_dmem_n10471, MEM_stage_inst_dmem_n10472, MEM_stage_inst_dmem_n10473, MEM_stage_inst_dmem_n10474, MEM_stage_inst_dmem_n10475, MEM_stage_inst_dmem_n10476, MEM_stage_inst_dmem_n10477, MEM_stage_inst_dmem_n10478, MEM_stage_inst_dmem_n10479, MEM_stage_inst_dmem_n10480, MEM_stage_inst_dmem_n10481, MEM_stage_inst_dmem_n10482, MEM_stage_inst_dmem_n10483, MEM_stage_inst_dmem_n10484, MEM_stage_inst_dmem_n10485, MEM_stage_inst_dmem_n10486, MEM_stage_inst_dmem_n10487, MEM_stage_inst_dmem_n10488, MEM_stage_inst_dmem_n10489, MEM_stage_inst_dmem_n10490, MEM_stage_inst_dmem_n10491, MEM_stage_inst_dmem_n10492, MEM_stage_inst_dmem_n10493, MEM_stage_inst_dmem_n10494, MEM_stage_inst_dmem_n10495, MEM_stage_inst_dmem_n10496, MEM_stage_inst_dmem_n10497, MEM_stage_inst_dmem_n10498, MEM_stage_inst_dmem_n10499, MEM_stage_inst_dmem_n10500, MEM_stage_inst_dmem_n10501, MEM_stage_inst_dmem_n10502, MEM_stage_inst_dmem_n10503, MEM_stage_inst_dmem_n10504, MEM_stage_inst_dmem_n10505, MEM_stage_inst_dmem_n10506, MEM_stage_inst_dmem_n10507, MEM_stage_inst_dmem_n10508, MEM_stage_inst_dmem_n10509, MEM_stage_inst_dmem_n10510, MEM_stage_inst_dmem_n10511, MEM_stage_inst_dmem_n10512, MEM_stage_inst_dmem_n10513, MEM_stage_inst_dmem_n10514, MEM_stage_inst_dmem_n10515, MEM_stage_inst_dmem_n10516, MEM_stage_inst_dmem_n10517, MEM_stage_inst_dmem_n10518, MEM_stage_inst_dmem_n10519, MEM_stage_inst_dmem_n10520, MEM_stage_inst_dmem_n10521, MEM_stage_inst_dmem_n10522, MEM_stage_inst_dmem_n10523, MEM_stage_inst_dmem_n10524, MEM_stage_inst_dmem_n10525, MEM_stage_inst_dmem_n10526, MEM_stage_inst_dmem_n10527, MEM_stage_inst_dmem_n10528, MEM_stage_inst_dmem_n10529, MEM_stage_inst_dmem_n10530, MEM_stage_inst_dmem_n10531, MEM_stage_inst_dmem_n10532, MEM_stage_inst_dmem_n10533, MEM_stage_inst_dmem_n10534, MEM_stage_inst_dmem_n10535, MEM_stage_inst_dmem_n10536, MEM_stage_inst_dmem_n10537, MEM_stage_inst_dmem_n10538, MEM_stage_inst_dmem_n10539, MEM_stage_inst_dmem_n10540, MEM_stage_inst_dmem_n10541, MEM_stage_inst_dmem_n10542, MEM_stage_inst_dmem_n10543, MEM_stage_inst_dmem_n10544, MEM_stage_inst_dmem_n10545, MEM_stage_inst_dmem_n10546, MEM_stage_inst_dmem_n10547, MEM_stage_inst_dmem_n10548, MEM_stage_inst_dmem_n10549, MEM_stage_inst_dmem_n10550, MEM_stage_inst_dmem_n10551, MEM_stage_inst_dmem_n10552, MEM_stage_inst_dmem_n10553, MEM_stage_inst_dmem_n10554, MEM_stage_inst_dmem_n10555, MEM_stage_inst_dmem_n10556, MEM_stage_inst_dmem_n10557, MEM_stage_inst_dmem_n10558, MEM_stage_inst_dmem_n10559, MEM_stage_inst_dmem_n10560, MEM_stage_inst_dmem_n10561, MEM_stage_inst_dmem_n10562, MEM_stage_inst_dmem_n10563, MEM_stage_inst_dmem_n10564, MEM_stage_inst_dmem_n10565, MEM_stage_inst_dmem_n10566, MEM_stage_inst_dmem_n10567, MEM_stage_inst_dmem_n10568, MEM_stage_inst_dmem_n10569, MEM_stage_inst_dmem_n10570, MEM_stage_inst_dmem_n10571, MEM_stage_inst_dmem_n10572, MEM_stage_inst_dmem_n10573, MEM_stage_inst_dmem_n10574, MEM_stage_inst_dmem_n10575, MEM_stage_inst_dmem_n10576, MEM_stage_inst_dmem_n10577, MEM_stage_inst_dmem_n10578, MEM_stage_inst_dmem_n10579, MEM_stage_inst_dmem_n10580, MEM_stage_inst_dmem_n10581, MEM_stage_inst_dmem_n10582, MEM_stage_inst_dmem_n10583, MEM_stage_inst_dmem_n10584, MEM_stage_inst_dmem_n10585, MEM_stage_inst_dmem_n10586, MEM_stage_inst_dmem_n10587, MEM_stage_inst_dmem_n10588, MEM_stage_inst_dmem_n10589, MEM_stage_inst_dmem_n10590, MEM_stage_inst_dmem_n10591, MEM_stage_inst_dmem_n10592, MEM_stage_inst_dmem_n10593, MEM_stage_inst_dmem_n10594, MEM_stage_inst_dmem_n10595, MEM_stage_inst_dmem_n10596, MEM_stage_inst_dmem_n10597, MEM_stage_inst_dmem_n10598, MEM_stage_inst_dmem_n10599, MEM_stage_inst_dmem_n10600, MEM_stage_inst_dmem_n10601, MEM_stage_inst_dmem_n10602, MEM_stage_inst_dmem_n10603, MEM_stage_inst_dmem_n10604, MEM_stage_inst_dmem_n10605, MEM_stage_inst_dmem_n10606, MEM_stage_inst_dmem_n10607, MEM_stage_inst_dmem_n10608, MEM_stage_inst_dmem_n10609, MEM_stage_inst_dmem_n10610, MEM_stage_inst_dmem_n10611, MEM_stage_inst_dmem_n10612, MEM_stage_inst_dmem_n10613, MEM_stage_inst_dmem_n10614, MEM_stage_inst_dmem_n10615, MEM_stage_inst_dmem_n10616, MEM_stage_inst_dmem_n10617, MEM_stage_inst_dmem_n10618, MEM_stage_inst_dmem_n10619, MEM_stage_inst_dmem_n10620, MEM_stage_inst_dmem_n10621, MEM_stage_inst_dmem_n10622, MEM_stage_inst_dmem_n10623, MEM_stage_inst_dmem_n10624, MEM_stage_inst_dmem_n10625, MEM_stage_inst_dmem_n10626, MEM_stage_inst_dmem_n10627, MEM_stage_inst_dmem_n10628, MEM_stage_inst_dmem_n10629, MEM_stage_inst_dmem_n10630, MEM_stage_inst_dmem_n10631, MEM_stage_inst_dmem_n10632, MEM_stage_inst_dmem_n10633, MEM_stage_inst_dmem_n10634, MEM_stage_inst_dmem_n10635, MEM_stage_inst_dmem_n10636, MEM_stage_inst_dmem_n10637, MEM_stage_inst_dmem_n10638, MEM_stage_inst_dmem_n10639, MEM_stage_inst_dmem_n10640, MEM_stage_inst_dmem_n10641, MEM_stage_inst_dmem_n10642, MEM_stage_inst_dmem_n10643, MEM_stage_inst_dmem_n10644, MEM_stage_inst_dmem_n10645, MEM_stage_inst_dmem_n10646, MEM_stage_inst_dmem_n10647, MEM_stage_inst_dmem_n10648, MEM_stage_inst_dmem_n10649, MEM_stage_inst_dmem_n10650, MEM_stage_inst_dmem_n10651, MEM_stage_inst_dmem_n10652, MEM_stage_inst_dmem_n10653, MEM_stage_inst_dmem_n10654, MEM_stage_inst_dmem_n10655, MEM_stage_inst_dmem_n10656, MEM_stage_inst_dmem_n10657, MEM_stage_inst_dmem_n10658, MEM_stage_inst_dmem_n10659, MEM_stage_inst_dmem_n10660, MEM_stage_inst_dmem_n10661, MEM_stage_inst_dmem_n10662, MEM_stage_inst_dmem_n10663, MEM_stage_inst_dmem_n10664, MEM_stage_inst_dmem_n10665, MEM_stage_inst_dmem_n10666, MEM_stage_inst_dmem_n10667, MEM_stage_inst_dmem_n10668, MEM_stage_inst_dmem_n10669, MEM_stage_inst_dmem_n10670, MEM_stage_inst_dmem_n10671, MEM_stage_inst_dmem_n10672, MEM_stage_inst_dmem_n10673, MEM_stage_inst_dmem_n10674, MEM_stage_inst_dmem_n10675, MEM_stage_inst_dmem_n10676, MEM_stage_inst_dmem_n10677, MEM_stage_inst_dmem_n10678, MEM_stage_inst_dmem_n10679, MEM_stage_inst_dmem_n10680, MEM_stage_inst_dmem_n10681, MEM_stage_inst_dmem_n10682, MEM_stage_inst_dmem_n10683, MEM_stage_inst_dmem_n10684, MEM_stage_inst_dmem_n10685, MEM_stage_inst_dmem_n10686, MEM_stage_inst_dmem_n10687, MEM_stage_inst_dmem_n10688, MEM_stage_inst_dmem_n10689, MEM_stage_inst_dmem_n10690, MEM_stage_inst_dmem_n10691, MEM_stage_inst_dmem_n10692, MEM_stage_inst_dmem_n10693, MEM_stage_inst_dmem_n10694, MEM_stage_inst_dmem_n10695, MEM_stage_inst_dmem_n10696, MEM_stage_inst_dmem_n10697, MEM_stage_inst_dmem_n10698, MEM_stage_inst_dmem_n10699, MEM_stage_inst_dmem_n10700, MEM_stage_inst_dmem_n10701, MEM_stage_inst_dmem_n10702, MEM_stage_inst_dmem_n10703, MEM_stage_inst_dmem_n10704, MEM_stage_inst_dmem_n10705, MEM_stage_inst_dmem_n10706, MEM_stage_inst_dmem_n10707, MEM_stage_inst_dmem_n10708, MEM_stage_inst_dmem_n10709, MEM_stage_inst_dmem_n10710, MEM_stage_inst_dmem_n10711, MEM_stage_inst_dmem_n10712, MEM_stage_inst_dmem_n10713, MEM_stage_inst_dmem_n10714, MEM_stage_inst_dmem_n10715, MEM_stage_inst_dmem_n10716, MEM_stage_inst_dmem_n10717, MEM_stage_inst_dmem_n10718, MEM_stage_inst_dmem_n10719, MEM_stage_inst_dmem_n10720, MEM_stage_inst_dmem_n10721, MEM_stage_inst_dmem_n10722, MEM_stage_inst_dmem_n10723, MEM_stage_inst_dmem_n10724, MEM_stage_inst_dmem_n10725, MEM_stage_inst_dmem_n10726, MEM_stage_inst_dmem_n10727, MEM_stage_inst_dmem_n10728, MEM_stage_inst_dmem_n10729, MEM_stage_inst_dmem_n10730, MEM_stage_inst_dmem_n10731, MEM_stage_inst_dmem_n10732, MEM_stage_inst_dmem_n10733, MEM_stage_inst_dmem_n10734, MEM_stage_inst_dmem_n10735, MEM_stage_inst_dmem_n10736, MEM_stage_inst_dmem_n10737, MEM_stage_inst_dmem_n10738, MEM_stage_inst_dmem_n10739, MEM_stage_inst_dmem_n10740, MEM_stage_inst_dmem_n10741, MEM_stage_inst_dmem_n10742, MEM_stage_inst_dmem_n10743, MEM_stage_inst_dmem_n10744, MEM_stage_inst_dmem_n10745, MEM_stage_inst_dmem_n10746, MEM_stage_inst_dmem_n10747, MEM_stage_inst_dmem_n10748, MEM_stage_inst_dmem_n10749, MEM_stage_inst_dmem_n10750, MEM_stage_inst_dmem_n10751, MEM_stage_inst_dmem_n10752, MEM_stage_inst_dmem_n10753, MEM_stage_inst_dmem_n10754, MEM_stage_inst_dmem_n10755, MEM_stage_inst_dmem_n10756, MEM_stage_inst_dmem_n10757, MEM_stage_inst_dmem_n10758, MEM_stage_inst_dmem_n10759, MEM_stage_inst_dmem_n10760, MEM_stage_inst_dmem_n10761, MEM_stage_inst_dmem_n10762, MEM_stage_inst_dmem_n10763, MEM_stage_inst_dmem_n10764, MEM_stage_inst_dmem_n10765, MEM_stage_inst_dmem_n10766, MEM_stage_inst_dmem_n10767, MEM_stage_inst_dmem_n10768, MEM_stage_inst_dmem_n10769, MEM_stage_inst_dmem_n10770, MEM_stage_inst_dmem_n10771, MEM_stage_inst_dmem_n10772, MEM_stage_inst_dmem_n10773, MEM_stage_inst_dmem_n10774, MEM_stage_inst_dmem_n10775, MEM_stage_inst_dmem_n10776, MEM_stage_inst_dmem_n10777, MEM_stage_inst_dmem_n10778, MEM_stage_inst_dmem_n10779, MEM_stage_inst_dmem_n10780, MEM_stage_inst_dmem_n10781, MEM_stage_inst_dmem_n10782, MEM_stage_inst_dmem_n10783, MEM_stage_inst_dmem_n10784, MEM_stage_inst_dmem_n10785, MEM_stage_inst_dmem_n10786, MEM_stage_inst_dmem_n10787, MEM_stage_inst_dmem_n10788, MEM_stage_inst_dmem_n10789, MEM_stage_inst_dmem_n10790, MEM_stage_inst_dmem_n10791, MEM_stage_inst_dmem_n10792, MEM_stage_inst_dmem_n10793, MEM_stage_inst_dmem_n10794, MEM_stage_inst_dmem_n10795, MEM_stage_inst_dmem_n10796, MEM_stage_inst_dmem_n10797, MEM_stage_inst_dmem_n10798, MEM_stage_inst_dmem_n10799, MEM_stage_inst_dmem_n10800, MEM_stage_inst_dmem_n10801, MEM_stage_inst_dmem_n10802, MEM_stage_inst_dmem_n10803, MEM_stage_inst_dmem_n10804, MEM_stage_inst_dmem_n10805, MEM_stage_inst_dmem_n10806, MEM_stage_inst_dmem_n10807, MEM_stage_inst_dmem_n10808, MEM_stage_inst_dmem_n10809, MEM_stage_inst_dmem_n10810, MEM_stage_inst_dmem_n10811, MEM_stage_inst_dmem_n10812, MEM_stage_inst_dmem_n10813, MEM_stage_inst_dmem_n10814, MEM_stage_inst_dmem_n10815, MEM_stage_inst_dmem_n10816, MEM_stage_inst_dmem_n10817, MEM_stage_inst_dmem_n10818, MEM_stage_inst_dmem_n10819, MEM_stage_inst_dmem_n10820, MEM_stage_inst_dmem_n10821, MEM_stage_inst_dmem_n10822, MEM_stage_inst_dmem_n10823, MEM_stage_inst_dmem_n10824, MEM_stage_inst_dmem_n10825, MEM_stage_inst_dmem_n10826, MEM_stage_inst_dmem_n10827, MEM_stage_inst_dmem_n10828, MEM_stage_inst_dmem_n10829, MEM_stage_inst_dmem_n10830, MEM_stage_inst_dmem_n10831, MEM_stage_inst_dmem_n10832, MEM_stage_inst_dmem_n10833, MEM_stage_inst_dmem_n10834, MEM_stage_inst_dmem_n10835, MEM_stage_inst_dmem_n10836, MEM_stage_inst_dmem_n10837, MEM_stage_inst_dmem_n10838, MEM_stage_inst_dmem_n10839, MEM_stage_inst_dmem_n10840, MEM_stage_inst_dmem_n10841, MEM_stage_inst_dmem_n10842, MEM_stage_inst_dmem_n10843, MEM_stage_inst_dmem_n10844, MEM_stage_inst_dmem_n10845, MEM_stage_inst_dmem_n10846, MEM_stage_inst_dmem_n10847, MEM_stage_inst_dmem_n10848, MEM_stage_inst_dmem_n10849, MEM_stage_inst_dmem_n10850, MEM_stage_inst_dmem_n10851, MEM_stage_inst_dmem_n10852, MEM_stage_inst_dmem_n10853, MEM_stage_inst_dmem_n10854, MEM_stage_inst_dmem_n10855, MEM_stage_inst_dmem_n10856, MEM_stage_inst_dmem_n10857, MEM_stage_inst_dmem_n10858, MEM_stage_inst_dmem_n10859, MEM_stage_inst_dmem_n10860, MEM_stage_inst_dmem_n10861, MEM_stage_inst_dmem_n10862, MEM_stage_inst_dmem_n10863, MEM_stage_inst_dmem_n10864, MEM_stage_inst_dmem_n10865, MEM_stage_inst_dmem_n10866, MEM_stage_inst_dmem_n10867, MEM_stage_inst_dmem_n10868, MEM_stage_inst_dmem_n10869, MEM_stage_inst_dmem_n10870, MEM_stage_inst_dmem_n10871, MEM_stage_inst_dmem_n10872, MEM_stage_inst_dmem_n10873, MEM_stage_inst_dmem_n10874, MEM_stage_inst_dmem_n10875, MEM_stage_inst_dmem_n10876, MEM_stage_inst_dmem_n10877, MEM_stage_inst_dmem_n10878, MEM_stage_inst_dmem_n10879, MEM_stage_inst_dmem_n10880, MEM_stage_inst_dmem_n10881, MEM_stage_inst_dmem_n10882, MEM_stage_inst_dmem_n10883, MEM_stage_inst_dmem_n10884, MEM_stage_inst_dmem_n10885, MEM_stage_inst_dmem_n10886, MEM_stage_inst_dmem_n10887, MEM_stage_inst_dmem_n10888, MEM_stage_inst_dmem_n10889, MEM_stage_inst_dmem_n10890, MEM_stage_inst_dmem_n10891, MEM_stage_inst_dmem_n10892, MEM_stage_inst_dmem_n10893, MEM_stage_inst_dmem_n10894, MEM_stage_inst_dmem_n10895, MEM_stage_inst_dmem_n10896, MEM_stage_inst_dmem_n10897, MEM_stage_inst_dmem_n10898, MEM_stage_inst_dmem_n10899, MEM_stage_inst_dmem_n10900, MEM_stage_inst_dmem_n10901, MEM_stage_inst_dmem_n10902, MEM_stage_inst_dmem_n10903, MEM_stage_inst_dmem_n10904, MEM_stage_inst_dmem_n10905, MEM_stage_inst_dmem_n10906, MEM_stage_inst_dmem_n10907, MEM_stage_inst_dmem_n10908, MEM_stage_inst_dmem_n10909, MEM_stage_inst_dmem_n10910, MEM_stage_inst_dmem_n10911, MEM_stage_inst_dmem_n10912, MEM_stage_inst_dmem_n10913, MEM_stage_inst_dmem_n10914, MEM_stage_inst_dmem_n10915, MEM_stage_inst_dmem_n10916, MEM_stage_inst_dmem_n10917, MEM_stage_inst_dmem_n10918, MEM_stage_inst_dmem_n10919, MEM_stage_inst_dmem_n10920, MEM_stage_inst_dmem_n10921, MEM_stage_inst_dmem_n10922, MEM_stage_inst_dmem_n10923, MEM_stage_inst_dmem_n10924, MEM_stage_inst_dmem_n10925, MEM_stage_inst_dmem_n10926, MEM_stage_inst_dmem_n10927, MEM_stage_inst_dmem_n10928, MEM_stage_inst_dmem_n10929, MEM_stage_inst_dmem_n10930, MEM_stage_inst_dmem_n10931, MEM_stage_inst_dmem_n10932, MEM_stage_inst_dmem_n10933, MEM_stage_inst_dmem_n10934, MEM_stage_inst_dmem_n10935, MEM_stage_inst_dmem_n10936, MEM_stage_inst_dmem_n10937, MEM_stage_inst_dmem_n10938, MEM_stage_inst_dmem_n10939, MEM_stage_inst_dmem_n10940, MEM_stage_inst_dmem_n10941, MEM_stage_inst_dmem_n10942, MEM_stage_inst_dmem_n10943, MEM_stage_inst_dmem_n10944, MEM_stage_inst_dmem_n10945, MEM_stage_inst_dmem_n10946, MEM_stage_inst_dmem_n10947, MEM_stage_inst_dmem_n10948, MEM_stage_inst_dmem_n10949, MEM_stage_inst_dmem_n10950, MEM_stage_inst_dmem_n10951, MEM_stage_inst_dmem_n10952, MEM_stage_inst_dmem_n10953, MEM_stage_inst_dmem_n10954, MEM_stage_inst_dmem_n10955, MEM_stage_inst_dmem_n10956, MEM_stage_inst_dmem_n10957, MEM_stage_inst_dmem_n10958, MEM_stage_inst_dmem_n10959, MEM_stage_inst_dmem_n10960, MEM_stage_inst_dmem_n10961, MEM_stage_inst_dmem_n10962, MEM_stage_inst_dmem_n10963, MEM_stage_inst_dmem_n10964, MEM_stage_inst_dmem_n10965, MEM_stage_inst_dmem_n10966, MEM_stage_inst_dmem_n10967, MEM_stage_inst_dmem_n10968, MEM_stage_inst_dmem_n10969, MEM_stage_inst_dmem_n10970, MEM_stage_inst_dmem_n10971, MEM_stage_inst_dmem_n10972, MEM_stage_inst_dmem_n10973, MEM_stage_inst_dmem_n10974, MEM_stage_inst_dmem_n10975, MEM_stage_inst_dmem_n10976, MEM_stage_inst_dmem_n10977, MEM_stage_inst_dmem_n10978, MEM_stage_inst_dmem_n10979, MEM_stage_inst_dmem_n10980, MEM_stage_inst_dmem_n10981, MEM_stage_inst_dmem_n10982, MEM_stage_inst_dmem_n10983, MEM_stage_inst_dmem_n10984, MEM_stage_inst_dmem_n10985, MEM_stage_inst_dmem_n10986, MEM_stage_inst_dmem_n10987, MEM_stage_inst_dmem_n10988, MEM_stage_inst_dmem_n10989, MEM_stage_inst_dmem_n10990, MEM_stage_inst_dmem_n10991, MEM_stage_inst_dmem_n10992, MEM_stage_inst_dmem_n10993, MEM_stage_inst_dmem_n10994, MEM_stage_inst_dmem_n10995, MEM_stage_inst_dmem_n10996, MEM_stage_inst_dmem_n10997, MEM_stage_inst_dmem_n10998, MEM_stage_inst_dmem_n10999, MEM_stage_inst_dmem_n11000, MEM_stage_inst_dmem_n11001, MEM_stage_inst_dmem_n11002, MEM_stage_inst_dmem_n11003, MEM_stage_inst_dmem_n11004, MEM_stage_inst_dmem_n11005, MEM_stage_inst_dmem_n11006, MEM_stage_inst_dmem_n11007, MEM_stage_inst_dmem_n11008, MEM_stage_inst_dmem_n11009, MEM_stage_inst_dmem_n11010, MEM_stage_inst_dmem_n11011, MEM_stage_inst_dmem_n11012, MEM_stage_inst_dmem_n11013, MEM_stage_inst_dmem_n11014, MEM_stage_inst_dmem_n11015, MEM_stage_inst_dmem_n11016, MEM_stage_inst_dmem_n11017, MEM_stage_inst_dmem_n11018, MEM_stage_inst_dmem_n11019, MEM_stage_inst_dmem_n11020, MEM_stage_inst_dmem_n11021, MEM_stage_inst_dmem_n11022, MEM_stage_inst_dmem_n11023, MEM_stage_inst_dmem_n11024, MEM_stage_inst_dmem_n11025, MEM_stage_inst_dmem_n11026, MEM_stage_inst_dmem_n11027, MEM_stage_inst_dmem_n11028, MEM_stage_inst_dmem_n11029, MEM_stage_inst_dmem_n11030, MEM_stage_inst_dmem_n11031, MEM_stage_inst_dmem_n11032, MEM_stage_inst_dmem_n11033, MEM_stage_inst_dmem_n11034, MEM_stage_inst_dmem_n11035, MEM_stage_inst_dmem_n11036, MEM_stage_inst_dmem_n11037, MEM_stage_inst_dmem_n11038, MEM_stage_inst_dmem_n11039, MEM_stage_inst_dmem_n11040, MEM_stage_inst_dmem_n11041, MEM_stage_inst_dmem_n11042, MEM_stage_inst_dmem_n11043, MEM_stage_inst_dmem_n11044, MEM_stage_inst_dmem_n11045, MEM_stage_inst_dmem_n11046, MEM_stage_inst_dmem_n11047, MEM_stage_inst_dmem_n11048, MEM_stage_inst_dmem_n11049, MEM_stage_inst_dmem_n11050, MEM_stage_inst_dmem_n11051, MEM_stage_inst_dmem_n11052, MEM_stage_inst_dmem_n11053, MEM_stage_inst_dmem_n11054, MEM_stage_inst_dmem_n11055, MEM_stage_inst_dmem_n11056, MEM_stage_inst_dmem_n11057, MEM_stage_inst_dmem_n11058, MEM_stage_inst_dmem_n11059, MEM_stage_inst_dmem_n11060, MEM_stage_inst_dmem_n11061, MEM_stage_inst_dmem_n11062, MEM_stage_inst_dmem_n11063, MEM_stage_inst_dmem_n11064, MEM_stage_inst_dmem_n11065, MEM_stage_inst_dmem_n11066, MEM_stage_inst_dmem_n11067, MEM_stage_inst_dmem_n11068, MEM_stage_inst_dmem_n11069, MEM_stage_inst_dmem_n11070, MEM_stage_inst_dmem_n11071, MEM_stage_inst_dmem_n11072, MEM_stage_inst_dmem_n11073, MEM_stage_inst_dmem_n11074, MEM_stage_inst_dmem_n11075, MEM_stage_inst_dmem_n11076, MEM_stage_inst_dmem_n11077, MEM_stage_inst_dmem_n11078, MEM_stage_inst_dmem_n11079, MEM_stage_inst_dmem_n11080, MEM_stage_inst_dmem_n11081, MEM_stage_inst_dmem_n11082, MEM_stage_inst_dmem_n11083, MEM_stage_inst_dmem_n11084, MEM_stage_inst_dmem_n11085, MEM_stage_inst_dmem_n11086, MEM_stage_inst_dmem_n11087, MEM_stage_inst_dmem_n11088, MEM_stage_inst_dmem_n11089, MEM_stage_inst_dmem_n11090, MEM_stage_inst_dmem_n11091, MEM_stage_inst_dmem_n11092, MEM_stage_inst_dmem_n11093, MEM_stage_inst_dmem_n11094, MEM_stage_inst_dmem_n11095, MEM_stage_inst_dmem_n11096, MEM_stage_inst_dmem_n11097, MEM_stage_inst_dmem_n11098, MEM_stage_inst_dmem_n11099, MEM_stage_inst_dmem_n11100, MEM_stage_inst_dmem_n11101, MEM_stage_inst_dmem_n11102, MEM_stage_inst_dmem_n11103, MEM_stage_inst_dmem_n11104, MEM_stage_inst_dmem_n11105, MEM_stage_inst_dmem_n11106, MEM_stage_inst_dmem_n11107, MEM_stage_inst_dmem_n11108, MEM_stage_inst_dmem_n11109, MEM_stage_inst_dmem_n11110, MEM_stage_inst_dmem_n11111, MEM_stage_inst_dmem_n11112, MEM_stage_inst_dmem_n11113, MEM_stage_inst_dmem_n11114, MEM_stage_inst_dmem_n11115, MEM_stage_inst_dmem_n11116, MEM_stage_inst_dmem_n11117, MEM_stage_inst_dmem_n11118, MEM_stage_inst_dmem_n11119, MEM_stage_inst_dmem_n11120, MEM_stage_inst_dmem_n11121, MEM_stage_inst_dmem_n11122, MEM_stage_inst_dmem_n11123, MEM_stage_inst_dmem_n11124, MEM_stage_inst_dmem_n11125, MEM_stage_inst_dmem_n11126, MEM_stage_inst_dmem_n11127, MEM_stage_inst_dmem_n11128, MEM_stage_inst_dmem_n11129, MEM_stage_inst_dmem_n11130, MEM_stage_inst_dmem_n11131, MEM_stage_inst_dmem_n11132, MEM_stage_inst_dmem_n11133, MEM_stage_inst_dmem_n11134, MEM_stage_inst_dmem_n11135, MEM_stage_inst_dmem_n11136, MEM_stage_inst_dmem_n11137, MEM_stage_inst_dmem_n11138, MEM_stage_inst_dmem_n11139, MEM_stage_inst_dmem_n11140, MEM_stage_inst_dmem_n11141, MEM_stage_inst_dmem_n11142, MEM_stage_inst_dmem_n11143, MEM_stage_inst_dmem_n11144, MEM_stage_inst_dmem_n11145, MEM_stage_inst_dmem_n11146, MEM_stage_inst_dmem_n11147, MEM_stage_inst_dmem_n11148, MEM_stage_inst_dmem_n11149, MEM_stage_inst_dmem_n11150, MEM_stage_inst_dmem_n11151, MEM_stage_inst_dmem_n11152, MEM_stage_inst_dmem_n11153, MEM_stage_inst_dmem_n11154, MEM_stage_inst_dmem_n11155, MEM_stage_inst_dmem_n11156, MEM_stage_inst_dmem_n11157, MEM_stage_inst_dmem_n11158, MEM_stage_inst_dmem_n11159, MEM_stage_inst_dmem_n11160, MEM_stage_inst_dmem_n11161, MEM_stage_inst_dmem_n11162, MEM_stage_inst_dmem_n11163, MEM_stage_inst_dmem_n11164, MEM_stage_inst_dmem_n11165, MEM_stage_inst_dmem_n11166, MEM_stage_inst_dmem_n11167, MEM_stage_inst_dmem_n11168, MEM_stage_inst_dmem_n11169, MEM_stage_inst_dmem_n11170, MEM_stage_inst_dmem_n11171, MEM_stage_inst_dmem_n11172, MEM_stage_inst_dmem_n11173, MEM_stage_inst_dmem_n11174, MEM_stage_inst_dmem_n11175, MEM_stage_inst_dmem_n11176, MEM_stage_inst_dmem_n11177, MEM_stage_inst_dmem_n11178, MEM_stage_inst_dmem_n11179, MEM_stage_inst_dmem_n11180, MEM_stage_inst_dmem_n11181, MEM_stage_inst_dmem_n11182, MEM_stage_inst_dmem_n11183, MEM_stage_inst_dmem_n11184, MEM_stage_inst_dmem_n11185, MEM_stage_inst_dmem_n11186, MEM_stage_inst_dmem_n11187, MEM_stage_inst_dmem_n11188, MEM_stage_inst_dmem_n11189, MEM_stage_inst_dmem_n11190, MEM_stage_inst_dmem_n11191, MEM_stage_inst_dmem_n11192, MEM_stage_inst_dmem_n11193, MEM_stage_inst_dmem_n11194, MEM_stage_inst_dmem_n11195, MEM_stage_inst_dmem_n11196, MEM_stage_inst_dmem_n11197, MEM_stage_inst_dmem_n11198, MEM_stage_inst_dmem_n11199, MEM_stage_inst_dmem_n11200, MEM_stage_inst_dmem_n11201, MEM_stage_inst_dmem_n11202, MEM_stage_inst_dmem_n11203, MEM_stage_inst_dmem_n11204, MEM_stage_inst_dmem_n11205, MEM_stage_inst_dmem_n11206, MEM_stage_inst_dmem_n11207, MEM_stage_inst_dmem_n11208, MEM_stage_inst_dmem_n11209, MEM_stage_inst_dmem_n11210, MEM_stage_inst_dmem_n11211, MEM_stage_inst_dmem_n11212, MEM_stage_inst_dmem_n11213, MEM_stage_inst_dmem_n11214, MEM_stage_inst_dmem_n11215, MEM_stage_inst_dmem_n11216, MEM_stage_inst_dmem_n11217, MEM_stage_inst_dmem_n11218, MEM_stage_inst_dmem_n11219, MEM_stage_inst_dmem_n11220, MEM_stage_inst_dmem_n11221, MEM_stage_inst_dmem_n11222, MEM_stage_inst_dmem_n11223, MEM_stage_inst_dmem_n11224, MEM_stage_inst_dmem_n11225, MEM_stage_inst_dmem_n11226, MEM_stage_inst_dmem_n11227, MEM_stage_inst_dmem_n11228, MEM_stage_inst_dmem_n11229, MEM_stage_inst_dmem_n11230, MEM_stage_inst_dmem_n11231, MEM_stage_inst_dmem_n11232, MEM_stage_inst_dmem_n11233, MEM_stage_inst_dmem_n11234, MEM_stage_inst_dmem_n11235, MEM_stage_inst_dmem_n11236, MEM_stage_inst_dmem_n11237, MEM_stage_inst_dmem_n11238, MEM_stage_inst_dmem_n11239, MEM_stage_inst_dmem_n11240, MEM_stage_inst_dmem_n11241, MEM_stage_inst_dmem_n11242, MEM_stage_inst_dmem_n11243, MEM_stage_inst_dmem_n11244, MEM_stage_inst_dmem_n11245, MEM_stage_inst_dmem_n11246, MEM_stage_inst_dmem_n11247, MEM_stage_inst_dmem_n11248, MEM_stage_inst_dmem_n11249, MEM_stage_inst_dmem_n11250, MEM_stage_inst_dmem_n11251, MEM_stage_inst_dmem_n11252, MEM_stage_inst_dmem_n11253, MEM_stage_inst_dmem_n11254, MEM_stage_inst_dmem_n11255, MEM_stage_inst_dmem_n11256, MEM_stage_inst_dmem_n11257, MEM_stage_inst_dmem_n11258, MEM_stage_inst_dmem_n11259, MEM_stage_inst_dmem_n11260, MEM_stage_inst_dmem_n11261, MEM_stage_inst_dmem_n11262, MEM_stage_inst_dmem_n11263, MEM_stage_inst_dmem_n11264, MEM_stage_inst_dmem_n11265, MEM_stage_inst_dmem_n11266, MEM_stage_inst_dmem_n11267, MEM_stage_inst_dmem_n11268, MEM_stage_inst_dmem_n11269, MEM_stage_inst_dmem_n11270, MEM_stage_inst_dmem_n11271, MEM_stage_inst_dmem_n11272, MEM_stage_inst_dmem_n11273, MEM_stage_inst_dmem_n11274, MEM_stage_inst_dmem_n11275, MEM_stage_inst_dmem_n11276, MEM_stage_inst_dmem_n11277, MEM_stage_inst_dmem_n11278, MEM_stage_inst_dmem_n11279, MEM_stage_inst_dmem_n11280, MEM_stage_inst_dmem_n11281, MEM_stage_inst_dmem_n11282, MEM_stage_inst_dmem_n11283, MEM_stage_inst_dmem_n11284, MEM_stage_inst_dmem_n11285, MEM_stage_inst_dmem_n11286, MEM_stage_inst_dmem_n11287, MEM_stage_inst_dmem_n11288, MEM_stage_inst_dmem_n11289, MEM_stage_inst_dmem_n11290, MEM_stage_inst_dmem_n11291, MEM_stage_inst_dmem_n11292, MEM_stage_inst_dmem_n11293, MEM_stage_inst_dmem_n11294, MEM_stage_inst_dmem_n11295, MEM_stage_inst_dmem_n11296, MEM_stage_inst_dmem_n11297, MEM_stage_inst_dmem_n11298, MEM_stage_inst_dmem_n11299, MEM_stage_inst_dmem_n11300, MEM_stage_inst_dmem_n11301, MEM_stage_inst_dmem_n11302, MEM_stage_inst_dmem_n11303, MEM_stage_inst_dmem_n11304, MEM_stage_inst_dmem_n11305, MEM_stage_inst_dmem_n11306, MEM_stage_inst_dmem_n11307, MEM_stage_inst_dmem_n11308, MEM_stage_inst_dmem_n11309, MEM_stage_inst_dmem_n11310, MEM_stage_inst_dmem_n11311, MEM_stage_inst_dmem_n11312, MEM_stage_inst_dmem_n11313, MEM_stage_inst_dmem_n11314, MEM_stage_inst_dmem_n11315, MEM_stage_inst_dmem_n11316, MEM_stage_inst_dmem_n11317, MEM_stage_inst_dmem_n11318, MEM_stage_inst_dmem_n11319, MEM_stage_inst_dmem_n11320, MEM_stage_inst_dmem_n11321, MEM_stage_inst_dmem_n11322, MEM_stage_inst_dmem_n11323, MEM_stage_inst_dmem_n11324, MEM_stage_inst_dmem_n11325, MEM_stage_inst_dmem_n11326, MEM_stage_inst_dmem_n11327, MEM_stage_inst_dmem_n11328, MEM_stage_inst_dmem_n11329, MEM_stage_inst_dmem_n11330, MEM_stage_inst_dmem_n11331, MEM_stage_inst_dmem_n11332, MEM_stage_inst_dmem_n11333, MEM_stage_inst_dmem_n11334, MEM_stage_inst_dmem_n11335, MEM_stage_inst_dmem_n11336, MEM_stage_inst_dmem_n11337, MEM_stage_inst_dmem_n11338, MEM_stage_inst_dmem_n11339, MEM_stage_inst_dmem_n11340, MEM_stage_inst_dmem_n11341, MEM_stage_inst_dmem_n11342, MEM_stage_inst_dmem_n11343, MEM_stage_inst_dmem_n11344, MEM_stage_inst_dmem_n11345, MEM_stage_inst_dmem_n11346, MEM_stage_inst_dmem_n11347, MEM_stage_inst_dmem_n11348, MEM_stage_inst_dmem_n11349, MEM_stage_inst_dmem_n11350, MEM_stage_inst_dmem_n11351, MEM_stage_inst_dmem_n11352, MEM_stage_inst_dmem_n11353, MEM_stage_inst_dmem_n11354, MEM_stage_inst_dmem_n11355, MEM_stage_inst_dmem_n11356, MEM_stage_inst_dmem_n11357, MEM_stage_inst_dmem_n11358, MEM_stage_inst_dmem_n11359, MEM_stage_inst_dmem_n11360, MEM_stage_inst_dmem_n11361, MEM_stage_inst_dmem_n11362, MEM_stage_inst_dmem_n11363, MEM_stage_inst_dmem_n11364, MEM_stage_inst_dmem_n11365, MEM_stage_inst_dmem_n11366, MEM_stage_inst_dmem_n11367, MEM_stage_inst_dmem_n11368, MEM_stage_inst_dmem_n11369, MEM_stage_inst_dmem_n11370, MEM_stage_inst_dmem_n11371, MEM_stage_inst_dmem_n11372, MEM_stage_inst_dmem_n11373, MEM_stage_inst_dmem_n11374, MEM_stage_inst_dmem_n11375, MEM_stage_inst_dmem_n11376, MEM_stage_inst_dmem_n11377, MEM_stage_inst_dmem_n11378, MEM_stage_inst_dmem_n11379, MEM_stage_inst_dmem_n11380, MEM_stage_inst_dmem_n11381, MEM_stage_inst_dmem_n11382, MEM_stage_inst_dmem_n11383, MEM_stage_inst_dmem_n11384, MEM_stage_inst_dmem_n11385, MEM_stage_inst_dmem_n11386, MEM_stage_inst_dmem_n11387, MEM_stage_inst_dmem_n11388, MEM_stage_inst_dmem_n11389, MEM_stage_inst_dmem_n11390, MEM_stage_inst_dmem_n11391, MEM_stage_inst_dmem_n11392, MEM_stage_inst_dmem_n11393, MEM_stage_inst_dmem_n11394, MEM_stage_inst_dmem_n11395, MEM_stage_inst_dmem_n11396, MEM_stage_inst_dmem_n11397, MEM_stage_inst_dmem_n11398, MEM_stage_inst_dmem_n11399, MEM_stage_inst_dmem_n11400, MEM_stage_inst_dmem_n11401, MEM_stage_inst_dmem_n11402, MEM_stage_inst_dmem_n11403, MEM_stage_inst_dmem_n11404, MEM_stage_inst_dmem_n11405, MEM_stage_inst_dmem_n11406, MEM_stage_inst_dmem_n11407, MEM_stage_inst_dmem_n11408, MEM_stage_inst_dmem_n11409, MEM_stage_inst_dmem_n11410, MEM_stage_inst_dmem_n11411, MEM_stage_inst_dmem_n11412, MEM_stage_inst_dmem_n11413, MEM_stage_inst_dmem_n11414, MEM_stage_inst_dmem_n11415, MEM_stage_inst_dmem_n11416, MEM_stage_inst_dmem_n11417, MEM_stage_inst_dmem_n11418, MEM_stage_inst_dmem_n11419, MEM_stage_inst_dmem_n11420, MEM_stage_inst_dmem_n11421, MEM_stage_inst_dmem_n11422, MEM_stage_inst_dmem_n11423, MEM_stage_inst_dmem_n11424, MEM_stage_inst_dmem_n11425, MEM_stage_inst_dmem_n11426, MEM_stage_inst_dmem_n11427, MEM_stage_inst_dmem_n11428, MEM_stage_inst_dmem_n11429, MEM_stage_inst_dmem_n11430, MEM_stage_inst_dmem_n11431, MEM_stage_inst_dmem_n11432, MEM_stage_inst_dmem_n11433, MEM_stage_inst_dmem_n11434, MEM_stage_inst_dmem_n11435, MEM_stage_inst_dmem_n11436, MEM_stage_inst_dmem_n11437, MEM_stage_inst_dmem_n11438, MEM_stage_inst_dmem_n11439, MEM_stage_inst_dmem_n11440, MEM_stage_inst_dmem_n11441, MEM_stage_inst_dmem_n11442, MEM_stage_inst_dmem_n11443, MEM_stage_inst_dmem_n11444, MEM_stage_inst_dmem_n11445, MEM_stage_inst_dmem_n11446, MEM_stage_inst_dmem_n11447, MEM_stage_inst_dmem_n11448, MEM_stage_inst_dmem_n11449, MEM_stage_inst_dmem_n11450, MEM_stage_inst_dmem_n11451, MEM_stage_inst_dmem_n11452, MEM_stage_inst_dmem_n11453, MEM_stage_inst_dmem_n11454, MEM_stage_inst_dmem_n11455, MEM_stage_inst_dmem_n11456, MEM_stage_inst_dmem_n11457, MEM_stage_inst_dmem_n11458, MEM_stage_inst_dmem_n11459, MEM_stage_inst_dmem_n11460, MEM_stage_inst_dmem_n11461, MEM_stage_inst_dmem_n11462, MEM_stage_inst_dmem_n11463, MEM_stage_inst_dmem_n11464, MEM_stage_inst_dmem_n11465, MEM_stage_inst_dmem_n11466, MEM_stage_inst_dmem_n11467, MEM_stage_inst_dmem_n11468, MEM_stage_inst_dmem_n11469, MEM_stage_inst_dmem_n11470, MEM_stage_inst_dmem_n11471, MEM_stage_inst_dmem_n11472, MEM_stage_inst_dmem_n11473, MEM_stage_inst_dmem_n11474, MEM_stage_inst_dmem_n11475, MEM_stage_inst_dmem_n11476, MEM_stage_inst_dmem_n11477, MEM_stage_inst_dmem_n11478, MEM_stage_inst_dmem_n11479, MEM_stage_inst_dmem_n11480, MEM_stage_inst_dmem_n11481, MEM_stage_inst_dmem_n11482, MEM_stage_inst_dmem_n11483, MEM_stage_inst_dmem_n11484, MEM_stage_inst_dmem_n11485, MEM_stage_inst_dmem_n11486, MEM_stage_inst_dmem_n11487, MEM_stage_inst_dmem_n11488, MEM_stage_inst_dmem_n11489, MEM_stage_inst_dmem_n11490, MEM_stage_inst_dmem_n11491, MEM_stage_inst_dmem_n11492, MEM_stage_inst_dmem_n11493, MEM_stage_inst_dmem_n11494, MEM_stage_inst_dmem_n11495, MEM_stage_inst_dmem_n11496, MEM_stage_inst_dmem_n11497, MEM_stage_inst_dmem_n11498, MEM_stage_inst_dmem_n11499, MEM_stage_inst_dmem_n11500, MEM_stage_inst_dmem_n11501, MEM_stage_inst_dmem_n11502, MEM_stage_inst_dmem_n11503, MEM_stage_inst_dmem_n11504, MEM_stage_inst_dmem_n11505, MEM_stage_inst_dmem_n11506, MEM_stage_inst_dmem_n11507, MEM_stage_inst_dmem_n11508, MEM_stage_inst_dmem_n11509, MEM_stage_inst_dmem_n11510, MEM_stage_inst_dmem_n11511, MEM_stage_inst_dmem_n11512, MEM_stage_inst_dmem_n11513, MEM_stage_inst_dmem_n11514, MEM_stage_inst_dmem_n11515, MEM_stage_inst_dmem_n11516, MEM_stage_inst_dmem_n11517, MEM_stage_inst_dmem_n11518, MEM_stage_inst_dmem_n11519, MEM_stage_inst_dmem_n11520, MEM_stage_inst_dmem_n11521, MEM_stage_inst_dmem_n11522, MEM_stage_inst_dmem_n11523, MEM_stage_inst_dmem_n11524, MEM_stage_inst_dmem_n11525, MEM_stage_inst_dmem_n11526, MEM_stage_inst_dmem_n11527, MEM_stage_inst_dmem_n11528, MEM_stage_inst_dmem_n11529, MEM_stage_inst_dmem_n11530, MEM_stage_inst_dmem_n11531, MEM_stage_inst_dmem_n11532, MEM_stage_inst_dmem_n11533, MEM_stage_inst_dmem_n11534, MEM_stage_inst_dmem_n11535, MEM_stage_inst_dmem_n11536, MEM_stage_inst_dmem_n11537, MEM_stage_inst_dmem_n11538, MEM_stage_inst_dmem_n11539, MEM_stage_inst_dmem_n11540, MEM_stage_inst_dmem_n11541, MEM_stage_inst_dmem_n11542, MEM_stage_inst_dmem_n11543, MEM_stage_inst_dmem_n11544, MEM_stage_inst_dmem_n11545, MEM_stage_inst_dmem_n11546, MEM_stage_inst_dmem_n11547, MEM_stage_inst_dmem_n11548, MEM_stage_inst_dmem_n11549, MEM_stage_inst_dmem_n11550, MEM_stage_inst_dmem_n11551, MEM_stage_inst_dmem_n11552, MEM_stage_inst_dmem_n11553, MEM_stage_inst_dmem_n11554, MEM_stage_inst_dmem_n11555, MEM_stage_inst_dmem_n11556, MEM_stage_inst_dmem_n11557, MEM_stage_inst_dmem_n11558, MEM_stage_inst_dmem_n11559, MEM_stage_inst_dmem_n11560, MEM_stage_inst_dmem_n11561, MEM_stage_inst_dmem_n11562, MEM_stage_inst_dmem_n11563, MEM_stage_inst_dmem_n11564, MEM_stage_inst_dmem_n11565, MEM_stage_inst_dmem_n11566, MEM_stage_inst_dmem_n11567, MEM_stage_inst_dmem_n11568, MEM_stage_inst_dmem_n11569, MEM_stage_inst_dmem_n11570, MEM_stage_inst_dmem_n11571, MEM_stage_inst_dmem_n11572, MEM_stage_inst_dmem_n11573, MEM_stage_inst_dmem_n11574, MEM_stage_inst_dmem_n11575, MEM_stage_inst_dmem_n11576, MEM_stage_inst_dmem_n11577, MEM_stage_inst_dmem_n11578, MEM_stage_inst_dmem_n11579, MEM_stage_inst_dmem_n11580, MEM_stage_inst_dmem_n11581, MEM_stage_inst_dmem_n11582, MEM_stage_inst_dmem_n11583, MEM_stage_inst_dmem_n11584, MEM_stage_inst_dmem_n11585, MEM_stage_inst_dmem_n11586, MEM_stage_inst_dmem_n11587, MEM_stage_inst_dmem_n11588, MEM_stage_inst_dmem_n11589, MEM_stage_inst_dmem_n11590, MEM_stage_inst_dmem_n11591, MEM_stage_inst_dmem_n11592, MEM_stage_inst_dmem_n11593, MEM_stage_inst_dmem_n11594, MEM_stage_inst_dmem_n11595, MEM_stage_inst_dmem_n11596, MEM_stage_inst_dmem_n11597, MEM_stage_inst_dmem_n11598, MEM_stage_inst_dmem_n11599, MEM_stage_inst_dmem_n11600, MEM_stage_inst_dmem_n11601, MEM_stage_inst_dmem_n11602, MEM_stage_inst_dmem_n11603, MEM_stage_inst_dmem_n11604, MEM_stage_inst_dmem_n11605, MEM_stage_inst_dmem_n11606, MEM_stage_inst_dmem_n11607, MEM_stage_inst_dmem_n11608, MEM_stage_inst_dmem_n11609, MEM_stage_inst_dmem_n11610, MEM_stage_inst_dmem_n11611, MEM_stage_inst_dmem_n11612, MEM_stage_inst_dmem_n11613, MEM_stage_inst_dmem_n11614, MEM_stage_inst_dmem_n11615, MEM_stage_inst_dmem_n11616, MEM_stage_inst_dmem_n11617, MEM_stage_inst_dmem_n11618, MEM_stage_inst_dmem_n11619, MEM_stage_inst_dmem_n11620, MEM_stage_inst_dmem_n11621, MEM_stage_inst_dmem_n11622, MEM_stage_inst_dmem_n11623, MEM_stage_inst_dmem_n11624, MEM_stage_inst_dmem_n11625, MEM_stage_inst_dmem_n11626, MEM_stage_inst_dmem_n11627, MEM_stage_inst_dmem_n11628, MEM_stage_inst_dmem_n11629, MEM_stage_inst_dmem_n11630, MEM_stage_inst_dmem_n11631, MEM_stage_inst_dmem_n11632, MEM_stage_inst_dmem_n11633, MEM_stage_inst_dmem_n11634, MEM_stage_inst_dmem_n11635, MEM_stage_inst_dmem_n11636, MEM_stage_inst_dmem_n11637, MEM_stage_inst_dmem_n11638, MEM_stage_inst_dmem_n11639, MEM_stage_inst_dmem_n11640, MEM_stage_inst_dmem_n11641, MEM_stage_inst_dmem_n11642, MEM_stage_inst_dmem_n11643, MEM_stage_inst_dmem_n11644, MEM_stage_inst_dmem_n11645, MEM_stage_inst_dmem_n11646, MEM_stage_inst_dmem_n11647, MEM_stage_inst_dmem_n11648, MEM_stage_inst_dmem_n11649, MEM_stage_inst_dmem_n11650, MEM_stage_inst_dmem_n11651, MEM_stage_inst_dmem_n11652, MEM_stage_inst_dmem_n11653, MEM_stage_inst_dmem_n11654, MEM_stage_inst_dmem_n11655, MEM_stage_inst_dmem_n11656, MEM_stage_inst_dmem_n11657, MEM_stage_inst_dmem_n11658, MEM_stage_inst_dmem_n11659, MEM_stage_inst_dmem_n11660, MEM_stage_inst_dmem_n11661, MEM_stage_inst_dmem_n11662, MEM_stage_inst_dmem_n11663, MEM_stage_inst_dmem_n11664, MEM_stage_inst_dmem_n11665, MEM_stage_inst_dmem_n11666, MEM_stage_inst_dmem_n11667, MEM_stage_inst_dmem_n11668, MEM_stage_inst_dmem_n11669, MEM_stage_inst_dmem_n11670, MEM_stage_inst_dmem_n11671, MEM_stage_inst_dmem_n11672, MEM_stage_inst_dmem_n11673, MEM_stage_inst_dmem_n11674, MEM_stage_inst_dmem_n11675, MEM_stage_inst_dmem_n11676, MEM_stage_inst_dmem_n11677, MEM_stage_inst_dmem_n11678, MEM_stage_inst_dmem_n11679, MEM_stage_inst_dmem_n11680, MEM_stage_inst_dmem_n11681, MEM_stage_inst_dmem_n11682, MEM_stage_inst_dmem_n11683, MEM_stage_inst_dmem_n11684, MEM_stage_inst_dmem_n11685, MEM_stage_inst_dmem_n11686, MEM_stage_inst_dmem_n11687, MEM_stage_inst_dmem_n11688, MEM_stage_inst_dmem_n11689, MEM_stage_inst_dmem_n11690, MEM_stage_inst_dmem_n11691, MEM_stage_inst_dmem_n11692, MEM_stage_inst_dmem_n11693, MEM_stage_inst_dmem_n11694, MEM_stage_inst_dmem_n11695, MEM_stage_inst_dmem_n11696, MEM_stage_inst_dmem_n11697, MEM_stage_inst_dmem_n11698, MEM_stage_inst_dmem_n11699, MEM_stage_inst_dmem_n11700, MEM_stage_inst_dmem_n11701, MEM_stage_inst_dmem_n11702, MEM_stage_inst_dmem_n11703, MEM_stage_inst_dmem_n11704, MEM_stage_inst_dmem_n11705, MEM_stage_inst_dmem_n11706, MEM_stage_inst_dmem_n11707, MEM_stage_inst_dmem_n11708, MEM_stage_inst_dmem_n11709, MEM_stage_inst_dmem_n11710, MEM_stage_inst_dmem_n11711, MEM_stage_inst_dmem_n11712, MEM_stage_inst_dmem_n11713, MEM_stage_inst_dmem_n11714, MEM_stage_inst_dmem_n11715, MEM_stage_inst_dmem_n11716, MEM_stage_inst_dmem_n11717, MEM_stage_inst_dmem_n11718, MEM_stage_inst_dmem_n11719, MEM_stage_inst_dmem_n11720, MEM_stage_inst_dmem_n11721, MEM_stage_inst_dmem_n11722, MEM_stage_inst_dmem_n11723, MEM_stage_inst_dmem_n11724, MEM_stage_inst_dmem_n11725, MEM_stage_inst_dmem_n11726, MEM_stage_inst_dmem_n11727, MEM_stage_inst_dmem_n11728, MEM_stage_inst_dmem_n11729, MEM_stage_inst_dmem_n11730, MEM_stage_inst_dmem_n11731, MEM_stage_inst_dmem_n11732, MEM_stage_inst_dmem_n11733, MEM_stage_inst_dmem_n11734, MEM_stage_inst_dmem_n11735, MEM_stage_inst_dmem_n11736, MEM_stage_inst_dmem_n11737, MEM_stage_inst_dmem_n11738, MEM_stage_inst_dmem_n11739, MEM_stage_inst_dmem_n11740, MEM_stage_inst_dmem_n11741, MEM_stage_inst_dmem_n11742, MEM_stage_inst_dmem_n11743, MEM_stage_inst_dmem_n11744, MEM_stage_inst_dmem_n11745, MEM_stage_inst_dmem_n11746, MEM_stage_inst_dmem_n11747, MEM_stage_inst_dmem_n11748, MEM_stage_inst_dmem_n11749, MEM_stage_inst_dmem_n11750, MEM_stage_inst_dmem_n11751, MEM_stage_inst_dmem_n11752, MEM_stage_inst_dmem_n11753, MEM_stage_inst_dmem_n11754, MEM_stage_inst_dmem_n11755, MEM_stage_inst_dmem_n11756, MEM_stage_inst_dmem_n11757, MEM_stage_inst_dmem_n11758, MEM_stage_inst_dmem_n11759, MEM_stage_inst_dmem_n11760, MEM_stage_inst_dmem_n11761, MEM_stage_inst_dmem_n11762, MEM_stage_inst_dmem_n11763, MEM_stage_inst_dmem_n11764, MEM_stage_inst_dmem_n11765, MEM_stage_inst_dmem_n11766, MEM_stage_inst_dmem_n11767, MEM_stage_inst_dmem_n11768, MEM_stage_inst_dmem_n11769, MEM_stage_inst_dmem_n11770, MEM_stage_inst_dmem_n11771, MEM_stage_inst_dmem_n11772, MEM_stage_inst_dmem_n11773, MEM_stage_inst_dmem_n11774, MEM_stage_inst_dmem_n11775, MEM_stage_inst_dmem_n11776, MEM_stage_inst_dmem_n11777, MEM_stage_inst_dmem_n11778, MEM_stage_inst_dmem_n11779, MEM_stage_inst_dmem_n11780, MEM_stage_inst_dmem_n11781, MEM_stage_inst_dmem_n11782, MEM_stage_inst_dmem_n11783, MEM_stage_inst_dmem_n11784, MEM_stage_inst_dmem_n11785, MEM_stage_inst_dmem_n11786, MEM_stage_inst_dmem_n11787, MEM_stage_inst_dmem_n11788, MEM_stage_inst_dmem_n11789, MEM_stage_inst_dmem_n11790, MEM_stage_inst_dmem_n11791, MEM_stage_inst_dmem_n11792, MEM_stage_inst_dmem_n11793, MEM_stage_inst_dmem_n11794, MEM_stage_inst_dmem_n11795, MEM_stage_inst_dmem_n11796, MEM_stage_inst_dmem_n11797, MEM_stage_inst_dmem_n11798, MEM_stage_inst_dmem_n11799, MEM_stage_inst_dmem_n11800, MEM_stage_inst_dmem_n11801, MEM_stage_inst_dmem_n11802, MEM_stage_inst_dmem_n11803, MEM_stage_inst_dmem_n11804, MEM_stage_inst_dmem_n11805, MEM_stage_inst_dmem_n11806, MEM_stage_inst_dmem_n11807, MEM_stage_inst_dmem_n11808, MEM_stage_inst_dmem_n11809, MEM_stage_inst_dmem_n11810, MEM_stage_inst_dmem_n11811, MEM_stage_inst_dmem_n11812, MEM_stage_inst_dmem_n11813, MEM_stage_inst_dmem_n11814, MEM_stage_inst_dmem_n11815, MEM_stage_inst_dmem_n11816, MEM_stage_inst_dmem_n11817, MEM_stage_inst_dmem_n11818, MEM_stage_inst_dmem_n11819, MEM_stage_inst_dmem_n11820, MEM_stage_inst_dmem_n11821, MEM_stage_inst_dmem_n11822, MEM_stage_inst_dmem_n11823, MEM_stage_inst_dmem_n11824, MEM_stage_inst_dmem_n11825, MEM_stage_inst_dmem_n11826, MEM_stage_inst_dmem_n11827, MEM_stage_inst_dmem_n11828, MEM_stage_inst_dmem_n11829, MEM_stage_inst_dmem_n11830, MEM_stage_inst_dmem_n11831, MEM_stage_inst_dmem_n11832, MEM_stage_inst_dmem_n11833, MEM_stage_inst_dmem_n11834, MEM_stage_inst_dmem_n11835, MEM_stage_inst_dmem_n11836, MEM_stage_inst_dmem_n11837, MEM_stage_inst_dmem_n11838, MEM_stage_inst_dmem_n11839, MEM_stage_inst_dmem_n11840, MEM_stage_inst_dmem_n11841, MEM_stage_inst_dmem_n11842, MEM_stage_inst_dmem_n11843, MEM_stage_inst_dmem_n11844, MEM_stage_inst_dmem_n11845, MEM_stage_inst_dmem_n11846, MEM_stage_inst_dmem_n11847, MEM_stage_inst_dmem_n11848, MEM_stage_inst_dmem_n11849, MEM_stage_inst_dmem_n11850, MEM_stage_inst_dmem_n11851, MEM_stage_inst_dmem_n11852, MEM_stage_inst_dmem_n11853, MEM_stage_inst_dmem_n11854, MEM_stage_inst_dmem_n11855, MEM_stage_inst_dmem_n11856, MEM_stage_inst_dmem_n11857, MEM_stage_inst_dmem_n11858, MEM_stage_inst_dmem_n11859, MEM_stage_inst_dmem_n11860, MEM_stage_inst_dmem_n11861, MEM_stage_inst_dmem_n11862, MEM_stage_inst_dmem_n11863, MEM_stage_inst_dmem_n11864, MEM_stage_inst_dmem_n11865, MEM_stage_inst_dmem_n11866, MEM_stage_inst_dmem_n11867, MEM_stage_inst_dmem_n11868, MEM_stage_inst_dmem_n11869, MEM_stage_inst_dmem_n11870, MEM_stage_inst_dmem_n11871, MEM_stage_inst_dmem_n11872, MEM_stage_inst_dmem_n11873, MEM_stage_inst_dmem_n11874, MEM_stage_inst_dmem_n11875, MEM_stage_inst_dmem_n11876, MEM_stage_inst_dmem_n11877, MEM_stage_inst_dmem_n11878, MEM_stage_inst_dmem_n11879, MEM_stage_inst_dmem_n11880, MEM_stage_inst_dmem_n11881, MEM_stage_inst_dmem_n11882, MEM_stage_inst_dmem_n11883, MEM_stage_inst_dmem_n11884, MEM_stage_inst_dmem_n11885, MEM_stage_inst_dmem_n11886, MEM_stage_inst_dmem_n11887, MEM_stage_inst_dmem_n11888, MEM_stage_inst_dmem_n11889, MEM_stage_inst_dmem_n11890, MEM_stage_inst_dmem_n11891, MEM_stage_inst_dmem_n11892, MEM_stage_inst_dmem_n11893, MEM_stage_inst_dmem_n11894, MEM_stage_inst_dmem_n11895, MEM_stage_inst_dmem_n11896, MEM_stage_inst_dmem_n11897, MEM_stage_inst_dmem_n11898, MEM_stage_inst_dmem_n11899, MEM_stage_inst_dmem_n11900, MEM_stage_inst_dmem_n11901, MEM_stage_inst_dmem_n11902, MEM_stage_inst_dmem_n11903, MEM_stage_inst_dmem_n11904, MEM_stage_inst_dmem_n11905, MEM_stage_inst_dmem_n11906, MEM_stage_inst_dmem_n11907, MEM_stage_inst_dmem_n11908, MEM_stage_inst_dmem_n11909, MEM_stage_inst_dmem_n11910, MEM_stage_inst_dmem_n11911, MEM_stage_inst_dmem_n11912, MEM_stage_inst_dmem_n11913, MEM_stage_inst_dmem_n11914, MEM_stage_inst_dmem_n11915, MEM_stage_inst_dmem_n11916, MEM_stage_inst_dmem_n11917, MEM_stage_inst_dmem_n11918, MEM_stage_inst_dmem_n11919, MEM_stage_inst_dmem_n11920, MEM_stage_inst_dmem_n11921, MEM_stage_inst_dmem_n11922, MEM_stage_inst_dmem_n11923, MEM_stage_inst_dmem_n11924, MEM_stage_inst_dmem_n11925, MEM_stage_inst_dmem_n11926, MEM_stage_inst_dmem_n11927, MEM_stage_inst_dmem_n11928, MEM_stage_inst_dmem_n11929, MEM_stage_inst_dmem_n11930, MEM_stage_inst_dmem_n11931, MEM_stage_inst_dmem_n11932, MEM_stage_inst_dmem_n11933, MEM_stage_inst_dmem_n11934, MEM_stage_inst_dmem_n11935, MEM_stage_inst_dmem_n11936, MEM_stage_inst_dmem_n11937, MEM_stage_inst_dmem_n11938, MEM_stage_inst_dmem_n11939, MEM_stage_inst_dmem_n11940, MEM_stage_inst_dmem_n11941, MEM_stage_inst_dmem_n11942, MEM_stage_inst_dmem_n11943, MEM_stage_inst_dmem_n11944, MEM_stage_inst_dmem_n11945, MEM_stage_inst_dmem_n11946, MEM_stage_inst_dmem_n11947, MEM_stage_inst_dmem_n11948, MEM_stage_inst_dmem_n11949, MEM_stage_inst_dmem_n11950, MEM_stage_inst_dmem_n11951, MEM_stage_inst_dmem_n11952, MEM_stage_inst_dmem_n11953, MEM_stage_inst_dmem_n11954, MEM_stage_inst_dmem_n11955, MEM_stage_inst_dmem_n11956, MEM_stage_inst_dmem_n11957, MEM_stage_inst_dmem_n11958, MEM_stage_inst_dmem_n11959, MEM_stage_inst_dmem_n11960, MEM_stage_inst_dmem_n11961, MEM_stage_inst_dmem_n11962, MEM_stage_inst_dmem_n11963, MEM_stage_inst_dmem_n11964, MEM_stage_inst_dmem_n11965, MEM_stage_inst_dmem_n11966, MEM_stage_inst_dmem_n11967, MEM_stage_inst_dmem_n11968, MEM_stage_inst_dmem_n11969, MEM_stage_inst_dmem_n11970, MEM_stage_inst_dmem_n11971, MEM_stage_inst_dmem_n11972, MEM_stage_inst_dmem_n11973, MEM_stage_inst_dmem_n11974, MEM_stage_inst_dmem_n11975, MEM_stage_inst_dmem_n11976, MEM_stage_inst_dmem_n11977, MEM_stage_inst_dmem_n11978, MEM_stage_inst_dmem_n11979, MEM_stage_inst_dmem_n11980, MEM_stage_inst_dmem_n11981, MEM_stage_inst_dmem_n11982, MEM_stage_inst_dmem_n11983, MEM_stage_inst_dmem_n11984, MEM_stage_inst_dmem_n11985, MEM_stage_inst_dmem_n11986, MEM_stage_inst_dmem_n11987, MEM_stage_inst_dmem_n11988, MEM_stage_inst_dmem_n11989, MEM_stage_inst_dmem_n11990, MEM_stage_inst_dmem_n11991, MEM_stage_inst_dmem_n11992, MEM_stage_inst_dmem_n11993, MEM_stage_inst_dmem_n11994, MEM_stage_inst_dmem_n11995, MEM_stage_inst_dmem_n11996, MEM_stage_inst_dmem_n11997, MEM_stage_inst_dmem_n11998, MEM_stage_inst_dmem_n11999, MEM_stage_inst_dmem_n12000, MEM_stage_inst_dmem_n12001, MEM_stage_inst_dmem_n12002, MEM_stage_inst_dmem_n12003, MEM_stage_inst_dmem_n12004, MEM_stage_inst_dmem_n12005, MEM_stage_inst_dmem_n12006, MEM_stage_inst_dmem_n12007, MEM_stage_inst_dmem_n12008, MEM_stage_inst_dmem_n12009, MEM_stage_inst_dmem_n12010, MEM_stage_inst_dmem_n12011, MEM_stage_inst_dmem_n12012, MEM_stage_inst_dmem_n12013, MEM_stage_inst_dmem_n12014, MEM_stage_inst_dmem_n12015, MEM_stage_inst_dmem_n12016, MEM_stage_inst_dmem_n12017, MEM_stage_inst_dmem_n12018, MEM_stage_inst_dmem_n12019, MEM_stage_inst_dmem_n12020, MEM_stage_inst_dmem_n12021, MEM_stage_inst_dmem_n12022, MEM_stage_inst_dmem_n12023, MEM_stage_inst_dmem_n12024, MEM_stage_inst_dmem_n12025, MEM_stage_inst_dmem_n12026, MEM_stage_inst_dmem_n12027, MEM_stage_inst_dmem_n12028, MEM_stage_inst_dmem_n12029, MEM_stage_inst_dmem_n12030, MEM_stage_inst_dmem_n12031, MEM_stage_inst_dmem_n12032, MEM_stage_inst_dmem_n12033, MEM_stage_inst_dmem_n12034, MEM_stage_inst_dmem_n12035, MEM_stage_inst_dmem_n12036, MEM_stage_inst_dmem_n12037, MEM_stage_inst_dmem_n12038, MEM_stage_inst_dmem_n12039, MEM_stage_inst_dmem_n12040, MEM_stage_inst_dmem_n12041, MEM_stage_inst_dmem_n12042, MEM_stage_inst_dmem_n12043, MEM_stage_inst_dmem_n12044, MEM_stage_inst_dmem_n12045, MEM_stage_inst_dmem_n12046, MEM_stage_inst_dmem_n12047, MEM_stage_inst_dmem_n12048, MEM_stage_inst_dmem_n12049, MEM_stage_inst_dmem_n12050, MEM_stage_inst_dmem_n12051, MEM_stage_inst_dmem_n12052, MEM_stage_inst_dmem_n12053, MEM_stage_inst_dmem_n12054, MEM_stage_inst_dmem_n12055, MEM_stage_inst_dmem_n12056, MEM_stage_inst_dmem_n12057, MEM_stage_inst_dmem_n12058, MEM_stage_inst_dmem_n12059, MEM_stage_inst_dmem_n12060, MEM_stage_inst_dmem_n12061, MEM_stage_inst_dmem_n12062, MEM_stage_inst_dmem_n12063, MEM_stage_inst_dmem_n12064, MEM_stage_inst_dmem_n12065, MEM_stage_inst_dmem_n12066, MEM_stage_inst_dmem_n12067, MEM_stage_inst_dmem_n12068, MEM_stage_inst_dmem_n12069, MEM_stage_inst_dmem_n12070, MEM_stage_inst_dmem_n12071, MEM_stage_inst_dmem_n12072, MEM_stage_inst_dmem_n12073, MEM_stage_inst_dmem_n12074, MEM_stage_inst_dmem_n12075, MEM_stage_inst_dmem_n12076, MEM_stage_inst_dmem_n12077, MEM_stage_inst_dmem_n12078, MEM_stage_inst_dmem_n12079, MEM_stage_inst_dmem_n12080, MEM_stage_inst_dmem_n12081, MEM_stage_inst_dmem_n12082, MEM_stage_inst_dmem_n12083, MEM_stage_inst_dmem_n12084, MEM_stage_inst_dmem_n12085, MEM_stage_inst_dmem_n12086, MEM_stage_inst_dmem_n12087, MEM_stage_inst_dmem_n12088, MEM_stage_inst_dmem_n12089, MEM_stage_inst_dmem_n12090, MEM_stage_inst_dmem_n12091, MEM_stage_inst_dmem_n12092, MEM_stage_inst_dmem_n12093, MEM_stage_inst_dmem_n12094, MEM_stage_inst_dmem_n12095, MEM_stage_inst_dmem_n12096, MEM_stage_inst_dmem_n12097, MEM_stage_inst_dmem_n12098, MEM_stage_inst_dmem_n12099, MEM_stage_inst_dmem_n12100, MEM_stage_inst_dmem_n12101, MEM_stage_inst_dmem_n12102, MEM_stage_inst_dmem_n12103, MEM_stage_inst_dmem_n12104, MEM_stage_inst_dmem_n12105, MEM_stage_inst_dmem_n12106, MEM_stage_inst_dmem_n12107, MEM_stage_inst_dmem_n12108, MEM_stage_inst_dmem_n12109, MEM_stage_inst_dmem_n12110, MEM_stage_inst_dmem_n12111, MEM_stage_inst_dmem_n12112, MEM_stage_inst_dmem_n12113, MEM_stage_inst_dmem_n12114, MEM_stage_inst_dmem_n12115, MEM_stage_inst_dmem_n12116, MEM_stage_inst_dmem_n12117, MEM_stage_inst_dmem_n12118, MEM_stage_inst_dmem_n12119, MEM_stage_inst_dmem_n12120, MEM_stage_inst_dmem_n12121, MEM_stage_inst_dmem_n12122, MEM_stage_inst_dmem_n12123, MEM_stage_inst_dmem_n12124, MEM_stage_inst_dmem_n12125, MEM_stage_inst_dmem_n12126, MEM_stage_inst_dmem_n12127, MEM_stage_inst_dmem_n12128, MEM_stage_inst_dmem_n12129, MEM_stage_inst_dmem_n12130, MEM_stage_inst_dmem_n12131, MEM_stage_inst_dmem_n12132, MEM_stage_inst_dmem_n12133, MEM_stage_inst_dmem_n12134, MEM_stage_inst_dmem_n12135, MEM_stage_inst_dmem_n12136, MEM_stage_inst_dmem_n12137, MEM_stage_inst_dmem_n12138, MEM_stage_inst_dmem_n12139, MEM_stage_inst_dmem_n12140, MEM_stage_inst_dmem_n12141, MEM_stage_inst_dmem_n12142, MEM_stage_inst_dmem_n12143, MEM_stage_inst_dmem_n12144, MEM_stage_inst_dmem_n12145, MEM_stage_inst_dmem_n12146, MEM_stage_inst_dmem_n12147, MEM_stage_inst_dmem_n12148, MEM_stage_inst_dmem_n12149, MEM_stage_inst_dmem_n12150, MEM_stage_inst_dmem_n12151, MEM_stage_inst_dmem_n12152, MEM_stage_inst_dmem_n12153, MEM_stage_inst_dmem_n12154, MEM_stage_inst_dmem_n12155, MEM_stage_inst_dmem_n12156, MEM_stage_inst_dmem_n12157, MEM_stage_inst_dmem_n12158, MEM_stage_inst_dmem_n12159, MEM_stage_inst_dmem_n12160, MEM_stage_inst_dmem_n12161, MEM_stage_inst_dmem_n12162, MEM_stage_inst_dmem_n12163, MEM_stage_inst_dmem_n12164, MEM_stage_inst_dmem_n12165, MEM_stage_inst_dmem_n12166, MEM_stage_inst_dmem_n12167, MEM_stage_inst_dmem_n12168, MEM_stage_inst_dmem_n12169, MEM_stage_inst_dmem_n12170, MEM_stage_inst_dmem_n12171, MEM_stage_inst_dmem_n12172, MEM_stage_inst_dmem_n12173, MEM_stage_inst_dmem_n12174, MEM_stage_inst_dmem_n12175, MEM_stage_inst_dmem_n12176, MEM_stage_inst_dmem_n12177, MEM_stage_inst_dmem_n12178, MEM_stage_inst_dmem_n12179, MEM_stage_inst_dmem_n12180, MEM_stage_inst_dmem_n12181, MEM_stage_inst_dmem_n12182, MEM_stage_inst_dmem_n12183, MEM_stage_inst_dmem_n12184, MEM_stage_inst_dmem_n12185, MEM_stage_inst_dmem_n12186, MEM_stage_inst_dmem_n12187, MEM_stage_inst_dmem_n12188, MEM_stage_inst_dmem_n12189, MEM_stage_inst_dmem_n12190, MEM_stage_inst_dmem_n12191, MEM_stage_inst_dmem_n12192, MEM_stage_inst_dmem_n12193, MEM_stage_inst_dmem_n12194, MEM_stage_inst_dmem_n12195, MEM_stage_inst_dmem_n12196, MEM_stage_inst_dmem_n12197, MEM_stage_inst_dmem_n12198, MEM_stage_inst_dmem_n12199, MEM_stage_inst_dmem_n12200, MEM_stage_inst_dmem_n12201, MEM_stage_inst_dmem_n12202, MEM_stage_inst_dmem_n12203, MEM_stage_inst_dmem_n12204, MEM_stage_inst_dmem_n12205, MEM_stage_inst_dmem_n12206, MEM_stage_inst_dmem_n12207, MEM_stage_inst_dmem_n12208, MEM_stage_inst_dmem_n12209, MEM_stage_inst_dmem_n12210, MEM_stage_inst_dmem_n12211, MEM_stage_inst_dmem_n12212, MEM_stage_inst_dmem_n12213, MEM_stage_inst_dmem_n12214, MEM_stage_inst_dmem_n12215, MEM_stage_inst_dmem_n12216, MEM_stage_inst_dmem_n12217, MEM_stage_inst_dmem_n12218, MEM_stage_inst_dmem_n12219, MEM_stage_inst_dmem_n12220, MEM_stage_inst_dmem_n12221, MEM_stage_inst_dmem_n12222, MEM_stage_inst_dmem_n12223, MEM_stage_inst_dmem_n12224, MEM_stage_inst_dmem_n12225, MEM_stage_inst_dmem_n12226, MEM_stage_inst_dmem_n12227, MEM_stage_inst_dmem_n12228, MEM_stage_inst_dmem_n12229, MEM_stage_inst_dmem_n12230, MEM_stage_inst_dmem_n12231, MEM_stage_inst_dmem_n12232, MEM_stage_inst_dmem_n12233, MEM_stage_inst_dmem_n12234, MEM_stage_inst_dmem_n12235, MEM_stage_inst_dmem_n12236, MEM_stage_inst_dmem_n12237, MEM_stage_inst_dmem_n12238, MEM_stage_inst_dmem_n12239, MEM_stage_inst_dmem_n12240, MEM_stage_inst_dmem_n12241, MEM_stage_inst_dmem_n12242, MEM_stage_inst_dmem_n12243, MEM_stage_inst_dmem_n12244, MEM_stage_inst_dmem_n12245, MEM_stage_inst_dmem_n12246, MEM_stage_inst_dmem_n12247, MEM_stage_inst_dmem_n12248, MEM_stage_inst_dmem_n12249, MEM_stage_inst_dmem_n12250, MEM_stage_inst_dmem_n12251, MEM_stage_inst_dmem_n12252, MEM_stage_inst_dmem_n12253, MEM_stage_inst_dmem_n12254, MEM_stage_inst_dmem_n12255, MEM_stage_inst_dmem_n12256, MEM_stage_inst_dmem_n12257, MEM_stage_inst_dmem_n12258, MEM_stage_inst_dmem_n12259, MEM_stage_inst_dmem_n12260, MEM_stage_inst_dmem_n12261, MEM_stage_inst_dmem_n12262, MEM_stage_inst_dmem_n12263, MEM_stage_inst_dmem_n12264, MEM_stage_inst_dmem_n12265, MEM_stage_inst_dmem_n12266, MEM_stage_inst_dmem_n12267, MEM_stage_inst_dmem_n12268, MEM_stage_inst_dmem_n12269, MEM_stage_inst_dmem_n12270, MEM_stage_inst_dmem_n12271, MEM_stage_inst_dmem_n12272, MEM_stage_inst_dmem_n12273, MEM_stage_inst_dmem_n12274, MEM_stage_inst_dmem_n12275, MEM_stage_inst_dmem_n12276, MEM_stage_inst_dmem_n12277, MEM_stage_inst_dmem_n12278, MEM_stage_inst_dmem_n12279, MEM_stage_inst_dmem_n12280, MEM_stage_inst_dmem_n12281, MEM_stage_inst_dmem_n12282, MEM_stage_inst_dmem_n12283, MEM_stage_inst_dmem_n12284, MEM_stage_inst_dmem_n12285, MEM_stage_inst_dmem_n12286, MEM_stage_inst_dmem_n12287, MEM_stage_inst_dmem_n12288, MEM_stage_inst_dmem_n12289, MEM_stage_inst_dmem_n12290, MEM_stage_inst_dmem_n12291, MEM_stage_inst_dmem_n12292, MEM_stage_inst_dmem_n12293, MEM_stage_inst_dmem_n12294, MEM_stage_inst_dmem_n12295, MEM_stage_inst_dmem_n12296, MEM_stage_inst_dmem_n12297, MEM_stage_inst_dmem_n12298, MEM_stage_inst_dmem_n12299, MEM_stage_inst_dmem_n12300, MEM_stage_inst_dmem_n12301, MEM_stage_inst_dmem_n12302, MEM_stage_inst_dmem_n12303, MEM_stage_inst_dmem_n12304, MEM_stage_inst_dmem_n12305, MEM_stage_inst_dmem_n12306, MEM_stage_inst_dmem_n12307, MEM_stage_inst_dmem_n12308, MEM_stage_inst_dmem_n12309, MEM_stage_inst_dmem_n12310, MEM_stage_inst_dmem_n12311, MEM_stage_inst_dmem_n12312, MEM_stage_inst_dmem_n12313, MEM_stage_inst_dmem_n12314, MEM_stage_inst_dmem_n12315, MEM_stage_inst_dmem_n12316, MEM_stage_inst_dmem_n12317, MEM_stage_inst_dmem_n12318, MEM_stage_inst_dmem_n12319, MEM_stage_inst_dmem_n12320, MEM_stage_inst_dmem_n12321, MEM_stage_inst_dmem_n12322, MEM_stage_inst_dmem_n12323, MEM_stage_inst_dmem_n12324, MEM_stage_inst_dmem_n12325, MEM_stage_inst_dmem_n12326, MEM_stage_inst_dmem_n12327, MEM_stage_inst_dmem_n12328, MEM_stage_inst_dmem_n12329, MEM_stage_inst_dmem_n12330, MEM_stage_inst_dmem_n12331, MEM_stage_inst_dmem_n12332, MEM_stage_inst_dmem_n12333, MEM_stage_inst_dmem_n12334, MEM_stage_inst_dmem_n12335, MEM_stage_inst_dmem_n12336, MEM_stage_inst_dmem_n12337, MEM_stage_inst_dmem_n12338, MEM_stage_inst_dmem_n12339, MEM_stage_inst_dmem_n12340, MEM_stage_inst_dmem_n12341, MEM_stage_inst_dmem_n12342, MEM_stage_inst_dmem_n12343, MEM_stage_inst_dmem_n12344, MEM_stage_inst_dmem_n12345, MEM_stage_inst_dmem_n12346, MEM_stage_inst_dmem_n12347, MEM_stage_inst_dmem_n12348, MEM_stage_inst_dmem_n12349, MEM_stage_inst_dmem_n12350, MEM_stage_inst_dmem_n12351, MEM_stage_inst_dmem_n12352, MEM_stage_inst_dmem_n12353, MEM_stage_inst_dmem_n12354, MEM_stage_inst_dmem_n12355, MEM_stage_inst_dmem_n12356, MEM_stage_inst_dmem_n12357, MEM_stage_inst_dmem_n12358, MEM_stage_inst_dmem_n12359, MEM_stage_inst_dmem_n12360, MEM_stage_inst_dmem_n12361, MEM_stage_inst_dmem_n12362, MEM_stage_inst_dmem_n12363, MEM_stage_inst_dmem_n12364, MEM_stage_inst_dmem_n12365, MEM_stage_inst_dmem_n12366, MEM_stage_inst_dmem_n12367, MEM_stage_inst_dmem_n12368, MEM_stage_inst_dmem_n12369, MEM_stage_inst_dmem_n12370, MEM_stage_inst_dmem_n12371, MEM_stage_inst_dmem_n12372, MEM_stage_inst_dmem_n12373, MEM_stage_inst_dmem_n12374, MEM_stage_inst_dmem_n12375, MEM_stage_inst_dmem_n12376, MEM_stage_inst_dmem_n12377, MEM_stage_inst_dmem_n12378, MEM_stage_inst_dmem_n12379, MEM_stage_inst_dmem_n12380, MEM_stage_inst_dmem_n12381, MEM_stage_inst_dmem_n12382, MEM_stage_inst_dmem_n12383, MEM_stage_inst_dmem_n12384, MEM_stage_inst_dmem_n12385, MEM_stage_inst_dmem_n12386, MEM_stage_inst_dmem_n12387, MEM_stage_inst_dmem_n12388, MEM_stage_inst_dmem_n12389, MEM_stage_inst_dmem_n12390, MEM_stage_inst_dmem_n12391, MEM_stage_inst_dmem_n12392, MEM_stage_inst_dmem_n12393, MEM_stage_inst_dmem_n12394, MEM_stage_inst_dmem_n12395, MEM_stage_inst_dmem_n12396, MEM_stage_inst_dmem_n12397, MEM_stage_inst_dmem_n12398, MEM_stage_inst_dmem_n12399, MEM_stage_inst_dmem_n12400, MEM_stage_inst_dmem_n12401, MEM_stage_inst_dmem_n12402, MEM_stage_inst_dmem_n12403, MEM_stage_inst_dmem_n12404, MEM_stage_inst_dmem_n12405, MEM_stage_inst_dmem_n12406, MEM_stage_inst_dmem_n12407, MEM_stage_inst_dmem_n12408, MEM_stage_inst_dmem_n12409, MEM_stage_inst_dmem_n12410, MEM_stage_inst_dmem_n12411, MEM_stage_inst_dmem_n12412, MEM_stage_inst_dmem_n12413, MEM_stage_inst_dmem_n12414, MEM_stage_inst_dmem_n12415, MEM_stage_inst_dmem_n12416, MEM_stage_inst_dmem_n12417, MEM_stage_inst_dmem_n12418, MEM_stage_inst_dmem_n12419, MEM_stage_inst_dmem_n12420, MEM_stage_inst_dmem_n12421, MEM_stage_inst_dmem_n12422, MEM_stage_inst_dmem_n12423, MEM_stage_inst_dmem_n12424, MEM_stage_inst_dmem_n12425, MEM_stage_inst_dmem_n12426, MEM_stage_inst_dmem_n12427, MEM_stage_inst_dmem_n12428, MEM_stage_inst_dmem_n12429, MEM_stage_inst_dmem_n12430, MEM_stage_inst_dmem_n12431, MEM_stage_inst_dmem_n12432, MEM_stage_inst_dmem_n12433, MEM_stage_inst_dmem_n12434, MEM_stage_inst_dmem_n12435, MEM_stage_inst_dmem_n12436, MEM_stage_inst_dmem_n12437, MEM_stage_inst_dmem_n12438, MEM_stage_inst_dmem_n12439, MEM_stage_inst_dmem_n12440, MEM_stage_inst_dmem_n12441, MEM_stage_inst_dmem_n12442, MEM_stage_inst_dmem_n12443, MEM_stage_inst_dmem_n12444, MEM_stage_inst_dmem_n12445, MEM_stage_inst_dmem_n12446, MEM_stage_inst_dmem_n12447, MEM_stage_inst_dmem_n12448, MEM_stage_inst_dmem_n12449, MEM_stage_inst_dmem_n12450, MEM_stage_inst_dmem_n12451, MEM_stage_inst_dmem_n12452, MEM_stage_inst_dmem_n12453, MEM_stage_inst_dmem_n12454, MEM_stage_inst_dmem_n12455, MEM_stage_inst_dmem_n12456, MEM_stage_inst_dmem_n12457, MEM_stage_inst_dmem_n12458, MEM_stage_inst_dmem_n12459, MEM_stage_inst_dmem_n12460, MEM_stage_inst_dmem_n12461, MEM_stage_inst_dmem_n12462, MEM_stage_inst_dmem_n12463, MEM_stage_inst_dmem_n12464, MEM_stage_inst_dmem_n12465, MEM_stage_inst_dmem_n12466, MEM_stage_inst_dmem_n12467, MEM_stage_inst_dmem_n12468, MEM_stage_inst_dmem_n12469, MEM_stage_inst_dmem_n12470, MEM_stage_inst_dmem_n12471, MEM_stage_inst_dmem_n12472, MEM_stage_inst_dmem_n12473, MEM_stage_inst_dmem_n12474, MEM_stage_inst_dmem_n12475, MEM_stage_inst_dmem_n12476, MEM_stage_inst_dmem_n12477, MEM_stage_inst_dmem_n12478, MEM_stage_inst_dmem_n12479, MEM_stage_inst_dmem_n12480, MEM_stage_inst_dmem_n12481, MEM_stage_inst_dmem_n12482, MEM_stage_inst_dmem_n12483, MEM_stage_inst_dmem_n12484, MEM_stage_inst_dmem_n12485, MEM_stage_inst_dmem_n12486, MEM_stage_inst_dmem_n12487, MEM_stage_inst_dmem_n12488, MEM_stage_inst_dmem_n12489, MEM_stage_inst_dmem_n12490, MEM_stage_inst_dmem_n12491, MEM_stage_inst_dmem_n12492, MEM_stage_inst_dmem_n12493, MEM_stage_inst_dmem_n12494, MEM_stage_inst_dmem_n12495, MEM_stage_inst_dmem_n12496, MEM_stage_inst_dmem_n12497, MEM_stage_inst_dmem_n12498, MEM_stage_inst_dmem_n12499, MEM_stage_inst_dmem_n12500, MEM_stage_inst_dmem_n12501, MEM_stage_inst_dmem_n12502, MEM_stage_inst_dmem_n12503, MEM_stage_inst_dmem_n12504, MEM_stage_inst_dmem_n12505, MEM_stage_inst_dmem_n12506, MEM_stage_inst_dmem_n12507, MEM_stage_inst_dmem_n12508, MEM_stage_inst_dmem_n12509, MEM_stage_inst_dmem_n12510, MEM_stage_inst_dmem_n12511, MEM_stage_inst_dmem_n12512, MEM_stage_inst_dmem_n12513, MEM_stage_inst_dmem_n12514, MEM_stage_inst_dmem_n12515, MEM_stage_inst_dmem_n12516, MEM_stage_inst_dmem_n12517, MEM_stage_inst_dmem_n12518, MEM_stage_inst_dmem_n12519, MEM_stage_inst_dmem_n12520, MEM_stage_inst_dmem_n12521, MEM_stage_inst_dmem_n12522, MEM_stage_inst_dmem_n12523, MEM_stage_inst_dmem_n12524, MEM_stage_inst_dmem_n12525, MEM_stage_inst_dmem_n12526, MEM_stage_inst_dmem_n12527, MEM_stage_inst_dmem_n12528, MEM_stage_inst_dmem_n12529, MEM_stage_inst_dmem_n12530, MEM_stage_inst_dmem_n12531, MEM_stage_inst_dmem_n12532, MEM_stage_inst_dmem_n12533, MEM_stage_inst_dmem_n12534, MEM_stage_inst_dmem_n12535, MEM_stage_inst_dmem_n12536, MEM_stage_inst_dmem_n12537, MEM_stage_inst_dmem_n12538, MEM_stage_inst_dmem_n12539, MEM_stage_inst_dmem_n12540, MEM_stage_inst_dmem_n12541, MEM_stage_inst_dmem_n12542, MEM_stage_inst_dmem_n12543, MEM_stage_inst_dmem_n12544, MEM_stage_inst_dmem_n12545, MEM_stage_inst_dmem_n12546, MEM_stage_inst_dmem_n12547, MEM_stage_inst_dmem_n12548, MEM_stage_inst_dmem_n12549, MEM_stage_inst_dmem_n12550, MEM_stage_inst_dmem_n12551, MEM_stage_inst_dmem_n12552, MEM_stage_inst_dmem_n12553, MEM_stage_inst_dmem_n12554, MEM_stage_inst_dmem_n12555, MEM_stage_inst_dmem_n12556, MEM_stage_inst_dmem_n12557, MEM_stage_inst_dmem_n12558, MEM_stage_inst_dmem_n12559, MEM_stage_inst_dmem_n12560, MEM_stage_inst_dmem_n12561, MEM_stage_inst_dmem_n12562, MEM_stage_inst_dmem_n12563, MEM_stage_inst_dmem_n12564, MEM_stage_inst_dmem_n12565, MEM_stage_inst_dmem_n12566, MEM_stage_inst_dmem_n12567, MEM_stage_inst_dmem_n12568, MEM_stage_inst_dmem_n12569, MEM_stage_inst_dmem_n12570, MEM_stage_inst_dmem_n12571, MEM_stage_inst_dmem_n12572, MEM_stage_inst_dmem_n12573, MEM_stage_inst_dmem_n12574, MEM_stage_inst_dmem_n12575, MEM_stage_inst_dmem_n12576, MEM_stage_inst_dmem_n12577, MEM_stage_inst_dmem_n12578, MEM_stage_inst_dmem_n12579, MEM_stage_inst_dmem_n12580, MEM_stage_inst_dmem_n12581, MEM_stage_inst_dmem_n12582, MEM_stage_inst_dmem_n12583, MEM_stage_inst_dmem_n12584, MEM_stage_inst_dmem_n12585, MEM_stage_inst_dmem_n12586, MEM_stage_inst_dmem_n12587, MEM_stage_inst_dmem_n12588, MEM_stage_inst_dmem_n12589, MEM_stage_inst_dmem_n12590, MEM_stage_inst_dmem_n12591, MEM_stage_inst_dmem_n12592, MEM_stage_inst_dmem_n12593, MEM_stage_inst_dmem_n12594, MEM_stage_inst_dmem_n12595, MEM_stage_inst_dmem_n12596, MEM_stage_inst_dmem_n12597, MEM_stage_inst_dmem_n12598, MEM_stage_inst_dmem_n12599, MEM_stage_inst_dmem_n12600, MEM_stage_inst_dmem_n12601, MEM_stage_inst_dmem_n12602, MEM_stage_inst_dmem_n12603, MEM_stage_inst_dmem_n12604, MEM_stage_inst_dmem_n12605, MEM_stage_inst_dmem_n12606, MEM_stage_inst_dmem_n12607, MEM_stage_inst_dmem_n12608, MEM_stage_inst_dmem_n12609, MEM_stage_inst_dmem_n12610, MEM_stage_inst_dmem_n12611, MEM_stage_inst_dmem_n12612, MEM_stage_inst_dmem_n12613, MEM_stage_inst_dmem_n12614, MEM_stage_inst_dmem_n12615, MEM_stage_inst_dmem_n12616, MEM_stage_inst_dmem_n12617, MEM_stage_inst_dmem_n12618, MEM_stage_inst_dmem_n12619, MEM_stage_inst_dmem_n12620, MEM_stage_inst_dmem_n12621, MEM_stage_inst_dmem_n12622, MEM_stage_inst_dmem_n12623, MEM_stage_inst_dmem_n12624, MEM_stage_inst_dmem_n12625, MEM_stage_inst_dmem_n12626, MEM_stage_inst_dmem_n12627, MEM_stage_inst_dmem_n12628, MEM_stage_inst_dmem_n12629, MEM_stage_inst_dmem_n12630, MEM_stage_inst_dmem_n12631, MEM_stage_inst_dmem_n12632, MEM_stage_inst_dmem_n12633, MEM_stage_inst_dmem_n12634, MEM_stage_inst_dmem_n12635, MEM_stage_inst_dmem_n12636, MEM_stage_inst_dmem_n12637, MEM_stage_inst_dmem_n12638, MEM_stage_inst_dmem_n12639, MEM_stage_inst_dmem_n12640, MEM_stage_inst_dmem_n12641, MEM_stage_inst_dmem_n12642, MEM_stage_inst_dmem_n12643, MEM_stage_inst_dmem_n12644, MEM_stage_inst_dmem_n12645, MEM_stage_inst_dmem_n12646, MEM_stage_inst_dmem_n12647, MEM_stage_inst_dmem_n12648, MEM_stage_inst_dmem_n12649, MEM_stage_inst_dmem_n12650, MEM_stage_inst_dmem_n12651, MEM_stage_inst_dmem_n12652, MEM_stage_inst_dmem_n12653, MEM_stage_inst_dmem_n12654, MEM_stage_inst_dmem_n12655, MEM_stage_inst_dmem_n12656, MEM_stage_inst_dmem_n12657, MEM_stage_inst_dmem_n12658, MEM_stage_inst_dmem_n12659, MEM_stage_inst_dmem_n12660, MEM_stage_inst_dmem_n12661, MEM_stage_inst_dmem_n12662, MEM_stage_inst_dmem_n12663, MEM_stage_inst_dmem_n12664, MEM_stage_inst_dmem_n12665, MEM_stage_inst_dmem_n12666, MEM_stage_inst_dmem_n12667, MEM_stage_inst_dmem_n12668, MEM_stage_inst_dmem_n12669, MEM_stage_inst_dmem_n12670, MEM_stage_inst_dmem_n12671, MEM_stage_inst_dmem_n12672, MEM_stage_inst_dmem_n12673, MEM_stage_inst_dmem_n12674, MEM_stage_inst_dmem_n12675, MEM_stage_inst_dmem_n12676, MEM_stage_inst_dmem_n12677, MEM_stage_inst_dmem_n12678, MEM_stage_inst_dmem_n12679, MEM_stage_inst_dmem_n12680, MEM_stage_inst_dmem_n12681, MEM_stage_inst_dmem_n12682, MEM_stage_inst_dmem_n12683, MEM_stage_inst_dmem_n12684, MEM_stage_inst_dmem_n12685, MEM_stage_inst_dmem_n12686, MEM_stage_inst_dmem_n12687, MEM_stage_inst_dmem_n12688, MEM_stage_inst_dmem_n12689, MEM_stage_inst_dmem_n12690, MEM_stage_inst_dmem_n12691, MEM_stage_inst_dmem_n12692, MEM_stage_inst_dmem_n12693, MEM_stage_inst_dmem_n12694, MEM_stage_inst_dmem_n12695, MEM_stage_inst_dmem_n12696, MEM_stage_inst_dmem_n12697, MEM_stage_inst_dmem_n12698, MEM_stage_inst_dmem_n12699, MEM_stage_inst_dmem_n12700, MEM_stage_inst_dmem_n12701, MEM_stage_inst_dmem_n12702, MEM_stage_inst_dmem_n12703, MEM_stage_inst_dmem_n12704, MEM_stage_inst_dmem_n12705, MEM_stage_inst_dmem_n12706, MEM_stage_inst_dmem_n12707, MEM_stage_inst_dmem_n12708, MEM_stage_inst_dmem_n12709, MEM_stage_inst_dmem_n12710, MEM_stage_inst_dmem_n12711, MEM_stage_inst_dmem_n12712, MEM_stage_inst_dmem_n12713, MEM_stage_inst_dmem_n12714, MEM_stage_inst_dmem_n12715, MEM_stage_inst_dmem_n12716, MEM_stage_inst_dmem_n12717, MEM_stage_inst_dmem_n12718, MEM_stage_inst_dmem_n12719, MEM_stage_inst_dmem_n12720, MEM_stage_inst_dmem_n12721, MEM_stage_inst_dmem_n12722, MEM_stage_inst_dmem_n12723, MEM_stage_inst_dmem_n12724, MEM_stage_inst_dmem_n12725, MEM_stage_inst_dmem_n12726, MEM_stage_inst_dmem_n12727, MEM_stage_inst_dmem_n12728, MEM_stage_inst_dmem_n12729, MEM_stage_inst_dmem_n12730, MEM_stage_inst_dmem_n12731, MEM_stage_inst_dmem_n12732, MEM_stage_inst_dmem_n12733, MEM_stage_inst_dmem_n12734, MEM_stage_inst_dmem_n12735, MEM_stage_inst_dmem_n12736, MEM_stage_inst_dmem_n12737, MEM_stage_inst_dmem_n12738, MEM_stage_inst_dmem_n12739, MEM_stage_inst_dmem_n12740, MEM_stage_inst_dmem_n12741, MEM_stage_inst_dmem_n12742, MEM_stage_inst_dmem_n12743, MEM_stage_inst_dmem_n12744, MEM_stage_inst_dmem_n12745, MEM_stage_inst_dmem_n12746, MEM_stage_inst_dmem_n12747, MEM_stage_inst_dmem_n12748, MEM_stage_inst_dmem_n12749, MEM_stage_inst_dmem_n12750, MEM_stage_inst_dmem_n12751, MEM_stage_inst_dmem_n12752, MEM_stage_inst_dmem_n12753, MEM_stage_inst_dmem_n12754, MEM_stage_inst_dmem_n12755, MEM_stage_inst_dmem_n12756, MEM_stage_inst_dmem_n12757, MEM_stage_inst_dmem_n12758, MEM_stage_inst_dmem_n12759, MEM_stage_inst_dmem_n12760, MEM_stage_inst_dmem_n12761, MEM_stage_inst_dmem_n12762, MEM_stage_inst_dmem_n12763, MEM_stage_inst_dmem_n12764, MEM_stage_inst_dmem_n12765, MEM_stage_inst_dmem_n12766, MEM_stage_inst_dmem_n12767, MEM_stage_inst_dmem_n12768, MEM_stage_inst_dmem_n12769, MEM_stage_inst_dmem_n12770, MEM_stage_inst_dmem_n12771, MEM_stage_inst_dmem_n12772, MEM_stage_inst_dmem_n12773, MEM_stage_inst_dmem_n12774, MEM_stage_inst_dmem_n12775, MEM_stage_inst_dmem_n12776, MEM_stage_inst_dmem_n12777, MEM_stage_inst_dmem_n12778, MEM_stage_inst_dmem_n12779, MEM_stage_inst_dmem_n12780, MEM_stage_inst_dmem_n12781, MEM_stage_inst_dmem_n12782, MEM_stage_inst_dmem_n12783, MEM_stage_inst_dmem_n12784, MEM_stage_inst_dmem_n12785, MEM_stage_inst_dmem_n12786, MEM_stage_inst_dmem_n12787, MEM_stage_inst_dmem_n12788, MEM_stage_inst_dmem_n12789, MEM_stage_inst_dmem_n12790, MEM_stage_inst_dmem_n12791, MEM_stage_inst_dmem_n12792, MEM_stage_inst_dmem_n12793, MEM_stage_inst_dmem_n12794, MEM_stage_inst_dmem_n12795, MEM_stage_inst_dmem_n12796, MEM_stage_inst_dmem_n12797, MEM_stage_inst_dmem_n12798, MEM_stage_inst_dmem_n12799, MEM_stage_inst_dmem_n12800, MEM_stage_inst_dmem_n12801, MEM_stage_inst_dmem_n12802, MEM_stage_inst_dmem_n12803, MEM_stage_inst_dmem_n12804, MEM_stage_inst_dmem_n12805, MEM_stage_inst_dmem_n12806, MEM_stage_inst_dmem_n12807, MEM_stage_inst_dmem_n12808, MEM_stage_inst_dmem_n12809, MEM_stage_inst_dmem_n12810, MEM_stage_inst_dmem_n12811, MEM_stage_inst_dmem_n12812, MEM_stage_inst_dmem_n12813, MEM_stage_inst_dmem_n12814, MEM_stage_inst_dmem_n12815, MEM_stage_inst_dmem_n12816, MEM_stage_inst_dmem_n12817, MEM_stage_inst_dmem_n12818, MEM_stage_inst_dmem_n12819, MEM_stage_inst_dmem_n12820, MEM_stage_inst_dmem_n12821, MEM_stage_inst_dmem_n12822, MEM_stage_inst_dmem_n12823, MEM_stage_inst_dmem_n12824, MEM_stage_inst_dmem_n12825, MEM_stage_inst_dmem_n12826, MEM_stage_inst_dmem_n12827, MEM_stage_inst_dmem_n12828, MEM_stage_inst_dmem_n12829, MEM_stage_inst_dmem_n12830, MEM_stage_inst_dmem_n12831, MEM_stage_inst_dmem_n12832, MEM_stage_inst_dmem_n12833, MEM_stage_inst_dmem_n12834, MEM_stage_inst_dmem_n12835, MEM_stage_inst_dmem_n12836, MEM_stage_inst_dmem_n12837, MEM_stage_inst_dmem_n12838, MEM_stage_inst_dmem_n12839, MEM_stage_inst_dmem_n12840, MEM_stage_inst_dmem_n12841, MEM_stage_inst_dmem_n12842, MEM_stage_inst_dmem_n12843, MEM_stage_inst_dmem_n12844, MEM_stage_inst_dmem_n12845, MEM_stage_inst_dmem_n12846, MEM_stage_inst_dmem_n12847, MEM_stage_inst_dmem_n12848, MEM_stage_inst_dmem_n12849, MEM_stage_inst_dmem_n12850, MEM_stage_inst_dmem_n12851, MEM_stage_inst_dmem_n12852, MEM_stage_inst_dmem_n12853, MEM_stage_inst_dmem_n12854, MEM_stage_inst_dmem_n12855, MEM_stage_inst_dmem_n12856, MEM_stage_inst_dmem_n12857, MEM_stage_inst_dmem_n12858, reg_write_dest_2, n3475, mem_op_dest_0, reg_write_dest_0, mem_op_dest_1, reg_write_dest_1, n3484, mem_op_dest_2, EX_pipeline_reg_out_0, EX_pipeline_reg_out_4, n3522, reg_write_en, n3516, EX_pipeline_reg_out_37, MEM_pipeline_reg_out_36, EX_pipeline_reg_out_20, EX_pipeline_reg_out_22, MEM_pipeline_reg_out_21, EX_pipeline_reg_out_5, EX_pipeline_reg_out_30, MEM_pipeline_reg_out_29, EX_pipeline_reg_out_13, EX_pipeline_reg_out_32, MEM_pipeline_reg_out_31, EX_pipeline_reg_out_15, EX_pipeline_reg_out_34, MEM_pipeline_reg_out_33, EX_pipeline_reg_out_17, EX_pipeline_reg_out_36, MEM_pipeline_reg_out_35, EX_pipeline_reg_out_19, EX_pipeline_reg_out_26, MEM_pipeline_reg_out_25, EX_pipeline_reg_out_9, EX_pipeline_reg_out_28, MEM_pipeline_reg_out_27, EX_pipeline_reg_out_11, EX_pipeline_reg_out_33, MEM_pipeline_reg_out_32, EX_pipeline_reg_out_16, EX_pipeline_reg_out_35, MEM_pipeline_reg_out_34, EX_pipeline_reg_out_18, EX_pipeline_reg_out_24, MEM_pipeline_reg_out_23, EX_pipeline_reg_out_7, EX_pipeline_reg_out_25, MEM_pipeline_reg_out_24, EX_pipeline_reg_out_8, EX_pipeline_reg_out_23, MEM_pipeline_reg_out_22, EX_pipeline_reg_out_6, EX_pipeline_reg_out_27, MEM_pipeline_reg_out_26, EX_pipeline_reg_out_10, EX_pipeline_reg_out_31, MEM_pipeline_reg_out_30, EX_pipeline_reg_out_14, EX_pipeline_reg_out_29, MEM_pipeline_reg_out_28, EX_pipeline_reg_out_12, MEM_pipeline_reg_out_5, MEM_pipeline_reg_out_6, MEM_pipeline_reg_out_7, MEM_pipeline_reg_out_8, MEM_pipeline_reg_out_9, MEM_pipeline_reg_out_10, MEM_pipeline_reg_out_11, MEM_pipeline_reg_out_12, MEM_pipeline_reg_out_13, MEM_pipeline_reg_out_14, MEM_pipeline_reg_out_15, MEM_pipeline_reg_out_16, MEM_pipeline_reg_out_17, MEM_pipeline_reg_out_18, MEM_pipeline_reg_out_19, MEM_pipeline_reg_out_20, n3511, branch_offset_imm_3, n3513, branch_offset_imm_5, n3509, branch_offset_imm_1, n3514, branch_offset_imm_4, n3512, ID_stage_inst_instruction_reg_14, n3510, ID_stage_inst_instruction_reg_13, branch_offset_imm_0, reg_read_addr_1_0, reg_read_addr_1_1, n3480, reg_read_addr_1_2, n3479, ID_stage_inst_instruction_reg_9, ex_op_dest_0, ID_stage_inst_instruction_reg_10, n3515, ex_op_dest_1, ID_stage_inst_instruction_reg_11, ex_op_dest_2, ID_stage_inst_instruction_reg_12, n3487, ID_stage_inst_instruction_reg_15, ID_pipeline_reg_out_55, ID_pipeline_reg_out_54, n3473, ID_pipeline_reg_out_56, n3488, ID_pipeline_reg_out_0, ID_pipeline_reg_out_4, ID_pipeline_reg_out_21, register_file_inst_reg_array_111, ID_pipeline_reg_out_53, n3485, register_file_inst_reg_array_95, register_file_inst_reg_array_79, register_file_inst_reg_array_63, n3492, register_file_inst_reg_array_47, register_file_inst_reg_array_31, register_file_inst_reg_array_15, ID_pipeline_reg_out_20, ID_pipeline_reg_out_37, register_file_inst_reg_array_96, register_file_inst_reg_array_80, register_file_inst_reg_array_64, register_file_inst_reg_array_48, n3491, register_file_inst_reg_array_32, register_file_inst_reg_array_16, register_file_inst_reg_array_0, ID_pipeline_reg_out_5, ID_pipeline_reg_out_38, n3486, register_file_inst_reg_array_104, register_file_inst_reg_array_88, register_file_inst_reg_array_72, register_file_inst_reg_array_56, n3500, register_file_inst_reg_array_40, register_file_inst_reg_array_24, register_file_inst_reg_array_8, ID_pipeline_reg_out_13, ID_pipeline_reg_out_30, ID_pipeline_reg_out_46, register_file_inst_reg_array_106, register_file_inst_reg_array_90, register_file_inst_reg_array_74, register_file_inst_reg_array_58, n3504, register_file_inst_reg_array_42, register_file_inst_reg_array_26, register_file_inst_reg_array_10, ID_pipeline_reg_out_15, ID_pipeline_reg_out_32, ID_pipeline_reg_out_48, register_file_inst_reg_array_108, register_file_inst_reg_array_92, register_file_inst_reg_array_76, register_file_inst_reg_array_60, n3495, register_file_inst_reg_array_44, register_file_inst_reg_array_28, register_file_inst_reg_array_12, ID_pipeline_reg_out_17, ID_pipeline_reg_out_34, ID_pipeline_reg_out_50, register_file_inst_reg_array_110, register_file_inst_reg_array_94, register_file_inst_reg_array_78, register_file_inst_reg_array_62, n3501, register_file_inst_reg_array_46, register_file_inst_reg_array_30, register_file_inst_reg_array_14, ID_pipeline_reg_out_19, ID_pipeline_reg_out_36, ID_pipeline_reg_out_52, register_file_inst_reg_array_100, register_file_inst_reg_array_84, register_file_inst_reg_array_68, register_file_inst_reg_array_52, n3496, register_file_inst_reg_array_36, register_file_inst_reg_array_20, register_file_inst_reg_array_4, ID_pipeline_reg_out_9, ID_pipeline_reg_out_26, n3474, ID_pipeline_reg_out_42, register_file_inst_reg_array_102, register_file_inst_reg_array_86, register_file_inst_reg_array_70, register_file_inst_reg_array_54, n3503, register_file_inst_reg_array_38, register_file_inst_reg_array_22, register_file_inst_reg_array_6, ID_pipeline_reg_out_11, ID_pipeline_reg_out_28, ID_pipeline_reg_out_44, register_file_inst_reg_array_107, register_file_inst_reg_array_91, register_file_inst_reg_array_75, register_file_inst_reg_array_59, n3498, register_file_inst_reg_array_43, register_file_inst_reg_array_27, register_file_inst_reg_array_11, ID_pipeline_reg_out_16, ID_pipeline_reg_out_33, ID_pipeline_reg_out_49, register_file_inst_reg_array_109, register_file_inst_reg_array_93, register_file_inst_reg_array_77, register_file_inst_reg_array_61, n3502, register_file_inst_reg_array_45, register_file_inst_reg_array_29, register_file_inst_reg_array_13, ID_pipeline_reg_out_18, ID_pipeline_reg_out_35, ID_pipeline_reg_out_51, n3483, register_file_inst_reg_array_98, register_file_inst_reg_array_82, register_file_inst_reg_array_66, register_file_inst_reg_array_50, n3494, register_file_inst_reg_array_34, register_file_inst_reg_array_18, register_file_inst_reg_array_2, ID_pipeline_reg_out_7, ID_pipeline_reg_out_40, n3508, register_file_inst_reg_array_99, register_file_inst_reg_array_83, register_file_inst_reg_array_67, register_file_inst_reg_array_51, n3506, register_file_inst_reg_array_35, register_file_inst_reg_array_19, register_file_inst_reg_array_3, ID_pipeline_reg_out_8, ID_pipeline_reg_out_41, n3482, register_file_inst_reg_array_97, register_file_inst_reg_array_81, register_file_inst_reg_array_65, register_file_inst_reg_array_49, n3499, register_file_inst_reg_array_33, register_file_inst_reg_array_17, register_file_inst_reg_array_1, ID_pipeline_reg_out_6, ID_pipeline_reg_out_39, register_file_inst_reg_array_101, register_file_inst_reg_array_85, register_file_inst_reg_array_69, register_file_inst_reg_array_53, n3497, register_file_inst_reg_array_37, register_file_inst_reg_array_21, register_file_inst_reg_array_5, ID_pipeline_reg_out_10, ID_pipeline_reg_out_27, ID_pipeline_reg_out_43, n3489, register_file_inst_reg_array_105, register_file_inst_reg_array_89, register_file_inst_reg_array_73, register_file_inst_reg_array_57, n3493, register_file_inst_reg_array_41, register_file_inst_reg_array_25, register_file_inst_reg_array_9, ID_pipeline_reg_out_14, ID_pipeline_reg_out_31, ID_pipeline_reg_out_47, n3490, register_file_inst_reg_array_103, register_file_inst_reg_array_87, register_file_inst_reg_array_71, register_file_inst_reg_array_55, n3505, register_file_inst_reg_array_39, register_file_inst_reg_array_23, register_file_inst_reg_array_7, ID_pipeline_reg_out_12, ID_pipeline_reg_out_29, ID_pipeline_reg_out_45, n3507, n3481, ID_pipeline_reg_out_23, n3478, MEM_pipeline_reg_out_0, n3477, ID_pipeline_reg_out_24, n3476, ID_pipeline_reg_out_22, n3472, ID_pipeline_reg_out_25, n3471, MEM_stage_inst_dmem_ram_3584, MEM_stage_inst_dmem_ram_3585, MEM_stage_inst_dmem_ram_3586, MEM_stage_inst_dmem_ram_3587, MEM_stage_inst_dmem_ram_3588, MEM_stage_inst_dmem_ram_3589, MEM_stage_inst_dmem_ram_3590, MEM_stage_inst_dmem_ram_3591, MEM_stage_inst_dmem_ram_3592, MEM_stage_inst_dmem_ram_3593, MEM_stage_inst_dmem_ram_3594, MEM_stage_inst_dmem_ram_3595, MEM_stage_inst_dmem_ram_3596, MEM_stage_inst_dmem_ram_3597, MEM_stage_inst_dmem_ram_3598, MEM_stage_inst_dmem_ram_3599, MEM_stage_inst_dmem_ram_3600, MEM_stage_inst_dmem_ram_3601, MEM_stage_inst_dmem_ram_3602, MEM_stage_inst_dmem_ram_3603, MEM_stage_inst_dmem_ram_3604, MEM_stage_inst_dmem_ram_3605, MEM_stage_inst_dmem_ram_3606, MEM_stage_inst_dmem_ram_3607, MEM_stage_inst_dmem_ram_3608, MEM_stage_inst_dmem_ram_3609, MEM_stage_inst_dmem_ram_3610, MEM_stage_inst_dmem_ram_3611, MEM_stage_inst_dmem_ram_3612, MEM_stage_inst_dmem_ram_3613, MEM_stage_inst_dmem_ram_3614, MEM_stage_inst_dmem_ram_3615, MEM_stage_inst_dmem_ram_3616, MEM_stage_inst_dmem_ram_3617, MEM_stage_inst_dmem_ram_3618, MEM_stage_inst_dmem_ram_3619, MEM_stage_inst_dmem_ram_3620, MEM_stage_inst_dmem_ram_3621, MEM_stage_inst_dmem_ram_3622, MEM_stage_inst_dmem_ram_3623, MEM_stage_inst_dmem_ram_3624, MEM_stage_inst_dmem_ram_3625, MEM_stage_inst_dmem_ram_3626, MEM_stage_inst_dmem_ram_3627, MEM_stage_inst_dmem_ram_3628, MEM_stage_inst_dmem_ram_3629, MEM_stage_inst_dmem_ram_3630, MEM_stage_inst_dmem_ram_3631, MEM_stage_inst_dmem_ram_3632, MEM_stage_inst_dmem_ram_3633, MEM_stage_inst_dmem_ram_3634, MEM_stage_inst_dmem_ram_3635, MEM_stage_inst_dmem_ram_3636, MEM_stage_inst_dmem_ram_3637, MEM_stage_inst_dmem_ram_3638, MEM_stage_inst_dmem_ram_3639, MEM_stage_inst_dmem_ram_3640, MEM_stage_inst_dmem_ram_3641, MEM_stage_inst_dmem_ram_3642, MEM_stage_inst_dmem_ram_3643, MEM_stage_inst_dmem_ram_3644, MEM_stage_inst_dmem_ram_3645, MEM_stage_inst_dmem_ram_3646, MEM_stage_inst_dmem_ram_3647, MEM_stage_inst_dmem_ram_3648, MEM_stage_inst_dmem_ram_3649, MEM_stage_inst_dmem_ram_3650, MEM_stage_inst_dmem_ram_3651, MEM_stage_inst_dmem_ram_3652, MEM_stage_inst_dmem_ram_3653, MEM_stage_inst_dmem_ram_3654, MEM_stage_inst_dmem_ram_3655, MEM_stage_inst_dmem_ram_3656, MEM_stage_inst_dmem_ram_3657, MEM_stage_inst_dmem_ram_3658, MEM_stage_inst_dmem_ram_3659, MEM_stage_inst_dmem_ram_3660, MEM_stage_inst_dmem_ram_3661, MEM_stage_inst_dmem_ram_3662, MEM_stage_inst_dmem_ram_3663, MEM_stage_inst_dmem_ram_3664, MEM_stage_inst_dmem_ram_3665, MEM_stage_inst_dmem_ram_3666, MEM_stage_inst_dmem_ram_3667, MEM_stage_inst_dmem_ram_3668, MEM_stage_inst_dmem_ram_3669, MEM_stage_inst_dmem_ram_3670, MEM_stage_inst_dmem_ram_3671, MEM_stage_inst_dmem_ram_3672, MEM_stage_inst_dmem_ram_3673, MEM_stage_inst_dmem_ram_3674, MEM_stage_inst_dmem_ram_3675, MEM_stage_inst_dmem_ram_3676, MEM_stage_inst_dmem_ram_3677, MEM_stage_inst_dmem_ram_3678, MEM_stage_inst_dmem_ram_3679, MEM_stage_inst_dmem_ram_3680, MEM_stage_inst_dmem_ram_3681, MEM_stage_inst_dmem_ram_3682, MEM_stage_inst_dmem_ram_3683, MEM_stage_inst_dmem_ram_3684, MEM_stage_inst_dmem_ram_3685, MEM_stage_inst_dmem_ram_3686, MEM_stage_inst_dmem_ram_3687, MEM_stage_inst_dmem_ram_3688, MEM_stage_inst_dmem_ram_3689, MEM_stage_inst_dmem_ram_3690, MEM_stage_inst_dmem_ram_3691, MEM_stage_inst_dmem_ram_3692, MEM_stage_inst_dmem_ram_3693, MEM_stage_inst_dmem_ram_3694, MEM_stage_inst_dmem_ram_3695, MEM_stage_inst_dmem_ram_3696, MEM_stage_inst_dmem_ram_3697, MEM_stage_inst_dmem_ram_3698, MEM_stage_inst_dmem_ram_3699, MEM_stage_inst_dmem_ram_3700, MEM_stage_inst_dmem_ram_3701, MEM_stage_inst_dmem_ram_3702, MEM_stage_inst_dmem_ram_3703, MEM_stage_inst_dmem_ram_3704, MEM_stage_inst_dmem_ram_3705, MEM_stage_inst_dmem_ram_3706, MEM_stage_inst_dmem_ram_3707, MEM_stage_inst_dmem_ram_3708, MEM_stage_inst_dmem_ram_3709, MEM_stage_inst_dmem_ram_3710, MEM_stage_inst_dmem_ram_3711, MEM_stage_inst_dmem_ram_3712, MEM_stage_inst_dmem_ram_3713, MEM_stage_inst_dmem_ram_3714, MEM_stage_inst_dmem_ram_3715, MEM_stage_inst_dmem_ram_3716, MEM_stage_inst_dmem_ram_3717, MEM_stage_inst_dmem_ram_3718, MEM_stage_inst_dmem_ram_3719, MEM_stage_inst_dmem_ram_3720, MEM_stage_inst_dmem_ram_3721, MEM_stage_inst_dmem_ram_3722, MEM_stage_inst_dmem_ram_3723, MEM_stage_inst_dmem_ram_3724, MEM_stage_inst_dmem_ram_3725, MEM_stage_inst_dmem_ram_3726, MEM_stage_inst_dmem_ram_3727, MEM_stage_inst_dmem_ram_3728, MEM_stage_inst_dmem_ram_3729, MEM_stage_inst_dmem_ram_3730, MEM_stage_inst_dmem_ram_3731, MEM_stage_inst_dmem_ram_3732, MEM_stage_inst_dmem_ram_3733, MEM_stage_inst_dmem_ram_3734, MEM_stage_inst_dmem_ram_3735, MEM_stage_inst_dmem_ram_3736, MEM_stage_inst_dmem_ram_3737, MEM_stage_inst_dmem_ram_3738, MEM_stage_inst_dmem_ram_3739, MEM_stage_inst_dmem_ram_3740, MEM_stage_inst_dmem_ram_3741, MEM_stage_inst_dmem_ram_3742, MEM_stage_inst_dmem_ram_3743, MEM_stage_inst_dmem_ram_3744, MEM_stage_inst_dmem_ram_3745, MEM_stage_inst_dmem_ram_3746, MEM_stage_inst_dmem_ram_3747, MEM_stage_inst_dmem_ram_3748, MEM_stage_inst_dmem_ram_3749, MEM_stage_inst_dmem_ram_3750, MEM_stage_inst_dmem_ram_3751, MEM_stage_inst_dmem_ram_3752, MEM_stage_inst_dmem_ram_3753, MEM_stage_inst_dmem_ram_3754, MEM_stage_inst_dmem_ram_3755, MEM_stage_inst_dmem_ram_3756, MEM_stage_inst_dmem_ram_3757, MEM_stage_inst_dmem_ram_3758, MEM_stage_inst_dmem_ram_3759, MEM_stage_inst_dmem_ram_3760, MEM_stage_inst_dmem_ram_3761, MEM_stage_inst_dmem_ram_3762, MEM_stage_inst_dmem_ram_3763, MEM_stage_inst_dmem_ram_3764, MEM_stage_inst_dmem_ram_3765, MEM_stage_inst_dmem_ram_3766, MEM_stage_inst_dmem_ram_3767, MEM_stage_inst_dmem_ram_3768, MEM_stage_inst_dmem_ram_3769, MEM_stage_inst_dmem_ram_3770, MEM_stage_inst_dmem_ram_3771, MEM_stage_inst_dmem_ram_3772, MEM_stage_inst_dmem_ram_3773, MEM_stage_inst_dmem_ram_3774, MEM_stage_inst_dmem_ram_3775, MEM_stage_inst_dmem_ram_3776, MEM_stage_inst_dmem_ram_3777, MEM_stage_inst_dmem_ram_3778, MEM_stage_inst_dmem_ram_3779, MEM_stage_inst_dmem_ram_3780, MEM_stage_inst_dmem_ram_3781, MEM_stage_inst_dmem_ram_3782, MEM_stage_inst_dmem_ram_3783, MEM_stage_inst_dmem_ram_3784, MEM_stage_inst_dmem_ram_3785, MEM_stage_inst_dmem_ram_3786, MEM_stage_inst_dmem_ram_3787, MEM_stage_inst_dmem_ram_3788, MEM_stage_inst_dmem_ram_3789, MEM_stage_inst_dmem_ram_3790, MEM_stage_inst_dmem_ram_3791, MEM_stage_inst_dmem_ram_3792, MEM_stage_inst_dmem_ram_3793, MEM_stage_inst_dmem_ram_3794, MEM_stage_inst_dmem_ram_3795, MEM_stage_inst_dmem_ram_3796, MEM_stage_inst_dmem_ram_3797, MEM_stage_inst_dmem_ram_3798, MEM_stage_inst_dmem_ram_3799, MEM_stage_inst_dmem_ram_3800, MEM_stage_inst_dmem_ram_3801, MEM_stage_inst_dmem_ram_3802, MEM_stage_inst_dmem_ram_3803, MEM_stage_inst_dmem_ram_3804, MEM_stage_inst_dmem_ram_3805, MEM_stage_inst_dmem_ram_3806, MEM_stage_inst_dmem_ram_3807, MEM_stage_inst_dmem_ram_3808, MEM_stage_inst_dmem_ram_3809, MEM_stage_inst_dmem_ram_3810, MEM_stage_inst_dmem_ram_3811, MEM_stage_inst_dmem_ram_3812, MEM_stage_inst_dmem_ram_3813, MEM_stage_inst_dmem_ram_3814, MEM_stage_inst_dmem_ram_3815, MEM_stage_inst_dmem_ram_3816, MEM_stage_inst_dmem_ram_3817, MEM_stage_inst_dmem_ram_3818, MEM_stage_inst_dmem_ram_3819, MEM_stage_inst_dmem_ram_3820, MEM_stage_inst_dmem_ram_3821, MEM_stage_inst_dmem_ram_3822, MEM_stage_inst_dmem_ram_3823, MEM_stage_inst_dmem_ram_3824, MEM_stage_inst_dmem_ram_3825, MEM_stage_inst_dmem_ram_3826, MEM_stage_inst_dmem_ram_3827, MEM_stage_inst_dmem_ram_3828, MEM_stage_inst_dmem_ram_3829, MEM_stage_inst_dmem_ram_3830, MEM_stage_inst_dmem_ram_3831, MEM_stage_inst_dmem_ram_3832, MEM_stage_inst_dmem_ram_3833, MEM_stage_inst_dmem_ram_3834, MEM_stage_inst_dmem_ram_3835, MEM_stage_inst_dmem_ram_3836, MEM_stage_inst_dmem_ram_3837, MEM_stage_inst_dmem_ram_3838, MEM_stage_inst_dmem_ram_3839, MEM_stage_inst_dmem_ram_3840, MEM_stage_inst_dmem_ram_3841, MEM_stage_inst_dmem_ram_3842, MEM_stage_inst_dmem_ram_3843, MEM_stage_inst_dmem_ram_3844, MEM_stage_inst_dmem_ram_3845, MEM_stage_inst_dmem_ram_3846, MEM_stage_inst_dmem_ram_3847, MEM_stage_inst_dmem_ram_3848, MEM_stage_inst_dmem_ram_3849, MEM_stage_inst_dmem_ram_3850, MEM_stage_inst_dmem_ram_3851, MEM_stage_inst_dmem_ram_3852, MEM_stage_inst_dmem_ram_3853, MEM_stage_inst_dmem_ram_3854, MEM_stage_inst_dmem_ram_3855, MEM_stage_inst_dmem_ram_3856, MEM_stage_inst_dmem_ram_3857, MEM_stage_inst_dmem_ram_3858, MEM_stage_inst_dmem_ram_3859, MEM_stage_inst_dmem_ram_3860, MEM_stage_inst_dmem_ram_3861, MEM_stage_inst_dmem_ram_3862, MEM_stage_inst_dmem_ram_3863, MEM_stage_inst_dmem_ram_3864, MEM_stage_inst_dmem_ram_3865, MEM_stage_inst_dmem_ram_3866, MEM_stage_inst_dmem_ram_3867, MEM_stage_inst_dmem_ram_3868, MEM_stage_inst_dmem_ram_3869, MEM_stage_inst_dmem_ram_3870, MEM_stage_inst_dmem_ram_3871, MEM_stage_inst_dmem_ram_3872, MEM_stage_inst_dmem_ram_3873, MEM_stage_inst_dmem_ram_3874, MEM_stage_inst_dmem_ram_3875, MEM_stage_inst_dmem_ram_3876, MEM_stage_inst_dmem_ram_3877, MEM_stage_inst_dmem_ram_3878, MEM_stage_inst_dmem_ram_3879, MEM_stage_inst_dmem_ram_3880, MEM_stage_inst_dmem_ram_3881, MEM_stage_inst_dmem_ram_3882, MEM_stage_inst_dmem_ram_3883, MEM_stage_inst_dmem_ram_3884, MEM_stage_inst_dmem_ram_3885, MEM_stage_inst_dmem_ram_3886, MEM_stage_inst_dmem_ram_3887, MEM_stage_inst_dmem_ram_3888, MEM_stage_inst_dmem_ram_3889, MEM_stage_inst_dmem_ram_3890, MEM_stage_inst_dmem_ram_3891, MEM_stage_inst_dmem_ram_3892, MEM_stage_inst_dmem_ram_3893, MEM_stage_inst_dmem_ram_3894, MEM_stage_inst_dmem_ram_3895, MEM_stage_inst_dmem_ram_3896, MEM_stage_inst_dmem_ram_3897, MEM_stage_inst_dmem_ram_3898, MEM_stage_inst_dmem_ram_3899, MEM_stage_inst_dmem_ram_3900, MEM_stage_inst_dmem_ram_3901, MEM_stage_inst_dmem_ram_3902, MEM_stage_inst_dmem_ram_3903, MEM_stage_inst_dmem_ram_3904, MEM_stage_inst_dmem_ram_3905, MEM_stage_inst_dmem_ram_3906, MEM_stage_inst_dmem_ram_3907, MEM_stage_inst_dmem_ram_3908, MEM_stage_inst_dmem_ram_3909, MEM_stage_inst_dmem_ram_3910, MEM_stage_inst_dmem_ram_3911, MEM_stage_inst_dmem_ram_3912, MEM_stage_inst_dmem_ram_3913, MEM_stage_inst_dmem_ram_3914, MEM_stage_inst_dmem_ram_3915, MEM_stage_inst_dmem_ram_3916, MEM_stage_inst_dmem_ram_3917, MEM_stage_inst_dmem_ram_3918, MEM_stage_inst_dmem_ram_3919, MEM_stage_inst_dmem_ram_3920, MEM_stage_inst_dmem_ram_3921, MEM_stage_inst_dmem_ram_3922, MEM_stage_inst_dmem_ram_3923, MEM_stage_inst_dmem_ram_3924, MEM_stage_inst_dmem_ram_3925, MEM_stage_inst_dmem_ram_3926, MEM_stage_inst_dmem_ram_3927, MEM_stage_inst_dmem_ram_3928, MEM_stage_inst_dmem_ram_3929, MEM_stage_inst_dmem_ram_3930, MEM_stage_inst_dmem_ram_3931, MEM_stage_inst_dmem_ram_3932, MEM_stage_inst_dmem_ram_3933, MEM_stage_inst_dmem_ram_3934, MEM_stage_inst_dmem_ram_3935, MEM_stage_inst_dmem_ram_3936, MEM_stage_inst_dmem_ram_3937, MEM_stage_inst_dmem_ram_3938, MEM_stage_inst_dmem_ram_3939, MEM_stage_inst_dmem_ram_3940, MEM_stage_inst_dmem_ram_3941, MEM_stage_inst_dmem_ram_3942, MEM_stage_inst_dmem_ram_3943, MEM_stage_inst_dmem_ram_3944, MEM_stage_inst_dmem_ram_3945, MEM_stage_inst_dmem_ram_3946, MEM_stage_inst_dmem_ram_3947, MEM_stage_inst_dmem_ram_3948, MEM_stage_inst_dmem_ram_3949, MEM_stage_inst_dmem_ram_3950, MEM_stage_inst_dmem_ram_3951, MEM_stage_inst_dmem_ram_3952, MEM_stage_inst_dmem_ram_3953, MEM_stage_inst_dmem_ram_3954, MEM_stage_inst_dmem_ram_3955, MEM_stage_inst_dmem_ram_3956, MEM_stage_inst_dmem_ram_3957, MEM_stage_inst_dmem_ram_3958, MEM_stage_inst_dmem_ram_3959, MEM_stage_inst_dmem_ram_3960, MEM_stage_inst_dmem_ram_3961, MEM_stage_inst_dmem_ram_3962, MEM_stage_inst_dmem_ram_3963, MEM_stage_inst_dmem_ram_3964, MEM_stage_inst_dmem_ram_3965, MEM_stage_inst_dmem_ram_3966, MEM_stage_inst_dmem_ram_3967, MEM_stage_inst_dmem_ram_3968, MEM_stage_inst_dmem_ram_3969, MEM_stage_inst_dmem_ram_3970, MEM_stage_inst_dmem_ram_3971, MEM_stage_inst_dmem_ram_3972, MEM_stage_inst_dmem_ram_3973, MEM_stage_inst_dmem_ram_3974, MEM_stage_inst_dmem_ram_3975, MEM_stage_inst_dmem_ram_3976, MEM_stage_inst_dmem_ram_3977, MEM_stage_inst_dmem_ram_3978, MEM_stage_inst_dmem_ram_3979, MEM_stage_inst_dmem_ram_3980, MEM_stage_inst_dmem_ram_3981, MEM_stage_inst_dmem_ram_3982, MEM_stage_inst_dmem_ram_3983, MEM_stage_inst_dmem_ram_3984, MEM_stage_inst_dmem_ram_3985, MEM_stage_inst_dmem_ram_3986, MEM_stage_inst_dmem_ram_3987, MEM_stage_inst_dmem_ram_3988, MEM_stage_inst_dmem_ram_3989, MEM_stage_inst_dmem_ram_3990, MEM_stage_inst_dmem_ram_3991, MEM_stage_inst_dmem_ram_3992, MEM_stage_inst_dmem_ram_3993, MEM_stage_inst_dmem_ram_3994, MEM_stage_inst_dmem_ram_3995, MEM_stage_inst_dmem_ram_3996, MEM_stage_inst_dmem_ram_3997, MEM_stage_inst_dmem_ram_3998, MEM_stage_inst_dmem_ram_3999, MEM_stage_inst_dmem_ram_4000, MEM_stage_inst_dmem_ram_4001, MEM_stage_inst_dmem_ram_4002, MEM_stage_inst_dmem_ram_4003, MEM_stage_inst_dmem_ram_4004, MEM_stage_inst_dmem_ram_4005, MEM_stage_inst_dmem_ram_4006, MEM_stage_inst_dmem_ram_4007, MEM_stage_inst_dmem_ram_4008, MEM_stage_inst_dmem_ram_4009, MEM_stage_inst_dmem_ram_4010, MEM_stage_inst_dmem_ram_4011, MEM_stage_inst_dmem_ram_4012, MEM_stage_inst_dmem_ram_4013, MEM_stage_inst_dmem_ram_4014, MEM_stage_inst_dmem_ram_4015, MEM_stage_inst_dmem_ram_4016, MEM_stage_inst_dmem_ram_4017, MEM_stage_inst_dmem_ram_4018, MEM_stage_inst_dmem_ram_4019, MEM_stage_inst_dmem_ram_4020, MEM_stage_inst_dmem_ram_4021, MEM_stage_inst_dmem_ram_4022, MEM_stage_inst_dmem_ram_4023, MEM_stage_inst_dmem_ram_4024, MEM_stage_inst_dmem_ram_4025, MEM_stage_inst_dmem_ram_4026, MEM_stage_inst_dmem_ram_4027, MEM_stage_inst_dmem_ram_4028, MEM_stage_inst_dmem_ram_4029, MEM_stage_inst_dmem_ram_4030, MEM_stage_inst_dmem_ram_4031, MEM_stage_inst_dmem_ram_4032, MEM_stage_inst_dmem_ram_4033, MEM_stage_inst_dmem_ram_4034, MEM_stage_inst_dmem_ram_4035, MEM_stage_inst_dmem_ram_4036, MEM_stage_inst_dmem_ram_4037, MEM_stage_inst_dmem_ram_4038, MEM_stage_inst_dmem_ram_4039, MEM_stage_inst_dmem_ram_4040, MEM_stage_inst_dmem_ram_4041, MEM_stage_inst_dmem_ram_4042, MEM_stage_inst_dmem_ram_4043, MEM_stage_inst_dmem_ram_4044, MEM_stage_inst_dmem_ram_4045, MEM_stage_inst_dmem_ram_4046, MEM_stage_inst_dmem_ram_4047, MEM_stage_inst_dmem_ram_4048, MEM_stage_inst_dmem_ram_4049, MEM_stage_inst_dmem_ram_4050, MEM_stage_inst_dmem_ram_4051, MEM_stage_inst_dmem_ram_4052, MEM_stage_inst_dmem_ram_4053, MEM_stage_inst_dmem_ram_4054, MEM_stage_inst_dmem_ram_4055, MEM_stage_inst_dmem_ram_4056, MEM_stage_inst_dmem_ram_4057, MEM_stage_inst_dmem_ram_4058, MEM_stage_inst_dmem_ram_4059, MEM_stage_inst_dmem_ram_4060, MEM_stage_inst_dmem_ram_4061, MEM_stage_inst_dmem_ram_4062, MEM_stage_inst_dmem_ram_4063, MEM_stage_inst_dmem_ram_4064, MEM_stage_inst_dmem_ram_4065, MEM_stage_inst_dmem_ram_4066, MEM_stage_inst_dmem_ram_4067, MEM_stage_inst_dmem_ram_4068, MEM_stage_inst_dmem_ram_4069, MEM_stage_inst_dmem_ram_4070, MEM_stage_inst_dmem_ram_4071, MEM_stage_inst_dmem_ram_4072, MEM_stage_inst_dmem_ram_4073, MEM_stage_inst_dmem_ram_4074, MEM_stage_inst_dmem_ram_4075, MEM_stage_inst_dmem_ram_4076, MEM_stage_inst_dmem_ram_4077, MEM_stage_inst_dmem_ram_4078, MEM_stage_inst_dmem_ram_4079, MEM_stage_inst_dmem_ram_4080, MEM_stage_inst_dmem_ram_4081, MEM_stage_inst_dmem_ram_4082, MEM_stage_inst_dmem_ram_4083, MEM_stage_inst_dmem_ram_4084, MEM_stage_inst_dmem_ram_4085, MEM_stage_inst_dmem_ram_4086, MEM_stage_inst_dmem_ram_4087, MEM_stage_inst_dmem_ram_4088, MEM_stage_inst_dmem_ram_4089, MEM_stage_inst_dmem_ram_4090, MEM_stage_inst_dmem_ram_4091, MEM_stage_inst_dmem_ram_4092, MEM_stage_inst_dmem_ram_4093, MEM_stage_inst_dmem_ram_4094, MEM_stage_inst_dmem_ram_4095, MEM_stage_inst_dmem_ram_3072, MEM_stage_inst_dmem_ram_3073, MEM_stage_inst_dmem_ram_3074, MEM_stage_inst_dmem_ram_3075, MEM_stage_inst_dmem_ram_3076, MEM_stage_inst_dmem_ram_3077, MEM_stage_inst_dmem_ram_3078, MEM_stage_inst_dmem_ram_3079, MEM_stage_inst_dmem_ram_3080, MEM_stage_inst_dmem_ram_3081, MEM_stage_inst_dmem_ram_3082, MEM_stage_inst_dmem_ram_3083, MEM_stage_inst_dmem_ram_3084, MEM_stage_inst_dmem_ram_3085, MEM_stage_inst_dmem_ram_3086, MEM_stage_inst_dmem_ram_3087, MEM_stage_inst_dmem_ram_3088, MEM_stage_inst_dmem_ram_3089, MEM_stage_inst_dmem_ram_3090, MEM_stage_inst_dmem_ram_3091, MEM_stage_inst_dmem_ram_3092, MEM_stage_inst_dmem_ram_3093, MEM_stage_inst_dmem_ram_3094, MEM_stage_inst_dmem_ram_3095, MEM_stage_inst_dmem_ram_3096, MEM_stage_inst_dmem_ram_3097, MEM_stage_inst_dmem_ram_3098, MEM_stage_inst_dmem_ram_3099, MEM_stage_inst_dmem_ram_3100, MEM_stage_inst_dmem_ram_3101, MEM_stage_inst_dmem_ram_3102, MEM_stage_inst_dmem_ram_3103, MEM_stage_inst_dmem_ram_3104, MEM_stage_inst_dmem_ram_3105, MEM_stage_inst_dmem_ram_3106, MEM_stage_inst_dmem_ram_3107, MEM_stage_inst_dmem_ram_3108, MEM_stage_inst_dmem_ram_3109, MEM_stage_inst_dmem_ram_3110, MEM_stage_inst_dmem_ram_3111, MEM_stage_inst_dmem_ram_3112, MEM_stage_inst_dmem_ram_3113, MEM_stage_inst_dmem_ram_3114, MEM_stage_inst_dmem_ram_3115, MEM_stage_inst_dmem_ram_3116, MEM_stage_inst_dmem_ram_3117, MEM_stage_inst_dmem_ram_3118, MEM_stage_inst_dmem_ram_3119, MEM_stage_inst_dmem_ram_3120, MEM_stage_inst_dmem_ram_3121, MEM_stage_inst_dmem_ram_3122, MEM_stage_inst_dmem_ram_3123, MEM_stage_inst_dmem_ram_3124, MEM_stage_inst_dmem_ram_3125, MEM_stage_inst_dmem_ram_3126, MEM_stage_inst_dmem_ram_3127, MEM_stage_inst_dmem_ram_3128, MEM_stage_inst_dmem_ram_3129, MEM_stage_inst_dmem_ram_3130, MEM_stage_inst_dmem_ram_3131, MEM_stage_inst_dmem_ram_3132, MEM_stage_inst_dmem_ram_3133, MEM_stage_inst_dmem_ram_3134, MEM_stage_inst_dmem_ram_3135, MEM_stage_inst_dmem_ram_3136, MEM_stage_inst_dmem_ram_3137, MEM_stage_inst_dmem_ram_3138, MEM_stage_inst_dmem_ram_3139, MEM_stage_inst_dmem_ram_3140, MEM_stage_inst_dmem_ram_3141, MEM_stage_inst_dmem_ram_3142, MEM_stage_inst_dmem_ram_3143, MEM_stage_inst_dmem_ram_3144, MEM_stage_inst_dmem_ram_3145, MEM_stage_inst_dmem_ram_3146, MEM_stage_inst_dmem_ram_3147, MEM_stage_inst_dmem_ram_3148, MEM_stage_inst_dmem_ram_3149, MEM_stage_inst_dmem_ram_3150, MEM_stage_inst_dmem_ram_3151, MEM_stage_inst_dmem_ram_3152, MEM_stage_inst_dmem_ram_3153, MEM_stage_inst_dmem_ram_3154, MEM_stage_inst_dmem_ram_3155, MEM_stage_inst_dmem_ram_3156, MEM_stage_inst_dmem_ram_3157, MEM_stage_inst_dmem_ram_3158, MEM_stage_inst_dmem_ram_3159, MEM_stage_inst_dmem_ram_3160, MEM_stage_inst_dmem_ram_3161, MEM_stage_inst_dmem_ram_3162, MEM_stage_inst_dmem_ram_3163, MEM_stage_inst_dmem_ram_3164, MEM_stage_inst_dmem_ram_3165, MEM_stage_inst_dmem_ram_3166, MEM_stage_inst_dmem_ram_3167, MEM_stage_inst_dmem_ram_3168, MEM_stage_inst_dmem_ram_3169, MEM_stage_inst_dmem_ram_3170, MEM_stage_inst_dmem_ram_3171, MEM_stage_inst_dmem_ram_3172, MEM_stage_inst_dmem_ram_3173, MEM_stage_inst_dmem_ram_3174, MEM_stage_inst_dmem_ram_3175, MEM_stage_inst_dmem_ram_3176, MEM_stage_inst_dmem_ram_3177, MEM_stage_inst_dmem_ram_3178, MEM_stage_inst_dmem_ram_3179, MEM_stage_inst_dmem_ram_3180, MEM_stage_inst_dmem_ram_3181, MEM_stage_inst_dmem_ram_3182, MEM_stage_inst_dmem_ram_3183, MEM_stage_inst_dmem_ram_3184, MEM_stage_inst_dmem_ram_3185, MEM_stage_inst_dmem_ram_3186, MEM_stage_inst_dmem_ram_3187, MEM_stage_inst_dmem_ram_3188, MEM_stage_inst_dmem_ram_3189, MEM_stage_inst_dmem_ram_3190, MEM_stage_inst_dmem_ram_3191, MEM_stage_inst_dmem_ram_3192, MEM_stage_inst_dmem_ram_3193, MEM_stage_inst_dmem_ram_3194, MEM_stage_inst_dmem_ram_3195, MEM_stage_inst_dmem_ram_3196, MEM_stage_inst_dmem_ram_3197, MEM_stage_inst_dmem_ram_3198, MEM_stage_inst_dmem_ram_3199, MEM_stage_inst_dmem_ram_3200, MEM_stage_inst_dmem_ram_3201, MEM_stage_inst_dmem_ram_3202, MEM_stage_inst_dmem_ram_3203, MEM_stage_inst_dmem_ram_3204, MEM_stage_inst_dmem_ram_3205, MEM_stage_inst_dmem_ram_3206, MEM_stage_inst_dmem_ram_3207, MEM_stage_inst_dmem_ram_3208, MEM_stage_inst_dmem_ram_3209, MEM_stage_inst_dmem_ram_3210, MEM_stage_inst_dmem_ram_3211, MEM_stage_inst_dmem_ram_3212, MEM_stage_inst_dmem_ram_3213, MEM_stage_inst_dmem_ram_3214, MEM_stage_inst_dmem_ram_3215, MEM_stage_inst_dmem_ram_3216, MEM_stage_inst_dmem_ram_3217, MEM_stage_inst_dmem_ram_3218, MEM_stage_inst_dmem_ram_3219, MEM_stage_inst_dmem_ram_3220, MEM_stage_inst_dmem_ram_3221, MEM_stage_inst_dmem_ram_3222, MEM_stage_inst_dmem_ram_3223, MEM_stage_inst_dmem_ram_3224, MEM_stage_inst_dmem_ram_3225, MEM_stage_inst_dmem_ram_3226, MEM_stage_inst_dmem_ram_3227, MEM_stage_inst_dmem_ram_3228, MEM_stage_inst_dmem_ram_3229, MEM_stage_inst_dmem_ram_3230, MEM_stage_inst_dmem_ram_3231, MEM_stage_inst_dmem_ram_3232, MEM_stage_inst_dmem_ram_3233, MEM_stage_inst_dmem_ram_3234, MEM_stage_inst_dmem_ram_3235, MEM_stage_inst_dmem_ram_3236, MEM_stage_inst_dmem_ram_3237, MEM_stage_inst_dmem_ram_3238, MEM_stage_inst_dmem_ram_3239, MEM_stage_inst_dmem_ram_3240, MEM_stage_inst_dmem_ram_3241, MEM_stage_inst_dmem_ram_3242, MEM_stage_inst_dmem_ram_3243, MEM_stage_inst_dmem_ram_3244, MEM_stage_inst_dmem_ram_3245, MEM_stage_inst_dmem_ram_3246, MEM_stage_inst_dmem_ram_3247, MEM_stage_inst_dmem_ram_3248, MEM_stage_inst_dmem_ram_3249, MEM_stage_inst_dmem_ram_3250, MEM_stage_inst_dmem_ram_3251, MEM_stage_inst_dmem_ram_3252, MEM_stage_inst_dmem_ram_3253, MEM_stage_inst_dmem_ram_3254, MEM_stage_inst_dmem_ram_3255, MEM_stage_inst_dmem_ram_3256, MEM_stage_inst_dmem_ram_3257, MEM_stage_inst_dmem_ram_3258, MEM_stage_inst_dmem_ram_3259, MEM_stage_inst_dmem_ram_3260, MEM_stage_inst_dmem_ram_3261, MEM_stage_inst_dmem_ram_3262, MEM_stage_inst_dmem_ram_3263, MEM_stage_inst_dmem_ram_3264, MEM_stage_inst_dmem_ram_3265, MEM_stage_inst_dmem_ram_3266, MEM_stage_inst_dmem_ram_3267, MEM_stage_inst_dmem_ram_3268, MEM_stage_inst_dmem_ram_3269, MEM_stage_inst_dmem_ram_3270, MEM_stage_inst_dmem_ram_3271, MEM_stage_inst_dmem_ram_3272, MEM_stage_inst_dmem_ram_3273, MEM_stage_inst_dmem_ram_3274, MEM_stage_inst_dmem_ram_3275, MEM_stage_inst_dmem_ram_3276, MEM_stage_inst_dmem_ram_3277, MEM_stage_inst_dmem_ram_3278, MEM_stage_inst_dmem_ram_3279, MEM_stage_inst_dmem_ram_3280, MEM_stage_inst_dmem_ram_3281, MEM_stage_inst_dmem_ram_3282, MEM_stage_inst_dmem_ram_3283, MEM_stage_inst_dmem_ram_3284, MEM_stage_inst_dmem_ram_3285, MEM_stage_inst_dmem_ram_3286, MEM_stage_inst_dmem_ram_3287, MEM_stage_inst_dmem_ram_3288, MEM_stage_inst_dmem_ram_3289, MEM_stage_inst_dmem_ram_3290, MEM_stage_inst_dmem_ram_3291, MEM_stage_inst_dmem_ram_3292, MEM_stage_inst_dmem_ram_3293, MEM_stage_inst_dmem_ram_3294, MEM_stage_inst_dmem_ram_3295, MEM_stage_inst_dmem_ram_3296, MEM_stage_inst_dmem_ram_3297, MEM_stage_inst_dmem_ram_3298, MEM_stage_inst_dmem_ram_3299, MEM_stage_inst_dmem_ram_3300, MEM_stage_inst_dmem_ram_3301, MEM_stage_inst_dmem_ram_3302, MEM_stage_inst_dmem_ram_3303, MEM_stage_inst_dmem_ram_3304, MEM_stage_inst_dmem_ram_3305, MEM_stage_inst_dmem_ram_3306, MEM_stage_inst_dmem_ram_3307, MEM_stage_inst_dmem_ram_3308, MEM_stage_inst_dmem_ram_3309, MEM_stage_inst_dmem_ram_3310, MEM_stage_inst_dmem_ram_3311, MEM_stage_inst_dmem_ram_3312, MEM_stage_inst_dmem_ram_3313, MEM_stage_inst_dmem_ram_3314, MEM_stage_inst_dmem_ram_3315, MEM_stage_inst_dmem_ram_3316, MEM_stage_inst_dmem_ram_3317, MEM_stage_inst_dmem_ram_3318, MEM_stage_inst_dmem_ram_3319, MEM_stage_inst_dmem_ram_3320, MEM_stage_inst_dmem_ram_3321, MEM_stage_inst_dmem_ram_3322, MEM_stage_inst_dmem_ram_3323, MEM_stage_inst_dmem_ram_3324, MEM_stage_inst_dmem_ram_3325, MEM_stage_inst_dmem_ram_3326, MEM_stage_inst_dmem_ram_3327, MEM_stage_inst_dmem_ram_3328, MEM_stage_inst_dmem_ram_3329, MEM_stage_inst_dmem_ram_3330, MEM_stage_inst_dmem_ram_3331, MEM_stage_inst_dmem_ram_3332, MEM_stage_inst_dmem_ram_3333, MEM_stage_inst_dmem_ram_3334, MEM_stage_inst_dmem_ram_3335, MEM_stage_inst_dmem_ram_3336, MEM_stage_inst_dmem_ram_3337, MEM_stage_inst_dmem_ram_3338, MEM_stage_inst_dmem_ram_3339, MEM_stage_inst_dmem_ram_3340, MEM_stage_inst_dmem_ram_3341, MEM_stage_inst_dmem_ram_3342, MEM_stage_inst_dmem_ram_3343, MEM_stage_inst_dmem_ram_3344, MEM_stage_inst_dmem_ram_3345, MEM_stage_inst_dmem_ram_3346, MEM_stage_inst_dmem_ram_3347, MEM_stage_inst_dmem_ram_3348, MEM_stage_inst_dmem_ram_3349, MEM_stage_inst_dmem_ram_3350, MEM_stage_inst_dmem_ram_3351, MEM_stage_inst_dmem_ram_3352, MEM_stage_inst_dmem_ram_3353, MEM_stage_inst_dmem_ram_3354, MEM_stage_inst_dmem_ram_3355, MEM_stage_inst_dmem_ram_3356, MEM_stage_inst_dmem_ram_3357, MEM_stage_inst_dmem_ram_3358, MEM_stage_inst_dmem_ram_3359, MEM_stage_inst_dmem_ram_3360, MEM_stage_inst_dmem_ram_3361, MEM_stage_inst_dmem_ram_3362, MEM_stage_inst_dmem_ram_3363, MEM_stage_inst_dmem_ram_3364, MEM_stage_inst_dmem_ram_3365, MEM_stage_inst_dmem_ram_3366, MEM_stage_inst_dmem_ram_3367, MEM_stage_inst_dmem_ram_3368, MEM_stage_inst_dmem_ram_3369, MEM_stage_inst_dmem_ram_3370, MEM_stage_inst_dmem_ram_3371, MEM_stage_inst_dmem_ram_3372, MEM_stage_inst_dmem_ram_3373, MEM_stage_inst_dmem_ram_3374, MEM_stage_inst_dmem_ram_3375, MEM_stage_inst_dmem_ram_3376, MEM_stage_inst_dmem_ram_3377, MEM_stage_inst_dmem_ram_3378, MEM_stage_inst_dmem_ram_3379, MEM_stage_inst_dmem_ram_3380, MEM_stage_inst_dmem_ram_3381, MEM_stage_inst_dmem_ram_3382, MEM_stage_inst_dmem_ram_3383, MEM_stage_inst_dmem_ram_3384, MEM_stage_inst_dmem_ram_3385, MEM_stage_inst_dmem_ram_3386, MEM_stage_inst_dmem_ram_3387, MEM_stage_inst_dmem_ram_3388, MEM_stage_inst_dmem_ram_3389, MEM_stage_inst_dmem_ram_3390, MEM_stage_inst_dmem_ram_3391, MEM_stage_inst_dmem_ram_3392, MEM_stage_inst_dmem_ram_3393, MEM_stage_inst_dmem_ram_3394, MEM_stage_inst_dmem_ram_3395, MEM_stage_inst_dmem_ram_3396, MEM_stage_inst_dmem_ram_3397, MEM_stage_inst_dmem_ram_3398, MEM_stage_inst_dmem_ram_3399, MEM_stage_inst_dmem_ram_3400, MEM_stage_inst_dmem_ram_3401, MEM_stage_inst_dmem_ram_3402, MEM_stage_inst_dmem_ram_3403, MEM_stage_inst_dmem_ram_3404, MEM_stage_inst_dmem_ram_3405, MEM_stage_inst_dmem_ram_3406, MEM_stage_inst_dmem_ram_3407, MEM_stage_inst_dmem_ram_3408, MEM_stage_inst_dmem_ram_3409, MEM_stage_inst_dmem_ram_3410, MEM_stage_inst_dmem_ram_3411, MEM_stage_inst_dmem_ram_3412, MEM_stage_inst_dmem_ram_3413, MEM_stage_inst_dmem_ram_3414, MEM_stage_inst_dmem_ram_3415, MEM_stage_inst_dmem_ram_3416, MEM_stage_inst_dmem_ram_3417, MEM_stage_inst_dmem_ram_3418, MEM_stage_inst_dmem_ram_3419, MEM_stage_inst_dmem_ram_3420, MEM_stage_inst_dmem_ram_3421, MEM_stage_inst_dmem_ram_3422, MEM_stage_inst_dmem_ram_3423, MEM_stage_inst_dmem_ram_3424, MEM_stage_inst_dmem_ram_3425, MEM_stage_inst_dmem_ram_3426, MEM_stage_inst_dmem_ram_3427, MEM_stage_inst_dmem_ram_3428, MEM_stage_inst_dmem_ram_3429, MEM_stage_inst_dmem_ram_3430, MEM_stage_inst_dmem_ram_3431, MEM_stage_inst_dmem_ram_3432, MEM_stage_inst_dmem_ram_3433, MEM_stage_inst_dmem_ram_3434, MEM_stage_inst_dmem_ram_3435, MEM_stage_inst_dmem_ram_3436, MEM_stage_inst_dmem_ram_3437, MEM_stage_inst_dmem_ram_3438, MEM_stage_inst_dmem_ram_3439, MEM_stage_inst_dmem_ram_3440, MEM_stage_inst_dmem_ram_3441, MEM_stage_inst_dmem_ram_3442, MEM_stage_inst_dmem_ram_3443, MEM_stage_inst_dmem_ram_3444, MEM_stage_inst_dmem_ram_3445, MEM_stage_inst_dmem_ram_3446, MEM_stage_inst_dmem_ram_3447, MEM_stage_inst_dmem_ram_3448, MEM_stage_inst_dmem_ram_3449, MEM_stage_inst_dmem_ram_3450, MEM_stage_inst_dmem_ram_3451, MEM_stage_inst_dmem_ram_3452, MEM_stage_inst_dmem_ram_3453, MEM_stage_inst_dmem_ram_3454, MEM_stage_inst_dmem_ram_3455, MEM_stage_inst_dmem_ram_3456, MEM_stage_inst_dmem_ram_3457, MEM_stage_inst_dmem_ram_3458, MEM_stage_inst_dmem_ram_3459, MEM_stage_inst_dmem_ram_3460, MEM_stage_inst_dmem_ram_3461, MEM_stage_inst_dmem_ram_3462, MEM_stage_inst_dmem_ram_3463, MEM_stage_inst_dmem_ram_3464, MEM_stage_inst_dmem_ram_3465, MEM_stage_inst_dmem_ram_3466, MEM_stage_inst_dmem_ram_3467, MEM_stage_inst_dmem_ram_3468, MEM_stage_inst_dmem_ram_3469, MEM_stage_inst_dmem_ram_3470, MEM_stage_inst_dmem_ram_3471, MEM_stage_inst_dmem_ram_3472, MEM_stage_inst_dmem_ram_3473, MEM_stage_inst_dmem_ram_3474, MEM_stage_inst_dmem_ram_3475, MEM_stage_inst_dmem_ram_3476, MEM_stage_inst_dmem_ram_3477, MEM_stage_inst_dmem_ram_3478, MEM_stage_inst_dmem_ram_3479, MEM_stage_inst_dmem_ram_3480, MEM_stage_inst_dmem_ram_3481, MEM_stage_inst_dmem_ram_3482, MEM_stage_inst_dmem_ram_3483, MEM_stage_inst_dmem_ram_3484, MEM_stage_inst_dmem_ram_3485, MEM_stage_inst_dmem_ram_3486, MEM_stage_inst_dmem_ram_3487, MEM_stage_inst_dmem_ram_3488, MEM_stage_inst_dmem_ram_3489, MEM_stage_inst_dmem_ram_3490, MEM_stage_inst_dmem_ram_3491, MEM_stage_inst_dmem_ram_3492, MEM_stage_inst_dmem_ram_3493, MEM_stage_inst_dmem_ram_3494, MEM_stage_inst_dmem_ram_3495, MEM_stage_inst_dmem_ram_3496, MEM_stage_inst_dmem_ram_3497, MEM_stage_inst_dmem_ram_3498, MEM_stage_inst_dmem_ram_3499, MEM_stage_inst_dmem_ram_3500, MEM_stage_inst_dmem_ram_3501, MEM_stage_inst_dmem_ram_3502, MEM_stage_inst_dmem_ram_3503, MEM_stage_inst_dmem_ram_3504, MEM_stage_inst_dmem_ram_3505, MEM_stage_inst_dmem_ram_3506, MEM_stage_inst_dmem_ram_3507, MEM_stage_inst_dmem_ram_3508, MEM_stage_inst_dmem_ram_3509, MEM_stage_inst_dmem_ram_3510, MEM_stage_inst_dmem_ram_3511, MEM_stage_inst_dmem_ram_3512, MEM_stage_inst_dmem_ram_3513, MEM_stage_inst_dmem_ram_3514, MEM_stage_inst_dmem_ram_3515, MEM_stage_inst_dmem_ram_3516, MEM_stage_inst_dmem_ram_3517, MEM_stage_inst_dmem_ram_3518, MEM_stage_inst_dmem_ram_3519, MEM_stage_inst_dmem_ram_3520, MEM_stage_inst_dmem_ram_3521, MEM_stage_inst_dmem_ram_3522, MEM_stage_inst_dmem_ram_3523, MEM_stage_inst_dmem_ram_3524, MEM_stage_inst_dmem_ram_3525, MEM_stage_inst_dmem_ram_3526, MEM_stage_inst_dmem_ram_3527, MEM_stage_inst_dmem_ram_3528, MEM_stage_inst_dmem_ram_3529, MEM_stage_inst_dmem_ram_3530, MEM_stage_inst_dmem_ram_3531, MEM_stage_inst_dmem_ram_3532, MEM_stage_inst_dmem_ram_3533, MEM_stage_inst_dmem_ram_3534, MEM_stage_inst_dmem_ram_3535, MEM_stage_inst_dmem_ram_3536, MEM_stage_inst_dmem_ram_3537, MEM_stage_inst_dmem_ram_3538, MEM_stage_inst_dmem_ram_3539, MEM_stage_inst_dmem_ram_3540, MEM_stage_inst_dmem_ram_3541, MEM_stage_inst_dmem_ram_3542, MEM_stage_inst_dmem_ram_3543, MEM_stage_inst_dmem_ram_3544, MEM_stage_inst_dmem_ram_3545, MEM_stage_inst_dmem_ram_3546, MEM_stage_inst_dmem_ram_3547, MEM_stage_inst_dmem_ram_3548, MEM_stage_inst_dmem_ram_3549, MEM_stage_inst_dmem_ram_3550, MEM_stage_inst_dmem_ram_3551, MEM_stage_inst_dmem_ram_3552, MEM_stage_inst_dmem_ram_3553, MEM_stage_inst_dmem_ram_3554, MEM_stage_inst_dmem_ram_3555, MEM_stage_inst_dmem_ram_3556, MEM_stage_inst_dmem_ram_3557, MEM_stage_inst_dmem_ram_3558, MEM_stage_inst_dmem_ram_3559, MEM_stage_inst_dmem_ram_3560, MEM_stage_inst_dmem_ram_3561, MEM_stage_inst_dmem_ram_3562, MEM_stage_inst_dmem_ram_3563, MEM_stage_inst_dmem_ram_3564, MEM_stage_inst_dmem_ram_3565, MEM_stage_inst_dmem_ram_3566, MEM_stage_inst_dmem_ram_3567, MEM_stage_inst_dmem_ram_3568, MEM_stage_inst_dmem_ram_3569, MEM_stage_inst_dmem_ram_3570, MEM_stage_inst_dmem_ram_3571, MEM_stage_inst_dmem_ram_3572, MEM_stage_inst_dmem_ram_3573, MEM_stage_inst_dmem_ram_3574, MEM_stage_inst_dmem_ram_3575, MEM_stage_inst_dmem_ram_3576, MEM_stage_inst_dmem_ram_3577, MEM_stage_inst_dmem_ram_3578, MEM_stage_inst_dmem_ram_3579, MEM_stage_inst_dmem_ram_3580, MEM_stage_inst_dmem_ram_3581, MEM_stage_inst_dmem_ram_3582, MEM_stage_inst_dmem_ram_3583, MEM_stage_inst_dmem_ram_2560, MEM_stage_inst_dmem_ram_2561, MEM_stage_inst_dmem_ram_2562, MEM_stage_inst_dmem_ram_2563, MEM_stage_inst_dmem_ram_2564, MEM_stage_inst_dmem_ram_2565, MEM_stage_inst_dmem_ram_2566, MEM_stage_inst_dmem_ram_2567, MEM_stage_inst_dmem_ram_2568, MEM_stage_inst_dmem_ram_2569, MEM_stage_inst_dmem_ram_2570, MEM_stage_inst_dmem_ram_2571, MEM_stage_inst_dmem_ram_2572, MEM_stage_inst_dmem_ram_2573, MEM_stage_inst_dmem_ram_2574, MEM_stage_inst_dmem_ram_2575, MEM_stage_inst_dmem_ram_2576, MEM_stage_inst_dmem_ram_2577, MEM_stage_inst_dmem_ram_2578, MEM_stage_inst_dmem_ram_2579, MEM_stage_inst_dmem_ram_2580, MEM_stage_inst_dmem_ram_2581, MEM_stage_inst_dmem_ram_2582, MEM_stage_inst_dmem_ram_2583, MEM_stage_inst_dmem_ram_2584, MEM_stage_inst_dmem_ram_2585, MEM_stage_inst_dmem_ram_2586, MEM_stage_inst_dmem_ram_2587, MEM_stage_inst_dmem_ram_2588, MEM_stage_inst_dmem_ram_2589, MEM_stage_inst_dmem_ram_2590, MEM_stage_inst_dmem_ram_2591, MEM_stage_inst_dmem_ram_2592, MEM_stage_inst_dmem_ram_2593, MEM_stage_inst_dmem_ram_2594, MEM_stage_inst_dmem_ram_2595, MEM_stage_inst_dmem_ram_2596, MEM_stage_inst_dmem_ram_2597, MEM_stage_inst_dmem_ram_2598, MEM_stage_inst_dmem_ram_2599, MEM_stage_inst_dmem_ram_2600, MEM_stage_inst_dmem_ram_2601, MEM_stage_inst_dmem_ram_2602, MEM_stage_inst_dmem_ram_2603, MEM_stage_inst_dmem_ram_2604, MEM_stage_inst_dmem_ram_2605, MEM_stage_inst_dmem_ram_2606, MEM_stage_inst_dmem_ram_2607, MEM_stage_inst_dmem_ram_2608, MEM_stage_inst_dmem_ram_2609, MEM_stage_inst_dmem_ram_2610, MEM_stage_inst_dmem_ram_2611, MEM_stage_inst_dmem_ram_2612, MEM_stage_inst_dmem_ram_2613, MEM_stage_inst_dmem_ram_2614, MEM_stage_inst_dmem_ram_2615, MEM_stage_inst_dmem_ram_2616, MEM_stage_inst_dmem_ram_2617, MEM_stage_inst_dmem_ram_2618, MEM_stage_inst_dmem_ram_2619, MEM_stage_inst_dmem_ram_2620, MEM_stage_inst_dmem_ram_2621, MEM_stage_inst_dmem_ram_2622, MEM_stage_inst_dmem_ram_2623, MEM_stage_inst_dmem_ram_2624, MEM_stage_inst_dmem_ram_2625, MEM_stage_inst_dmem_ram_2626, MEM_stage_inst_dmem_ram_2627, MEM_stage_inst_dmem_ram_2628, MEM_stage_inst_dmem_ram_2629, MEM_stage_inst_dmem_ram_2630, MEM_stage_inst_dmem_ram_2631, MEM_stage_inst_dmem_ram_2632, MEM_stage_inst_dmem_ram_2633, MEM_stage_inst_dmem_ram_2634, MEM_stage_inst_dmem_ram_2635, MEM_stage_inst_dmem_ram_2636, MEM_stage_inst_dmem_ram_2637, MEM_stage_inst_dmem_ram_2638, MEM_stage_inst_dmem_ram_2639, MEM_stage_inst_dmem_ram_2640, MEM_stage_inst_dmem_ram_2641, MEM_stage_inst_dmem_ram_2642, MEM_stage_inst_dmem_ram_2643, MEM_stage_inst_dmem_ram_2644, MEM_stage_inst_dmem_ram_2645, MEM_stage_inst_dmem_ram_2646, MEM_stage_inst_dmem_ram_2647, MEM_stage_inst_dmem_ram_2648, MEM_stage_inst_dmem_ram_2649, MEM_stage_inst_dmem_ram_2650, MEM_stage_inst_dmem_ram_2651, MEM_stage_inst_dmem_ram_2652, MEM_stage_inst_dmem_ram_2653, MEM_stage_inst_dmem_ram_2654, MEM_stage_inst_dmem_ram_2655, MEM_stage_inst_dmem_ram_2656, MEM_stage_inst_dmem_ram_2657, MEM_stage_inst_dmem_ram_2658, MEM_stage_inst_dmem_ram_2659, MEM_stage_inst_dmem_ram_2660, MEM_stage_inst_dmem_ram_2661, MEM_stage_inst_dmem_ram_2662, MEM_stage_inst_dmem_ram_2663, MEM_stage_inst_dmem_ram_2664, MEM_stage_inst_dmem_ram_2665, MEM_stage_inst_dmem_ram_2666, MEM_stage_inst_dmem_ram_2667, MEM_stage_inst_dmem_ram_2668, MEM_stage_inst_dmem_ram_2669, MEM_stage_inst_dmem_ram_2670, MEM_stage_inst_dmem_ram_2671, MEM_stage_inst_dmem_ram_2672, MEM_stage_inst_dmem_ram_2673, MEM_stage_inst_dmem_ram_2674, MEM_stage_inst_dmem_ram_2675, MEM_stage_inst_dmem_ram_2676, MEM_stage_inst_dmem_ram_2677, MEM_stage_inst_dmem_ram_2678, MEM_stage_inst_dmem_ram_2679, MEM_stage_inst_dmem_ram_2680, MEM_stage_inst_dmem_ram_2681, MEM_stage_inst_dmem_ram_2682, MEM_stage_inst_dmem_ram_2683, MEM_stage_inst_dmem_ram_2684, MEM_stage_inst_dmem_ram_2685, MEM_stage_inst_dmem_ram_2686, MEM_stage_inst_dmem_ram_2687, MEM_stage_inst_dmem_ram_2688, MEM_stage_inst_dmem_ram_2689, MEM_stage_inst_dmem_ram_2690, MEM_stage_inst_dmem_ram_2691, MEM_stage_inst_dmem_ram_2692, MEM_stage_inst_dmem_ram_2693, MEM_stage_inst_dmem_ram_2694, MEM_stage_inst_dmem_ram_2695, MEM_stage_inst_dmem_ram_2696, MEM_stage_inst_dmem_ram_2697, MEM_stage_inst_dmem_ram_2698, MEM_stage_inst_dmem_ram_2699, MEM_stage_inst_dmem_ram_2700, MEM_stage_inst_dmem_ram_2701, MEM_stage_inst_dmem_ram_2702, MEM_stage_inst_dmem_ram_2703, MEM_stage_inst_dmem_ram_2704, MEM_stage_inst_dmem_ram_2705, MEM_stage_inst_dmem_ram_2706, MEM_stage_inst_dmem_ram_2707, MEM_stage_inst_dmem_ram_2708, MEM_stage_inst_dmem_ram_2709, MEM_stage_inst_dmem_ram_2710, MEM_stage_inst_dmem_ram_2711, MEM_stage_inst_dmem_ram_2712, MEM_stage_inst_dmem_ram_2713, MEM_stage_inst_dmem_ram_2714, MEM_stage_inst_dmem_ram_2715, MEM_stage_inst_dmem_ram_2716, MEM_stage_inst_dmem_ram_2717, MEM_stage_inst_dmem_ram_2718, MEM_stage_inst_dmem_ram_2719, MEM_stage_inst_dmem_ram_2720, MEM_stage_inst_dmem_ram_2721, MEM_stage_inst_dmem_ram_2722, MEM_stage_inst_dmem_ram_2723, MEM_stage_inst_dmem_ram_2724, MEM_stage_inst_dmem_ram_2725, MEM_stage_inst_dmem_ram_2726, MEM_stage_inst_dmem_ram_2727, MEM_stage_inst_dmem_ram_2728, MEM_stage_inst_dmem_ram_2729, MEM_stage_inst_dmem_ram_2730, MEM_stage_inst_dmem_ram_2731, MEM_stage_inst_dmem_ram_2732, MEM_stage_inst_dmem_ram_2733, MEM_stage_inst_dmem_ram_2734, MEM_stage_inst_dmem_ram_2735, MEM_stage_inst_dmem_ram_2736, MEM_stage_inst_dmem_ram_2737, MEM_stage_inst_dmem_ram_2738, MEM_stage_inst_dmem_ram_2739, MEM_stage_inst_dmem_ram_2740, MEM_stage_inst_dmem_ram_2741, MEM_stage_inst_dmem_ram_2742, MEM_stage_inst_dmem_ram_2743, MEM_stage_inst_dmem_ram_2744, MEM_stage_inst_dmem_ram_2745, MEM_stage_inst_dmem_ram_2746, MEM_stage_inst_dmem_ram_2747, MEM_stage_inst_dmem_ram_2748, MEM_stage_inst_dmem_ram_2749, MEM_stage_inst_dmem_ram_2750, MEM_stage_inst_dmem_ram_2751, MEM_stage_inst_dmem_ram_2752, MEM_stage_inst_dmem_ram_2753, MEM_stage_inst_dmem_ram_2754, MEM_stage_inst_dmem_ram_2755, MEM_stage_inst_dmem_ram_2756, MEM_stage_inst_dmem_ram_2757, MEM_stage_inst_dmem_ram_2758, MEM_stage_inst_dmem_ram_2759, MEM_stage_inst_dmem_ram_2760, MEM_stage_inst_dmem_ram_2761, MEM_stage_inst_dmem_ram_2762, MEM_stage_inst_dmem_ram_2763, MEM_stage_inst_dmem_ram_2764, MEM_stage_inst_dmem_ram_2765, MEM_stage_inst_dmem_ram_2766, MEM_stage_inst_dmem_ram_2767, MEM_stage_inst_dmem_ram_2768, MEM_stage_inst_dmem_ram_2769, MEM_stage_inst_dmem_ram_2770, MEM_stage_inst_dmem_ram_2771, MEM_stage_inst_dmem_ram_2772, MEM_stage_inst_dmem_ram_2773, MEM_stage_inst_dmem_ram_2774, MEM_stage_inst_dmem_ram_2775, MEM_stage_inst_dmem_ram_2776, MEM_stage_inst_dmem_ram_2777, MEM_stage_inst_dmem_ram_2778, MEM_stage_inst_dmem_ram_2779, MEM_stage_inst_dmem_ram_2780, MEM_stage_inst_dmem_ram_2781, MEM_stage_inst_dmem_ram_2782, MEM_stage_inst_dmem_ram_2783, MEM_stage_inst_dmem_ram_2784, MEM_stage_inst_dmem_ram_2785, MEM_stage_inst_dmem_ram_2786, MEM_stage_inst_dmem_ram_2787, MEM_stage_inst_dmem_ram_2788, MEM_stage_inst_dmem_ram_2789, MEM_stage_inst_dmem_ram_2790, MEM_stage_inst_dmem_ram_2791, MEM_stage_inst_dmem_ram_2792, MEM_stage_inst_dmem_ram_2793, MEM_stage_inst_dmem_ram_2794, MEM_stage_inst_dmem_ram_2795, MEM_stage_inst_dmem_ram_2796, MEM_stage_inst_dmem_ram_2797, MEM_stage_inst_dmem_ram_2798, MEM_stage_inst_dmem_ram_2799, MEM_stage_inst_dmem_ram_2800, MEM_stage_inst_dmem_ram_2801, MEM_stage_inst_dmem_ram_2802, MEM_stage_inst_dmem_ram_2803, MEM_stage_inst_dmem_ram_2804, MEM_stage_inst_dmem_ram_2805, MEM_stage_inst_dmem_ram_2806, MEM_stage_inst_dmem_ram_2807, MEM_stage_inst_dmem_ram_2808, MEM_stage_inst_dmem_ram_2809, MEM_stage_inst_dmem_ram_2810, MEM_stage_inst_dmem_ram_2811, MEM_stage_inst_dmem_ram_2812, MEM_stage_inst_dmem_ram_2813, MEM_stage_inst_dmem_ram_2814, MEM_stage_inst_dmem_ram_2815, MEM_stage_inst_dmem_ram_2816, MEM_stage_inst_dmem_ram_2817, MEM_stage_inst_dmem_ram_2818, MEM_stage_inst_dmem_ram_2819, MEM_stage_inst_dmem_ram_2820, MEM_stage_inst_dmem_ram_2821, MEM_stage_inst_dmem_ram_2822, MEM_stage_inst_dmem_ram_2823, MEM_stage_inst_dmem_ram_2824, MEM_stage_inst_dmem_ram_2825, MEM_stage_inst_dmem_ram_2826, MEM_stage_inst_dmem_ram_2827, MEM_stage_inst_dmem_ram_2828, MEM_stage_inst_dmem_ram_2829, MEM_stage_inst_dmem_ram_2830, MEM_stage_inst_dmem_ram_2831, MEM_stage_inst_dmem_ram_2832, MEM_stage_inst_dmem_ram_2833, MEM_stage_inst_dmem_ram_2834, MEM_stage_inst_dmem_ram_2835, MEM_stage_inst_dmem_ram_2836, MEM_stage_inst_dmem_ram_2837, MEM_stage_inst_dmem_ram_2838, MEM_stage_inst_dmem_ram_2839, MEM_stage_inst_dmem_ram_2840, MEM_stage_inst_dmem_ram_2841, MEM_stage_inst_dmem_ram_2842, MEM_stage_inst_dmem_ram_2843, MEM_stage_inst_dmem_ram_2844, MEM_stage_inst_dmem_ram_2845, MEM_stage_inst_dmem_ram_2846, MEM_stage_inst_dmem_ram_2847, MEM_stage_inst_dmem_ram_2848, MEM_stage_inst_dmem_ram_2849, MEM_stage_inst_dmem_ram_2850, MEM_stage_inst_dmem_ram_2851, MEM_stage_inst_dmem_ram_2852, MEM_stage_inst_dmem_ram_2853, MEM_stage_inst_dmem_ram_2854, MEM_stage_inst_dmem_ram_2855, MEM_stage_inst_dmem_ram_2856, MEM_stage_inst_dmem_ram_2857, MEM_stage_inst_dmem_ram_2858, MEM_stage_inst_dmem_ram_2859, MEM_stage_inst_dmem_ram_2860, MEM_stage_inst_dmem_ram_2861, MEM_stage_inst_dmem_ram_2862, MEM_stage_inst_dmem_ram_2863, MEM_stage_inst_dmem_ram_2864, MEM_stage_inst_dmem_ram_2865, MEM_stage_inst_dmem_ram_2866, MEM_stage_inst_dmem_ram_2867, MEM_stage_inst_dmem_ram_2868, MEM_stage_inst_dmem_ram_2869, MEM_stage_inst_dmem_ram_2870, MEM_stage_inst_dmem_ram_2871, MEM_stage_inst_dmem_ram_2872, MEM_stage_inst_dmem_ram_2873, MEM_stage_inst_dmem_ram_2874, MEM_stage_inst_dmem_ram_2875, MEM_stage_inst_dmem_ram_2876, MEM_stage_inst_dmem_ram_2877, MEM_stage_inst_dmem_ram_2878, MEM_stage_inst_dmem_ram_2879, MEM_stage_inst_dmem_ram_2880, MEM_stage_inst_dmem_ram_2881, MEM_stage_inst_dmem_ram_2882, MEM_stage_inst_dmem_ram_2883, MEM_stage_inst_dmem_ram_2884, MEM_stage_inst_dmem_ram_2885, MEM_stage_inst_dmem_ram_2886, MEM_stage_inst_dmem_ram_2887, MEM_stage_inst_dmem_ram_2888, MEM_stage_inst_dmem_ram_2889, MEM_stage_inst_dmem_ram_2890, MEM_stage_inst_dmem_ram_2891, MEM_stage_inst_dmem_ram_2892, MEM_stage_inst_dmem_ram_2893, MEM_stage_inst_dmem_ram_2894, MEM_stage_inst_dmem_ram_2895, MEM_stage_inst_dmem_ram_2896, MEM_stage_inst_dmem_ram_2897, MEM_stage_inst_dmem_ram_2898, MEM_stage_inst_dmem_ram_2899, MEM_stage_inst_dmem_ram_2900, MEM_stage_inst_dmem_ram_2901, MEM_stage_inst_dmem_ram_2902, MEM_stage_inst_dmem_ram_2903, MEM_stage_inst_dmem_ram_2904, MEM_stage_inst_dmem_ram_2905, MEM_stage_inst_dmem_ram_2906, MEM_stage_inst_dmem_ram_2907, MEM_stage_inst_dmem_ram_2908, MEM_stage_inst_dmem_ram_2909, MEM_stage_inst_dmem_ram_2910, MEM_stage_inst_dmem_ram_2911, MEM_stage_inst_dmem_ram_2912, MEM_stage_inst_dmem_ram_2913, MEM_stage_inst_dmem_ram_2914, MEM_stage_inst_dmem_ram_2915, MEM_stage_inst_dmem_ram_2916, MEM_stage_inst_dmem_ram_2917, MEM_stage_inst_dmem_ram_2918, MEM_stage_inst_dmem_ram_2919, MEM_stage_inst_dmem_ram_2920, MEM_stage_inst_dmem_ram_2921, MEM_stage_inst_dmem_ram_2922, MEM_stage_inst_dmem_ram_2923, MEM_stage_inst_dmem_ram_2924, MEM_stage_inst_dmem_ram_2925, MEM_stage_inst_dmem_ram_2926, MEM_stage_inst_dmem_ram_2927, MEM_stage_inst_dmem_ram_2928, MEM_stage_inst_dmem_ram_2929, MEM_stage_inst_dmem_ram_2930, MEM_stage_inst_dmem_ram_2931, MEM_stage_inst_dmem_ram_2932, MEM_stage_inst_dmem_ram_2933, MEM_stage_inst_dmem_ram_2934, MEM_stage_inst_dmem_ram_2935, MEM_stage_inst_dmem_ram_2936, MEM_stage_inst_dmem_ram_2937, MEM_stage_inst_dmem_ram_2938, MEM_stage_inst_dmem_ram_2939, MEM_stage_inst_dmem_ram_2940, MEM_stage_inst_dmem_ram_2941, MEM_stage_inst_dmem_ram_2942, MEM_stage_inst_dmem_ram_2943, MEM_stage_inst_dmem_ram_2944, MEM_stage_inst_dmem_ram_2945, MEM_stage_inst_dmem_ram_2946, MEM_stage_inst_dmem_ram_2947, MEM_stage_inst_dmem_ram_2948, MEM_stage_inst_dmem_ram_2949, MEM_stage_inst_dmem_ram_2950, MEM_stage_inst_dmem_ram_2951, MEM_stage_inst_dmem_ram_2952, MEM_stage_inst_dmem_ram_2953, MEM_stage_inst_dmem_ram_2954, MEM_stage_inst_dmem_ram_2955, MEM_stage_inst_dmem_ram_2956, MEM_stage_inst_dmem_ram_2957, MEM_stage_inst_dmem_ram_2958, MEM_stage_inst_dmem_ram_2959, MEM_stage_inst_dmem_ram_2960, MEM_stage_inst_dmem_ram_2961, MEM_stage_inst_dmem_ram_2962, MEM_stage_inst_dmem_ram_2963, MEM_stage_inst_dmem_ram_2964, MEM_stage_inst_dmem_ram_2965, MEM_stage_inst_dmem_ram_2966, MEM_stage_inst_dmem_ram_2967, MEM_stage_inst_dmem_ram_2968, MEM_stage_inst_dmem_ram_2969, MEM_stage_inst_dmem_ram_2970, MEM_stage_inst_dmem_ram_2971, MEM_stage_inst_dmem_ram_2972, MEM_stage_inst_dmem_ram_2973, MEM_stage_inst_dmem_ram_2974, MEM_stage_inst_dmem_ram_2975, MEM_stage_inst_dmem_ram_2976, MEM_stage_inst_dmem_ram_2977, MEM_stage_inst_dmem_ram_2978, MEM_stage_inst_dmem_ram_2979, MEM_stage_inst_dmem_ram_2980, MEM_stage_inst_dmem_ram_2981, MEM_stage_inst_dmem_ram_2982, MEM_stage_inst_dmem_ram_2983, MEM_stage_inst_dmem_ram_2984, MEM_stage_inst_dmem_ram_2985, MEM_stage_inst_dmem_ram_2986, MEM_stage_inst_dmem_ram_2987, MEM_stage_inst_dmem_ram_2988, MEM_stage_inst_dmem_ram_2989, MEM_stage_inst_dmem_ram_2990, MEM_stage_inst_dmem_ram_2991, MEM_stage_inst_dmem_ram_2992, MEM_stage_inst_dmem_ram_2993, MEM_stage_inst_dmem_ram_2994, MEM_stage_inst_dmem_ram_2995, MEM_stage_inst_dmem_ram_2996, MEM_stage_inst_dmem_ram_2997, MEM_stage_inst_dmem_ram_2998, MEM_stage_inst_dmem_ram_2999, MEM_stage_inst_dmem_ram_3000, MEM_stage_inst_dmem_ram_3001, MEM_stage_inst_dmem_ram_3002, MEM_stage_inst_dmem_ram_3003, MEM_stage_inst_dmem_ram_3004, MEM_stage_inst_dmem_ram_3005, MEM_stage_inst_dmem_ram_3006, MEM_stage_inst_dmem_ram_3007, MEM_stage_inst_dmem_ram_3008, MEM_stage_inst_dmem_ram_3009, MEM_stage_inst_dmem_ram_3010, MEM_stage_inst_dmem_ram_3011, MEM_stage_inst_dmem_ram_3012, MEM_stage_inst_dmem_ram_3013, MEM_stage_inst_dmem_ram_3014, MEM_stage_inst_dmem_ram_3015, MEM_stage_inst_dmem_ram_3016, MEM_stage_inst_dmem_ram_3017, MEM_stage_inst_dmem_ram_3018, MEM_stage_inst_dmem_ram_3019, MEM_stage_inst_dmem_ram_3020, MEM_stage_inst_dmem_ram_3021, MEM_stage_inst_dmem_ram_3022, MEM_stage_inst_dmem_ram_3023, MEM_stage_inst_dmem_ram_3024, MEM_stage_inst_dmem_ram_3025, MEM_stage_inst_dmem_ram_3026, MEM_stage_inst_dmem_ram_3027, MEM_stage_inst_dmem_ram_3028, MEM_stage_inst_dmem_ram_3029, MEM_stage_inst_dmem_ram_3030, MEM_stage_inst_dmem_ram_3031, MEM_stage_inst_dmem_ram_3032, MEM_stage_inst_dmem_ram_3033, MEM_stage_inst_dmem_ram_3034, MEM_stage_inst_dmem_ram_3035, MEM_stage_inst_dmem_ram_3036, MEM_stage_inst_dmem_ram_3037, MEM_stage_inst_dmem_ram_3038, MEM_stage_inst_dmem_ram_3039, MEM_stage_inst_dmem_ram_3040, MEM_stage_inst_dmem_ram_3041, MEM_stage_inst_dmem_ram_3042, MEM_stage_inst_dmem_ram_3043, MEM_stage_inst_dmem_ram_3044, MEM_stage_inst_dmem_ram_3045, MEM_stage_inst_dmem_ram_3046, MEM_stage_inst_dmem_ram_3047, MEM_stage_inst_dmem_ram_3048, MEM_stage_inst_dmem_ram_3049, MEM_stage_inst_dmem_ram_3050, MEM_stage_inst_dmem_ram_3051, MEM_stage_inst_dmem_ram_3052, MEM_stage_inst_dmem_ram_3053, MEM_stage_inst_dmem_ram_3054, MEM_stage_inst_dmem_ram_3055, MEM_stage_inst_dmem_ram_3056, MEM_stage_inst_dmem_ram_3057, MEM_stage_inst_dmem_ram_3058, MEM_stage_inst_dmem_ram_3059, MEM_stage_inst_dmem_ram_3060, MEM_stage_inst_dmem_ram_3061, MEM_stage_inst_dmem_ram_3062, MEM_stage_inst_dmem_ram_3063, MEM_stage_inst_dmem_ram_3064, MEM_stage_inst_dmem_ram_3065, MEM_stage_inst_dmem_ram_3066, MEM_stage_inst_dmem_ram_3067, MEM_stage_inst_dmem_ram_3068, MEM_stage_inst_dmem_ram_3069, MEM_stage_inst_dmem_ram_3070, MEM_stage_inst_dmem_ram_3071, MEM_stage_inst_dmem_ram_2048, MEM_stage_inst_dmem_ram_2049, MEM_stage_inst_dmem_ram_2050, MEM_stage_inst_dmem_ram_2051, MEM_stage_inst_dmem_ram_2052, MEM_stage_inst_dmem_ram_2053, MEM_stage_inst_dmem_ram_2054, MEM_stage_inst_dmem_ram_2055, MEM_stage_inst_dmem_ram_2056, MEM_stage_inst_dmem_ram_2057, MEM_stage_inst_dmem_ram_2058, MEM_stage_inst_dmem_ram_2059, MEM_stage_inst_dmem_ram_2060, MEM_stage_inst_dmem_ram_2061, MEM_stage_inst_dmem_ram_2062, MEM_stage_inst_dmem_ram_2063, MEM_stage_inst_dmem_ram_2064, MEM_stage_inst_dmem_ram_2065, MEM_stage_inst_dmem_ram_2066, MEM_stage_inst_dmem_ram_2067, MEM_stage_inst_dmem_ram_2068, MEM_stage_inst_dmem_ram_2069, MEM_stage_inst_dmem_ram_2070, MEM_stage_inst_dmem_ram_2071, MEM_stage_inst_dmem_ram_2072, MEM_stage_inst_dmem_ram_2073, MEM_stage_inst_dmem_ram_2074, MEM_stage_inst_dmem_ram_2075, MEM_stage_inst_dmem_ram_2076, MEM_stage_inst_dmem_ram_2077, MEM_stage_inst_dmem_ram_2078, MEM_stage_inst_dmem_ram_2079, MEM_stage_inst_dmem_ram_2080, MEM_stage_inst_dmem_ram_2081, MEM_stage_inst_dmem_ram_2082, MEM_stage_inst_dmem_ram_2083, MEM_stage_inst_dmem_ram_2084, MEM_stage_inst_dmem_ram_2085, MEM_stage_inst_dmem_ram_2086, MEM_stage_inst_dmem_ram_2087, MEM_stage_inst_dmem_ram_2088, MEM_stage_inst_dmem_ram_2089, MEM_stage_inst_dmem_ram_2090, MEM_stage_inst_dmem_ram_2091, MEM_stage_inst_dmem_ram_2092, MEM_stage_inst_dmem_ram_2093, MEM_stage_inst_dmem_ram_2094, MEM_stage_inst_dmem_ram_2095, MEM_stage_inst_dmem_ram_2096, MEM_stage_inst_dmem_ram_2097, MEM_stage_inst_dmem_ram_2098, MEM_stage_inst_dmem_ram_2099, MEM_stage_inst_dmem_ram_2100, MEM_stage_inst_dmem_ram_2101, MEM_stage_inst_dmem_ram_2102, MEM_stage_inst_dmem_ram_2103, MEM_stage_inst_dmem_ram_2104, MEM_stage_inst_dmem_ram_2105, MEM_stage_inst_dmem_ram_2106, MEM_stage_inst_dmem_ram_2107, MEM_stage_inst_dmem_ram_2108, MEM_stage_inst_dmem_ram_2109, MEM_stage_inst_dmem_ram_2110, MEM_stage_inst_dmem_ram_2111, MEM_stage_inst_dmem_ram_2112, MEM_stage_inst_dmem_ram_2113, MEM_stage_inst_dmem_ram_2114, MEM_stage_inst_dmem_ram_2115, MEM_stage_inst_dmem_ram_2116, MEM_stage_inst_dmem_ram_2117, MEM_stage_inst_dmem_ram_2118, MEM_stage_inst_dmem_ram_2119, MEM_stage_inst_dmem_ram_2120, MEM_stage_inst_dmem_ram_2121, MEM_stage_inst_dmem_ram_2122, MEM_stage_inst_dmem_ram_2123, MEM_stage_inst_dmem_ram_2124, MEM_stage_inst_dmem_ram_2125, MEM_stage_inst_dmem_ram_2126, MEM_stage_inst_dmem_ram_2127, MEM_stage_inst_dmem_ram_2128, MEM_stage_inst_dmem_ram_2129, MEM_stage_inst_dmem_ram_2130, MEM_stage_inst_dmem_ram_2131, MEM_stage_inst_dmem_ram_2132, MEM_stage_inst_dmem_ram_2133, MEM_stage_inst_dmem_ram_2134, MEM_stage_inst_dmem_ram_2135, MEM_stage_inst_dmem_ram_2136, MEM_stage_inst_dmem_ram_2137, MEM_stage_inst_dmem_ram_2138, MEM_stage_inst_dmem_ram_2139, MEM_stage_inst_dmem_ram_2140, MEM_stage_inst_dmem_ram_2141, MEM_stage_inst_dmem_ram_2142, MEM_stage_inst_dmem_ram_2143, MEM_stage_inst_dmem_ram_2144, MEM_stage_inst_dmem_ram_2145, MEM_stage_inst_dmem_ram_2146, MEM_stage_inst_dmem_ram_2147, MEM_stage_inst_dmem_ram_2148, MEM_stage_inst_dmem_ram_2149, MEM_stage_inst_dmem_ram_2150, MEM_stage_inst_dmem_ram_2151, MEM_stage_inst_dmem_ram_2152, MEM_stage_inst_dmem_ram_2153, MEM_stage_inst_dmem_ram_2154, MEM_stage_inst_dmem_ram_2155, MEM_stage_inst_dmem_ram_2156, MEM_stage_inst_dmem_ram_2157, MEM_stage_inst_dmem_ram_2158, MEM_stage_inst_dmem_ram_2159, MEM_stage_inst_dmem_ram_2160, MEM_stage_inst_dmem_ram_2161, MEM_stage_inst_dmem_ram_2162, MEM_stage_inst_dmem_ram_2163, MEM_stage_inst_dmem_ram_2164, MEM_stage_inst_dmem_ram_2165, MEM_stage_inst_dmem_ram_2166, MEM_stage_inst_dmem_ram_2167, MEM_stage_inst_dmem_ram_2168, MEM_stage_inst_dmem_ram_2169, MEM_stage_inst_dmem_ram_2170, MEM_stage_inst_dmem_ram_2171, MEM_stage_inst_dmem_ram_2172, MEM_stage_inst_dmem_ram_2173, MEM_stage_inst_dmem_ram_2174, MEM_stage_inst_dmem_ram_2175, MEM_stage_inst_dmem_ram_2176, MEM_stage_inst_dmem_ram_2177, MEM_stage_inst_dmem_ram_2178, MEM_stage_inst_dmem_ram_2179, MEM_stage_inst_dmem_ram_2180, MEM_stage_inst_dmem_ram_2181, MEM_stage_inst_dmem_ram_2182, MEM_stage_inst_dmem_ram_2183, MEM_stage_inst_dmem_ram_2184, MEM_stage_inst_dmem_ram_2185, MEM_stage_inst_dmem_ram_2186, MEM_stage_inst_dmem_ram_2187, MEM_stage_inst_dmem_ram_2188, MEM_stage_inst_dmem_ram_2189, MEM_stage_inst_dmem_ram_2190, MEM_stage_inst_dmem_ram_2191, MEM_stage_inst_dmem_ram_2192, MEM_stage_inst_dmem_ram_2193, MEM_stage_inst_dmem_ram_2194, MEM_stage_inst_dmem_ram_2195, MEM_stage_inst_dmem_ram_2196, MEM_stage_inst_dmem_ram_2197, MEM_stage_inst_dmem_ram_2198, MEM_stage_inst_dmem_ram_2199, MEM_stage_inst_dmem_ram_2200, MEM_stage_inst_dmem_ram_2201, MEM_stage_inst_dmem_ram_2202, MEM_stage_inst_dmem_ram_2203, MEM_stage_inst_dmem_ram_2204, MEM_stage_inst_dmem_ram_2205, MEM_stage_inst_dmem_ram_2206, MEM_stage_inst_dmem_ram_2207, MEM_stage_inst_dmem_ram_2208, MEM_stage_inst_dmem_ram_2209, MEM_stage_inst_dmem_ram_2210, MEM_stage_inst_dmem_ram_2211, MEM_stage_inst_dmem_ram_2212, MEM_stage_inst_dmem_ram_2213, MEM_stage_inst_dmem_ram_2214, MEM_stage_inst_dmem_ram_2215, MEM_stage_inst_dmem_ram_2216, MEM_stage_inst_dmem_ram_2217, MEM_stage_inst_dmem_ram_2218, MEM_stage_inst_dmem_ram_2219, MEM_stage_inst_dmem_ram_2220, MEM_stage_inst_dmem_ram_2221, MEM_stage_inst_dmem_ram_2222, MEM_stage_inst_dmem_ram_2223, MEM_stage_inst_dmem_ram_2224, MEM_stage_inst_dmem_ram_2225, MEM_stage_inst_dmem_ram_2226, MEM_stage_inst_dmem_ram_2227, MEM_stage_inst_dmem_ram_2228, MEM_stage_inst_dmem_ram_2229, MEM_stage_inst_dmem_ram_2230, MEM_stage_inst_dmem_ram_2231, MEM_stage_inst_dmem_ram_2232, MEM_stage_inst_dmem_ram_2233, MEM_stage_inst_dmem_ram_2234, MEM_stage_inst_dmem_ram_2235, MEM_stage_inst_dmem_ram_2236, MEM_stage_inst_dmem_ram_2237, MEM_stage_inst_dmem_ram_2238, MEM_stage_inst_dmem_ram_2239, MEM_stage_inst_dmem_ram_2240, MEM_stage_inst_dmem_ram_2241, MEM_stage_inst_dmem_ram_2242, MEM_stage_inst_dmem_ram_2243, MEM_stage_inst_dmem_ram_2244, MEM_stage_inst_dmem_ram_2245, MEM_stage_inst_dmem_ram_2246, MEM_stage_inst_dmem_ram_2247, MEM_stage_inst_dmem_ram_2248, MEM_stage_inst_dmem_ram_2249, MEM_stage_inst_dmem_ram_2250, MEM_stage_inst_dmem_ram_2251, MEM_stage_inst_dmem_ram_2252, MEM_stage_inst_dmem_ram_2253, MEM_stage_inst_dmem_ram_2254, MEM_stage_inst_dmem_ram_2255, MEM_stage_inst_dmem_ram_2256, MEM_stage_inst_dmem_ram_2257, MEM_stage_inst_dmem_ram_2258, MEM_stage_inst_dmem_ram_2259, MEM_stage_inst_dmem_ram_2260, MEM_stage_inst_dmem_ram_2261, MEM_stage_inst_dmem_ram_2262, MEM_stage_inst_dmem_ram_2263, MEM_stage_inst_dmem_ram_2264, MEM_stage_inst_dmem_ram_2265, MEM_stage_inst_dmem_ram_2266, MEM_stage_inst_dmem_ram_2267, MEM_stage_inst_dmem_ram_2268, MEM_stage_inst_dmem_ram_2269, MEM_stage_inst_dmem_ram_2270, MEM_stage_inst_dmem_ram_2271, MEM_stage_inst_dmem_ram_2272, MEM_stage_inst_dmem_ram_2273, MEM_stage_inst_dmem_ram_2274, MEM_stage_inst_dmem_ram_2275, MEM_stage_inst_dmem_ram_2276, MEM_stage_inst_dmem_ram_2277, MEM_stage_inst_dmem_ram_2278, MEM_stage_inst_dmem_ram_2279, MEM_stage_inst_dmem_ram_2280, MEM_stage_inst_dmem_ram_2281, MEM_stage_inst_dmem_ram_2282, MEM_stage_inst_dmem_ram_2283, MEM_stage_inst_dmem_ram_2284, MEM_stage_inst_dmem_ram_2285, MEM_stage_inst_dmem_ram_2286, MEM_stage_inst_dmem_ram_2287, MEM_stage_inst_dmem_ram_2288, MEM_stage_inst_dmem_ram_2289, MEM_stage_inst_dmem_ram_2290, MEM_stage_inst_dmem_ram_2291, MEM_stage_inst_dmem_ram_2292, MEM_stage_inst_dmem_ram_2293, MEM_stage_inst_dmem_ram_2294, MEM_stage_inst_dmem_ram_2295, MEM_stage_inst_dmem_ram_2296, MEM_stage_inst_dmem_ram_2297, MEM_stage_inst_dmem_ram_2298, MEM_stage_inst_dmem_ram_2299, MEM_stage_inst_dmem_ram_2300, MEM_stage_inst_dmem_ram_2301, MEM_stage_inst_dmem_ram_2302, MEM_stage_inst_dmem_ram_2303, MEM_stage_inst_dmem_ram_2304, MEM_stage_inst_dmem_ram_2305, MEM_stage_inst_dmem_ram_2306, MEM_stage_inst_dmem_ram_2307, MEM_stage_inst_dmem_ram_2308, MEM_stage_inst_dmem_ram_2309, MEM_stage_inst_dmem_ram_2310, MEM_stage_inst_dmem_ram_2311, MEM_stage_inst_dmem_ram_2312, MEM_stage_inst_dmem_ram_2313, MEM_stage_inst_dmem_ram_2314, MEM_stage_inst_dmem_ram_2315, MEM_stage_inst_dmem_ram_2316, MEM_stage_inst_dmem_ram_2317, MEM_stage_inst_dmem_ram_2318, MEM_stage_inst_dmem_ram_2319, MEM_stage_inst_dmem_ram_2320, MEM_stage_inst_dmem_ram_2321, MEM_stage_inst_dmem_ram_2322, MEM_stage_inst_dmem_ram_2323, MEM_stage_inst_dmem_ram_2324, MEM_stage_inst_dmem_ram_2325, MEM_stage_inst_dmem_ram_2326, MEM_stage_inst_dmem_ram_2327, MEM_stage_inst_dmem_ram_2328, MEM_stage_inst_dmem_ram_2329, MEM_stage_inst_dmem_ram_2330, MEM_stage_inst_dmem_ram_2331, MEM_stage_inst_dmem_ram_2332, MEM_stage_inst_dmem_ram_2333, MEM_stage_inst_dmem_ram_2334, MEM_stage_inst_dmem_ram_2335, MEM_stage_inst_dmem_ram_2336, MEM_stage_inst_dmem_ram_2337, MEM_stage_inst_dmem_ram_2338, MEM_stage_inst_dmem_ram_2339, MEM_stage_inst_dmem_ram_2340, MEM_stage_inst_dmem_ram_2341, MEM_stage_inst_dmem_ram_2342, MEM_stage_inst_dmem_ram_2343, MEM_stage_inst_dmem_ram_2344, MEM_stage_inst_dmem_ram_2345, MEM_stage_inst_dmem_ram_2346, MEM_stage_inst_dmem_ram_2347, MEM_stage_inst_dmem_ram_2348, MEM_stage_inst_dmem_ram_2349, MEM_stage_inst_dmem_ram_2350, MEM_stage_inst_dmem_ram_2351, MEM_stage_inst_dmem_ram_2352, MEM_stage_inst_dmem_ram_2353, MEM_stage_inst_dmem_ram_2354, MEM_stage_inst_dmem_ram_2355, MEM_stage_inst_dmem_ram_2356, MEM_stage_inst_dmem_ram_2357, MEM_stage_inst_dmem_ram_2358, MEM_stage_inst_dmem_ram_2359, MEM_stage_inst_dmem_ram_2360, MEM_stage_inst_dmem_ram_2361, MEM_stage_inst_dmem_ram_2362, MEM_stage_inst_dmem_ram_2363, MEM_stage_inst_dmem_ram_2364, MEM_stage_inst_dmem_ram_2365, MEM_stage_inst_dmem_ram_2366, MEM_stage_inst_dmem_ram_2367, MEM_stage_inst_dmem_ram_2368, MEM_stage_inst_dmem_ram_2369, MEM_stage_inst_dmem_ram_2370, MEM_stage_inst_dmem_ram_2371, MEM_stage_inst_dmem_ram_2372, MEM_stage_inst_dmem_ram_2373, MEM_stage_inst_dmem_ram_2374, MEM_stage_inst_dmem_ram_2375, MEM_stage_inst_dmem_ram_2376, MEM_stage_inst_dmem_ram_2377, MEM_stage_inst_dmem_ram_2378, MEM_stage_inst_dmem_ram_2379, MEM_stage_inst_dmem_ram_2380, MEM_stage_inst_dmem_ram_2381, MEM_stage_inst_dmem_ram_2382, MEM_stage_inst_dmem_ram_2383, MEM_stage_inst_dmem_ram_2384, MEM_stage_inst_dmem_ram_2385, MEM_stage_inst_dmem_ram_2386, MEM_stage_inst_dmem_ram_2387, MEM_stage_inst_dmem_ram_2388, MEM_stage_inst_dmem_ram_2389, MEM_stage_inst_dmem_ram_2390, MEM_stage_inst_dmem_ram_2391, MEM_stage_inst_dmem_ram_2392, MEM_stage_inst_dmem_ram_2393, MEM_stage_inst_dmem_ram_2394, MEM_stage_inst_dmem_ram_2395, MEM_stage_inst_dmem_ram_2396, MEM_stage_inst_dmem_ram_2397, MEM_stage_inst_dmem_ram_2398, MEM_stage_inst_dmem_ram_2399, MEM_stage_inst_dmem_ram_2400, MEM_stage_inst_dmem_ram_2401, MEM_stage_inst_dmem_ram_2402, MEM_stage_inst_dmem_ram_2403, MEM_stage_inst_dmem_ram_2404, MEM_stage_inst_dmem_ram_2405, MEM_stage_inst_dmem_ram_2406, MEM_stage_inst_dmem_ram_2407, MEM_stage_inst_dmem_ram_2408, MEM_stage_inst_dmem_ram_2409, MEM_stage_inst_dmem_ram_2410, MEM_stage_inst_dmem_ram_2411, MEM_stage_inst_dmem_ram_2412, MEM_stage_inst_dmem_ram_2413, MEM_stage_inst_dmem_ram_2414, MEM_stage_inst_dmem_ram_2415, MEM_stage_inst_dmem_ram_2416, MEM_stage_inst_dmem_ram_2417, MEM_stage_inst_dmem_ram_2418, MEM_stage_inst_dmem_ram_2419, MEM_stage_inst_dmem_ram_2420, MEM_stage_inst_dmem_ram_2421, MEM_stage_inst_dmem_ram_2422, MEM_stage_inst_dmem_ram_2423, MEM_stage_inst_dmem_ram_2424, MEM_stage_inst_dmem_ram_2425, MEM_stage_inst_dmem_ram_2426, MEM_stage_inst_dmem_ram_2427, MEM_stage_inst_dmem_ram_2428, MEM_stage_inst_dmem_ram_2429, MEM_stage_inst_dmem_ram_2430, MEM_stage_inst_dmem_ram_2431, MEM_stage_inst_dmem_ram_2432, MEM_stage_inst_dmem_ram_2433, MEM_stage_inst_dmem_ram_2434, MEM_stage_inst_dmem_ram_2435, MEM_stage_inst_dmem_ram_2436, MEM_stage_inst_dmem_ram_2437, MEM_stage_inst_dmem_ram_2438, MEM_stage_inst_dmem_ram_2439, MEM_stage_inst_dmem_ram_2440, MEM_stage_inst_dmem_ram_2441, MEM_stage_inst_dmem_ram_2442, MEM_stage_inst_dmem_ram_2443, MEM_stage_inst_dmem_ram_2444, MEM_stage_inst_dmem_ram_2445, MEM_stage_inst_dmem_ram_2446, MEM_stage_inst_dmem_ram_2447, MEM_stage_inst_dmem_ram_2448, MEM_stage_inst_dmem_ram_2449, MEM_stage_inst_dmem_ram_2450, MEM_stage_inst_dmem_ram_2451, MEM_stage_inst_dmem_ram_2452, MEM_stage_inst_dmem_ram_2453, MEM_stage_inst_dmem_ram_2454, MEM_stage_inst_dmem_ram_2455, MEM_stage_inst_dmem_ram_2456, MEM_stage_inst_dmem_ram_2457, MEM_stage_inst_dmem_ram_2458, MEM_stage_inst_dmem_ram_2459, MEM_stage_inst_dmem_ram_2460, MEM_stage_inst_dmem_ram_2461, MEM_stage_inst_dmem_ram_2462, MEM_stage_inst_dmem_ram_2463, MEM_stage_inst_dmem_ram_2464, MEM_stage_inst_dmem_ram_2465, MEM_stage_inst_dmem_ram_2466, MEM_stage_inst_dmem_ram_2467, MEM_stage_inst_dmem_ram_2468, MEM_stage_inst_dmem_ram_2469, MEM_stage_inst_dmem_ram_2470, MEM_stage_inst_dmem_ram_2471, MEM_stage_inst_dmem_ram_2472, MEM_stage_inst_dmem_ram_2473, MEM_stage_inst_dmem_ram_2474, MEM_stage_inst_dmem_ram_2475, MEM_stage_inst_dmem_ram_2476, MEM_stage_inst_dmem_ram_2477, MEM_stage_inst_dmem_ram_2478, MEM_stage_inst_dmem_ram_2479, MEM_stage_inst_dmem_ram_2480, MEM_stage_inst_dmem_ram_2481, MEM_stage_inst_dmem_ram_2482, MEM_stage_inst_dmem_ram_2483, MEM_stage_inst_dmem_ram_2484, MEM_stage_inst_dmem_ram_2485, MEM_stage_inst_dmem_ram_2486, MEM_stage_inst_dmem_ram_2487, MEM_stage_inst_dmem_ram_2488, MEM_stage_inst_dmem_ram_2489, MEM_stage_inst_dmem_ram_2490, MEM_stage_inst_dmem_ram_2491, MEM_stage_inst_dmem_ram_2492, MEM_stage_inst_dmem_ram_2493, MEM_stage_inst_dmem_ram_2494, MEM_stage_inst_dmem_ram_2495, MEM_stage_inst_dmem_ram_2496, MEM_stage_inst_dmem_ram_2497, MEM_stage_inst_dmem_ram_2498, MEM_stage_inst_dmem_ram_2499, MEM_stage_inst_dmem_ram_2500, MEM_stage_inst_dmem_ram_2501, MEM_stage_inst_dmem_ram_2502, MEM_stage_inst_dmem_ram_2503, MEM_stage_inst_dmem_ram_2504, MEM_stage_inst_dmem_ram_2505, MEM_stage_inst_dmem_ram_2506, MEM_stage_inst_dmem_ram_2507, MEM_stage_inst_dmem_ram_2508, MEM_stage_inst_dmem_ram_2509, MEM_stage_inst_dmem_ram_2510, MEM_stage_inst_dmem_ram_2511, MEM_stage_inst_dmem_ram_2512, MEM_stage_inst_dmem_ram_2513, MEM_stage_inst_dmem_ram_2514, MEM_stage_inst_dmem_ram_2515, MEM_stage_inst_dmem_ram_2516, MEM_stage_inst_dmem_ram_2517, MEM_stage_inst_dmem_ram_2518, MEM_stage_inst_dmem_ram_2519, MEM_stage_inst_dmem_ram_2520, MEM_stage_inst_dmem_ram_2521, MEM_stage_inst_dmem_ram_2522, MEM_stage_inst_dmem_ram_2523, MEM_stage_inst_dmem_ram_2524, MEM_stage_inst_dmem_ram_2525, MEM_stage_inst_dmem_ram_2526, MEM_stage_inst_dmem_ram_2527, MEM_stage_inst_dmem_ram_2528, MEM_stage_inst_dmem_ram_2529, MEM_stage_inst_dmem_ram_2530, MEM_stage_inst_dmem_ram_2531, MEM_stage_inst_dmem_ram_2532, MEM_stage_inst_dmem_ram_2533, MEM_stage_inst_dmem_ram_2534, MEM_stage_inst_dmem_ram_2535, MEM_stage_inst_dmem_ram_2536, MEM_stage_inst_dmem_ram_2537, MEM_stage_inst_dmem_ram_2538, MEM_stage_inst_dmem_ram_2539, MEM_stage_inst_dmem_ram_2540, MEM_stage_inst_dmem_ram_2541, MEM_stage_inst_dmem_ram_2542, MEM_stage_inst_dmem_ram_2543, MEM_stage_inst_dmem_ram_2544, MEM_stage_inst_dmem_ram_2545, MEM_stage_inst_dmem_ram_2546, MEM_stage_inst_dmem_ram_2547, MEM_stage_inst_dmem_ram_2548, MEM_stage_inst_dmem_ram_2549, MEM_stage_inst_dmem_ram_2550, MEM_stage_inst_dmem_ram_2551, MEM_stage_inst_dmem_ram_2552, MEM_stage_inst_dmem_ram_2553, MEM_stage_inst_dmem_ram_2554, MEM_stage_inst_dmem_ram_2555, MEM_stage_inst_dmem_ram_2556, MEM_stage_inst_dmem_ram_2557, MEM_stage_inst_dmem_ram_2558, MEM_stage_inst_dmem_ram_2559, MEM_stage_inst_dmem_ram_1536, MEM_stage_inst_dmem_ram_1537, MEM_stage_inst_dmem_ram_1538, MEM_stage_inst_dmem_ram_1539, MEM_stage_inst_dmem_ram_1540, MEM_stage_inst_dmem_ram_1541, MEM_stage_inst_dmem_ram_1542, MEM_stage_inst_dmem_ram_1543, MEM_stage_inst_dmem_ram_1544, MEM_stage_inst_dmem_ram_1545, MEM_stage_inst_dmem_ram_1546, MEM_stage_inst_dmem_ram_1547, MEM_stage_inst_dmem_ram_1548, MEM_stage_inst_dmem_ram_1549, MEM_stage_inst_dmem_ram_1550, MEM_stage_inst_dmem_ram_1551, MEM_stage_inst_dmem_ram_1552, MEM_stage_inst_dmem_ram_1553, MEM_stage_inst_dmem_ram_1554, MEM_stage_inst_dmem_ram_1555, MEM_stage_inst_dmem_ram_1556, MEM_stage_inst_dmem_ram_1557, MEM_stage_inst_dmem_ram_1558, MEM_stage_inst_dmem_ram_1559, MEM_stage_inst_dmem_ram_1560, MEM_stage_inst_dmem_ram_1561, MEM_stage_inst_dmem_ram_1562, MEM_stage_inst_dmem_ram_1563, MEM_stage_inst_dmem_ram_1564, MEM_stage_inst_dmem_ram_1565, MEM_stage_inst_dmem_ram_1566, MEM_stage_inst_dmem_ram_1567, MEM_stage_inst_dmem_ram_1568, MEM_stage_inst_dmem_ram_1569, MEM_stage_inst_dmem_ram_1570, MEM_stage_inst_dmem_ram_1571, MEM_stage_inst_dmem_ram_1572, MEM_stage_inst_dmem_ram_1573, MEM_stage_inst_dmem_ram_1574, MEM_stage_inst_dmem_ram_1575, MEM_stage_inst_dmem_ram_1576, MEM_stage_inst_dmem_ram_1577, MEM_stage_inst_dmem_ram_1578, MEM_stage_inst_dmem_ram_1579, MEM_stage_inst_dmem_ram_1580, MEM_stage_inst_dmem_ram_1581, MEM_stage_inst_dmem_ram_1582, MEM_stage_inst_dmem_ram_1583, MEM_stage_inst_dmem_ram_1584, MEM_stage_inst_dmem_ram_1585, MEM_stage_inst_dmem_ram_1586, MEM_stage_inst_dmem_ram_1587, MEM_stage_inst_dmem_ram_1588, MEM_stage_inst_dmem_ram_1589, MEM_stage_inst_dmem_ram_1590, MEM_stage_inst_dmem_ram_1591, MEM_stage_inst_dmem_ram_1592, MEM_stage_inst_dmem_ram_1593, MEM_stage_inst_dmem_ram_1594, MEM_stage_inst_dmem_ram_1595, MEM_stage_inst_dmem_ram_1596, MEM_stage_inst_dmem_ram_1597, MEM_stage_inst_dmem_ram_1598, MEM_stage_inst_dmem_ram_1599, MEM_stage_inst_dmem_ram_1600, MEM_stage_inst_dmem_ram_1601, MEM_stage_inst_dmem_ram_1602, MEM_stage_inst_dmem_ram_1603, MEM_stage_inst_dmem_ram_1604, MEM_stage_inst_dmem_ram_1605, MEM_stage_inst_dmem_ram_1606, MEM_stage_inst_dmem_ram_1607, MEM_stage_inst_dmem_ram_1608, MEM_stage_inst_dmem_ram_1609, MEM_stage_inst_dmem_ram_1610, MEM_stage_inst_dmem_ram_1611, MEM_stage_inst_dmem_ram_1612, MEM_stage_inst_dmem_ram_1613, MEM_stage_inst_dmem_ram_1614, MEM_stage_inst_dmem_ram_1615, MEM_stage_inst_dmem_ram_1616, MEM_stage_inst_dmem_ram_1617, MEM_stage_inst_dmem_ram_1618, MEM_stage_inst_dmem_ram_1619, MEM_stage_inst_dmem_ram_1620, MEM_stage_inst_dmem_ram_1621, MEM_stage_inst_dmem_ram_1622, MEM_stage_inst_dmem_ram_1623, MEM_stage_inst_dmem_ram_1624, MEM_stage_inst_dmem_ram_1625, MEM_stage_inst_dmem_ram_1626, MEM_stage_inst_dmem_ram_1627, MEM_stage_inst_dmem_ram_1628, MEM_stage_inst_dmem_ram_1629, MEM_stage_inst_dmem_ram_1630, MEM_stage_inst_dmem_ram_1631, MEM_stage_inst_dmem_ram_1632, MEM_stage_inst_dmem_ram_1633, MEM_stage_inst_dmem_ram_1634, MEM_stage_inst_dmem_ram_1635, MEM_stage_inst_dmem_ram_1636, MEM_stage_inst_dmem_ram_1637, MEM_stage_inst_dmem_ram_1638, MEM_stage_inst_dmem_ram_1639, MEM_stage_inst_dmem_ram_1640, MEM_stage_inst_dmem_ram_1641, MEM_stage_inst_dmem_ram_1642, MEM_stage_inst_dmem_ram_1643, MEM_stage_inst_dmem_ram_1644, MEM_stage_inst_dmem_ram_1645, MEM_stage_inst_dmem_ram_1646, MEM_stage_inst_dmem_ram_1647, MEM_stage_inst_dmem_ram_1648, MEM_stage_inst_dmem_ram_1649, MEM_stage_inst_dmem_ram_1650, MEM_stage_inst_dmem_ram_1651, MEM_stage_inst_dmem_ram_1652, MEM_stage_inst_dmem_ram_1653, MEM_stage_inst_dmem_ram_1654, MEM_stage_inst_dmem_ram_1655, MEM_stage_inst_dmem_ram_1656, MEM_stage_inst_dmem_ram_1657, MEM_stage_inst_dmem_ram_1658, MEM_stage_inst_dmem_ram_1659, MEM_stage_inst_dmem_ram_1660, MEM_stage_inst_dmem_ram_1661, MEM_stage_inst_dmem_ram_1662, MEM_stage_inst_dmem_ram_1663, MEM_stage_inst_dmem_ram_1664, MEM_stage_inst_dmem_ram_1665, MEM_stage_inst_dmem_ram_1666, MEM_stage_inst_dmem_ram_1667, MEM_stage_inst_dmem_ram_1668, MEM_stage_inst_dmem_ram_1669, MEM_stage_inst_dmem_ram_1670, MEM_stage_inst_dmem_ram_1671, MEM_stage_inst_dmem_ram_1672, MEM_stage_inst_dmem_ram_1673, MEM_stage_inst_dmem_ram_1674, MEM_stage_inst_dmem_ram_1675, MEM_stage_inst_dmem_ram_1676, MEM_stage_inst_dmem_ram_1677, MEM_stage_inst_dmem_ram_1678, MEM_stage_inst_dmem_ram_1679, MEM_stage_inst_dmem_ram_1680, MEM_stage_inst_dmem_ram_1681, MEM_stage_inst_dmem_ram_1682, MEM_stage_inst_dmem_ram_1683, MEM_stage_inst_dmem_ram_1684, MEM_stage_inst_dmem_ram_1685, MEM_stage_inst_dmem_ram_1686, MEM_stage_inst_dmem_ram_1687, MEM_stage_inst_dmem_ram_1688, MEM_stage_inst_dmem_ram_1689, MEM_stage_inst_dmem_ram_1690, MEM_stage_inst_dmem_ram_1691, MEM_stage_inst_dmem_ram_1692, MEM_stage_inst_dmem_ram_1693, MEM_stage_inst_dmem_ram_1694, MEM_stage_inst_dmem_ram_1695, MEM_stage_inst_dmem_ram_1696, MEM_stage_inst_dmem_ram_1697, MEM_stage_inst_dmem_ram_1698, MEM_stage_inst_dmem_ram_1699, MEM_stage_inst_dmem_ram_1700, MEM_stage_inst_dmem_ram_1701, MEM_stage_inst_dmem_ram_1702, MEM_stage_inst_dmem_ram_1703, MEM_stage_inst_dmem_ram_1704, MEM_stage_inst_dmem_ram_1705, MEM_stage_inst_dmem_ram_1706, MEM_stage_inst_dmem_ram_1707, MEM_stage_inst_dmem_ram_1708, MEM_stage_inst_dmem_ram_1709, MEM_stage_inst_dmem_ram_1710, MEM_stage_inst_dmem_ram_1711, MEM_stage_inst_dmem_ram_1712, MEM_stage_inst_dmem_ram_1713, MEM_stage_inst_dmem_ram_1714, MEM_stage_inst_dmem_ram_1715, MEM_stage_inst_dmem_ram_1716, MEM_stage_inst_dmem_ram_1717, MEM_stage_inst_dmem_ram_1718, MEM_stage_inst_dmem_ram_1719, MEM_stage_inst_dmem_ram_1720, MEM_stage_inst_dmem_ram_1721, MEM_stage_inst_dmem_ram_1722, MEM_stage_inst_dmem_ram_1723, MEM_stage_inst_dmem_ram_1724, MEM_stage_inst_dmem_ram_1725, MEM_stage_inst_dmem_ram_1726, MEM_stage_inst_dmem_ram_1727, MEM_stage_inst_dmem_ram_1728, MEM_stage_inst_dmem_ram_1729, MEM_stage_inst_dmem_ram_1730, MEM_stage_inst_dmem_ram_1731, MEM_stage_inst_dmem_ram_1732, MEM_stage_inst_dmem_ram_1733, MEM_stage_inst_dmem_ram_1734, MEM_stage_inst_dmem_ram_1735, MEM_stage_inst_dmem_ram_1736, MEM_stage_inst_dmem_ram_1737, MEM_stage_inst_dmem_ram_1738, MEM_stage_inst_dmem_ram_1739, MEM_stage_inst_dmem_ram_1740, MEM_stage_inst_dmem_ram_1741, MEM_stage_inst_dmem_ram_1742, MEM_stage_inst_dmem_ram_1743, MEM_stage_inst_dmem_ram_1744, MEM_stage_inst_dmem_ram_1745, MEM_stage_inst_dmem_ram_1746, MEM_stage_inst_dmem_ram_1747, MEM_stage_inst_dmem_ram_1748, MEM_stage_inst_dmem_ram_1749, MEM_stage_inst_dmem_ram_1750, MEM_stage_inst_dmem_ram_1751, MEM_stage_inst_dmem_ram_1752, MEM_stage_inst_dmem_ram_1753, MEM_stage_inst_dmem_ram_1754, MEM_stage_inst_dmem_ram_1755, MEM_stage_inst_dmem_ram_1756, MEM_stage_inst_dmem_ram_1757, MEM_stage_inst_dmem_ram_1758, MEM_stage_inst_dmem_ram_1759, MEM_stage_inst_dmem_ram_1760, MEM_stage_inst_dmem_ram_1761, MEM_stage_inst_dmem_ram_1762, MEM_stage_inst_dmem_ram_1763, MEM_stage_inst_dmem_ram_1764, MEM_stage_inst_dmem_ram_1765, MEM_stage_inst_dmem_ram_1766, MEM_stage_inst_dmem_ram_1767, MEM_stage_inst_dmem_ram_1768, MEM_stage_inst_dmem_ram_1769, MEM_stage_inst_dmem_ram_1770, MEM_stage_inst_dmem_ram_1771, MEM_stage_inst_dmem_ram_1772, MEM_stage_inst_dmem_ram_1773, MEM_stage_inst_dmem_ram_1774, MEM_stage_inst_dmem_ram_1775, MEM_stage_inst_dmem_ram_1776, MEM_stage_inst_dmem_ram_1777, MEM_stage_inst_dmem_ram_1778, MEM_stage_inst_dmem_ram_1779, MEM_stage_inst_dmem_ram_1780, MEM_stage_inst_dmem_ram_1781, MEM_stage_inst_dmem_ram_1782, MEM_stage_inst_dmem_ram_1783, MEM_stage_inst_dmem_ram_1784, MEM_stage_inst_dmem_ram_1785, MEM_stage_inst_dmem_ram_1786, MEM_stage_inst_dmem_ram_1787, MEM_stage_inst_dmem_ram_1788, MEM_stage_inst_dmem_ram_1789, MEM_stage_inst_dmem_ram_1790, MEM_stage_inst_dmem_ram_1791, MEM_stage_inst_dmem_ram_1792, MEM_stage_inst_dmem_ram_1793, MEM_stage_inst_dmem_ram_1794, MEM_stage_inst_dmem_ram_1795, MEM_stage_inst_dmem_ram_1796, MEM_stage_inst_dmem_ram_1797, MEM_stage_inst_dmem_ram_1798, MEM_stage_inst_dmem_ram_1799, MEM_stage_inst_dmem_ram_1800, MEM_stage_inst_dmem_ram_1801, MEM_stage_inst_dmem_ram_1802, MEM_stage_inst_dmem_ram_1803, MEM_stage_inst_dmem_ram_1804, MEM_stage_inst_dmem_ram_1805, MEM_stage_inst_dmem_ram_1806, MEM_stage_inst_dmem_ram_1807, MEM_stage_inst_dmem_ram_1808, MEM_stage_inst_dmem_ram_1809, MEM_stage_inst_dmem_ram_1810, MEM_stage_inst_dmem_ram_1811, MEM_stage_inst_dmem_ram_1812, MEM_stage_inst_dmem_ram_1813, MEM_stage_inst_dmem_ram_1814, MEM_stage_inst_dmem_ram_1815, MEM_stage_inst_dmem_ram_1816, MEM_stage_inst_dmem_ram_1817, MEM_stage_inst_dmem_ram_1818, MEM_stage_inst_dmem_ram_1819, MEM_stage_inst_dmem_ram_1820, MEM_stage_inst_dmem_ram_1821, MEM_stage_inst_dmem_ram_1822, MEM_stage_inst_dmem_ram_1823, MEM_stage_inst_dmem_ram_1824, MEM_stage_inst_dmem_ram_1825, MEM_stage_inst_dmem_ram_1826, MEM_stage_inst_dmem_ram_1827, MEM_stage_inst_dmem_ram_1828, MEM_stage_inst_dmem_ram_1829, MEM_stage_inst_dmem_ram_1830, MEM_stage_inst_dmem_ram_1831, MEM_stage_inst_dmem_ram_1832, MEM_stage_inst_dmem_ram_1833, MEM_stage_inst_dmem_ram_1834, MEM_stage_inst_dmem_ram_1835, MEM_stage_inst_dmem_ram_1836, MEM_stage_inst_dmem_ram_1837, MEM_stage_inst_dmem_ram_1838, MEM_stage_inst_dmem_ram_1839, MEM_stage_inst_dmem_ram_1840, MEM_stage_inst_dmem_ram_1841, MEM_stage_inst_dmem_ram_1842, MEM_stage_inst_dmem_ram_1843, MEM_stage_inst_dmem_ram_1844, MEM_stage_inst_dmem_ram_1845, MEM_stage_inst_dmem_ram_1846, MEM_stage_inst_dmem_ram_1847, MEM_stage_inst_dmem_ram_1848, MEM_stage_inst_dmem_ram_1849, MEM_stage_inst_dmem_ram_1850, MEM_stage_inst_dmem_ram_1851, MEM_stage_inst_dmem_ram_1852, MEM_stage_inst_dmem_ram_1853, MEM_stage_inst_dmem_ram_1854, MEM_stage_inst_dmem_ram_1855, MEM_stage_inst_dmem_ram_1856, MEM_stage_inst_dmem_ram_1857, MEM_stage_inst_dmem_ram_1858, MEM_stage_inst_dmem_ram_1859, MEM_stage_inst_dmem_ram_1860, MEM_stage_inst_dmem_ram_1861, MEM_stage_inst_dmem_ram_1862, MEM_stage_inst_dmem_ram_1863, MEM_stage_inst_dmem_ram_1864, MEM_stage_inst_dmem_ram_1865, MEM_stage_inst_dmem_ram_1866, MEM_stage_inst_dmem_ram_1867, MEM_stage_inst_dmem_ram_1868, MEM_stage_inst_dmem_ram_1869, MEM_stage_inst_dmem_ram_1870, MEM_stage_inst_dmem_ram_1871, MEM_stage_inst_dmem_ram_1872, MEM_stage_inst_dmem_ram_1873, MEM_stage_inst_dmem_ram_1874, MEM_stage_inst_dmem_ram_1875, MEM_stage_inst_dmem_ram_1876, MEM_stage_inst_dmem_ram_1877, MEM_stage_inst_dmem_ram_1878, MEM_stage_inst_dmem_ram_1879, MEM_stage_inst_dmem_ram_1880, MEM_stage_inst_dmem_ram_1881, MEM_stage_inst_dmem_ram_1882, MEM_stage_inst_dmem_ram_1883, MEM_stage_inst_dmem_ram_1884, MEM_stage_inst_dmem_ram_1885, MEM_stage_inst_dmem_ram_1886, MEM_stage_inst_dmem_ram_1887, MEM_stage_inst_dmem_ram_1888, MEM_stage_inst_dmem_ram_1889, MEM_stage_inst_dmem_ram_1890, MEM_stage_inst_dmem_ram_1891, MEM_stage_inst_dmem_ram_1892, MEM_stage_inst_dmem_ram_1893, MEM_stage_inst_dmem_ram_1894, MEM_stage_inst_dmem_ram_1895, MEM_stage_inst_dmem_ram_1896, MEM_stage_inst_dmem_ram_1897, MEM_stage_inst_dmem_ram_1898, MEM_stage_inst_dmem_ram_1899, MEM_stage_inst_dmem_ram_1900, MEM_stage_inst_dmem_ram_1901, MEM_stage_inst_dmem_ram_1902, MEM_stage_inst_dmem_ram_1903, MEM_stage_inst_dmem_ram_1904, MEM_stage_inst_dmem_ram_1905, MEM_stage_inst_dmem_ram_1906, MEM_stage_inst_dmem_ram_1907, MEM_stage_inst_dmem_ram_1908, MEM_stage_inst_dmem_ram_1909, MEM_stage_inst_dmem_ram_1910, MEM_stage_inst_dmem_ram_1911, MEM_stage_inst_dmem_ram_1912, MEM_stage_inst_dmem_ram_1913, MEM_stage_inst_dmem_ram_1914, MEM_stage_inst_dmem_ram_1915, MEM_stage_inst_dmem_ram_1916, MEM_stage_inst_dmem_ram_1917, MEM_stage_inst_dmem_ram_1918, MEM_stage_inst_dmem_ram_1919, MEM_stage_inst_dmem_ram_1920, MEM_stage_inst_dmem_ram_1921, MEM_stage_inst_dmem_ram_1922, MEM_stage_inst_dmem_ram_1923, MEM_stage_inst_dmem_ram_1924, MEM_stage_inst_dmem_ram_1925, MEM_stage_inst_dmem_ram_1926, MEM_stage_inst_dmem_ram_1927, MEM_stage_inst_dmem_ram_1928, MEM_stage_inst_dmem_ram_1929, MEM_stage_inst_dmem_ram_1930, MEM_stage_inst_dmem_ram_1931, MEM_stage_inst_dmem_ram_1932, MEM_stage_inst_dmem_ram_1933, MEM_stage_inst_dmem_ram_1934, MEM_stage_inst_dmem_ram_1935, MEM_stage_inst_dmem_ram_1936, MEM_stage_inst_dmem_ram_1937, MEM_stage_inst_dmem_ram_1938, MEM_stage_inst_dmem_ram_1939, MEM_stage_inst_dmem_ram_1940, MEM_stage_inst_dmem_ram_1941, MEM_stage_inst_dmem_ram_1942, MEM_stage_inst_dmem_ram_1943, MEM_stage_inst_dmem_ram_1944, MEM_stage_inst_dmem_ram_1945, MEM_stage_inst_dmem_ram_1946, MEM_stage_inst_dmem_ram_1947, MEM_stage_inst_dmem_ram_1948, MEM_stage_inst_dmem_ram_1949, MEM_stage_inst_dmem_ram_1950, MEM_stage_inst_dmem_ram_1951, MEM_stage_inst_dmem_ram_1952, MEM_stage_inst_dmem_ram_1953, MEM_stage_inst_dmem_ram_1954, MEM_stage_inst_dmem_ram_1955, MEM_stage_inst_dmem_ram_1956, MEM_stage_inst_dmem_ram_1957, MEM_stage_inst_dmem_ram_1958, MEM_stage_inst_dmem_ram_1959, MEM_stage_inst_dmem_ram_1960, MEM_stage_inst_dmem_ram_1961, MEM_stage_inst_dmem_ram_1962, MEM_stage_inst_dmem_ram_1963, MEM_stage_inst_dmem_ram_1964, MEM_stage_inst_dmem_ram_1965, MEM_stage_inst_dmem_ram_1966, MEM_stage_inst_dmem_ram_1967, MEM_stage_inst_dmem_ram_1968, MEM_stage_inst_dmem_ram_1969, MEM_stage_inst_dmem_ram_1970, MEM_stage_inst_dmem_ram_1971, MEM_stage_inst_dmem_ram_1972, MEM_stage_inst_dmem_ram_1973, MEM_stage_inst_dmem_ram_1974, MEM_stage_inst_dmem_ram_1975, MEM_stage_inst_dmem_ram_1976, MEM_stage_inst_dmem_ram_1977, MEM_stage_inst_dmem_ram_1978, MEM_stage_inst_dmem_ram_1979, MEM_stage_inst_dmem_ram_1980, MEM_stage_inst_dmem_ram_1981, MEM_stage_inst_dmem_ram_1982, MEM_stage_inst_dmem_ram_1983, MEM_stage_inst_dmem_ram_1984, MEM_stage_inst_dmem_ram_1985, MEM_stage_inst_dmem_ram_1986, MEM_stage_inst_dmem_ram_1987, MEM_stage_inst_dmem_ram_1988, MEM_stage_inst_dmem_ram_1989, MEM_stage_inst_dmem_ram_1990, MEM_stage_inst_dmem_ram_1991, MEM_stage_inst_dmem_ram_1992, MEM_stage_inst_dmem_ram_1993, MEM_stage_inst_dmem_ram_1994, MEM_stage_inst_dmem_ram_1995, MEM_stage_inst_dmem_ram_1996, MEM_stage_inst_dmem_ram_1997, MEM_stage_inst_dmem_ram_1998, MEM_stage_inst_dmem_ram_1999, MEM_stage_inst_dmem_ram_2000, MEM_stage_inst_dmem_ram_2001, MEM_stage_inst_dmem_ram_2002, MEM_stage_inst_dmem_ram_2003, MEM_stage_inst_dmem_ram_2004, MEM_stage_inst_dmem_ram_2005, MEM_stage_inst_dmem_ram_2006, MEM_stage_inst_dmem_ram_2007, MEM_stage_inst_dmem_ram_2008, MEM_stage_inst_dmem_ram_2009, MEM_stage_inst_dmem_ram_2010, MEM_stage_inst_dmem_ram_2011, MEM_stage_inst_dmem_ram_2012, MEM_stage_inst_dmem_ram_2013, MEM_stage_inst_dmem_ram_2014, MEM_stage_inst_dmem_ram_2015, MEM_stage_inst_dmem_ram_2016, MEM_stage_inst_dmem_ram_2017, MEM_stage_inst_dmem_ram_2018, MEM_stage_inst_dmem_ram_2019, MEM_stage_inst_dmem_ram_2020, MEM_stage_inst_dmem_ram_2021, MEM_stage_inst_dmem_ram_2022, MEM_stage_inst_dmem_ram_2023, MEM_stage_inst_dmem_ram_2024, MEM_stage_inst_dmem_ram_2025, MEM_stage_inst_dmem_ram_2026, MEM_stage_inst_dmem_ram_2027, MEM_stage_inst_dmem_ram_2028, MEM_stage_inst_dmem_ram_2029, MEM_stage_inst_dmem_ram_2030, MEM_stage_inst_dmem_ram_2031, MEM_stage_inst_dmem_ram_2032, MEM_stage_inst_dmem_ram_2033, MEM_stage_inst_dmem_ram_2034, MEM_stage_inst_dmem_ram_2035, MEM_stage_inst_dmem_ram_2036, MEM_stage_inst_dmem_ram_2037, MEM_stage_inst_dmem_ram_2038, MEM_stage_inst_dmem_ram_2039, MEM_stage_inst_dmem_ram_2040, MEM_stage_inst_dmem_ram_2041, MEM_stage_inst_dmem_ram_2042, MEM_stage_inst_dmem_ram_2043, MEM_stage_inst_dmem_ram_2044, MEM_stage_inst_dmem_ram_2045, MEM_stage_inst_dmem_ram_2046, MEM_stage_inst_dmem_ram_2047, MEM_stage_inst_dmem_ram_1024, MEM_stage_inst_dmem_ram_1025, MEM_stage_inst_dmem_ram_1026, MEM_stage_inst_dmem_ram_1027, MEM_stage_inst_dmem_ram_1028, MEM_stage_inst_dmem_ram_1029, MEM_stage_inst_dmem_ram_1030, MEM_stage_inst_dmem_ram_1031, MEM_stage_inst_dmem_ram_1032, MEM_stage_inst_dmem_ram_1033, MEM_stage_inst_dmem_ram_1034, MEM_stage_inst_dmem_ram_1035, MEM_stage_inst_dmem_ram_1036, MEM_stage_inst_dmem_ram_1037, MEM_stage_inst_dmem_ram_1038, MEM_stage_inst_dmem_ram_1039, MEM_stage_inst_dmem_ram_1040, MEM_stage_inst_dmem_ram_1041, MEM_stage_inst_dmem_ram_1042, MEM_stage_inst_dmem_ram_1043, MEM_stage_inst_dmem_ram_1044, MEM_stage_inst_dmem_ram_1045, MEM_stage_inst_dmem_ram_1046, MEM_stage_inst_dmem_ram_1047, MEM_stage_inst_dmem_ram_1048, MEM_stage_inst_dmem_ram_1049, MEM_stage_inst_dmem_ram_1050, MEM_stage_inst_dmem_ram_1051, MEM_stage_inst_dmem_ram_1052, MEM_stage_inst_dmem_ram_1053, MEM_stage_inst_dmem_ram_1054, MEM_stage_inst_dmem_ram_1055, MEM_stage_inst_dmem_ram_1056, MEM_stage_inst_dmem_ram_1057, MEM_stage_inst_dmem_ram_1058, MEM_stage_inst_dmem_ram_1059, MEM_stage_inst_dmem_ram_1060, MEM_stage_inst_dmem_ram_1061, MEM_stage_inst_dmem_ram_1062, MEM_stage_inst_dmem_ram_1063, MEM_stage_inst_dmem_ram_1064, MEM_stage_inst_dmem_ram_1065, MEM_stage_inst_dmem_ram_1066, MEM_stage_inst_dmem_ram_1067, MEM_stage_inst_dmem_ram_1068, MEM_stage_inst_dmem_ram_1069, MEM_stage_inst_dmem_ram_1070, MEM_stage_inst_dmem_ram_1071, MEM_stage_inst_dmem_ram_1072, MEM_stage_inst_dmem_ram_1073, MEM_stage_inst_dmem_ram_1074, MEM_stage_inst_dmem_ram_1075, MEM_stage_inst_dmem_ram_1076, MEM_stage_inst_dmem_ram_1077, MEM_stage_inst_dmem_ram_1078, MEM_stage_inst_dmem_ram_1079, MEM_stage_inst_dmem_ram_1080, MEM_stage_inst_dmem_ram_1081, MEM_stage_inst_dmem_ram_1082, MEM_stage_inst_dmem_ram_1083, MEM_stage_inst_dmem_ram_1084, MEM_stage_inst_dmem_ram_1085, MEM_stage_inst_dmem_ram_1086, MEM_stage_inst_dmem_ram_1087, MEM_stage_inst_dmem_ram_1088, MEM_stage_inst_dmem_ram_1089, MEM_stage_inst_dmem_ram_1090, MEM_stage_inst_dmem_ram_1091, MEM_stage_inst_dmem_ram_1092, MEM_stage_inst_dmem_ram_1093, MEM_stage_inst_dmem_ram_1094, MEM_stage_inst_dmem_ram_1095, MEM_stage_inst_dmem_ram_1096, MEM_stage_inst_dmem_ram_1097, MEM_stage_inst_dmem_ram_1098, MEM_stage_inst_dmem_ram_1099, MEM_stage_inst_dmem_ram_1100, MEM_stage_inst_dmem_ram_1101, MEM_stage_inst_dmem_ram_1102, MEM_stage_inst_dmem_ram_1103, MEM_stage_inst_dmem_ram_1104, MEM_stage_inst_dmem_ram_1105, MEM_stage_inst_dmem_ram_1106, MEM_stage_inst_dmem_ram_1107, MEM_stage_inst_dmem_ram_1108, MEM_stage_inst_dmem_ram_1109, MEM_stage_inst_dmem_ram_1110, MEM_stage_inst_dmem_ram_1111, MEM_stage_inst_dmem_ram_1112, MEM_stage_inst_dmem_ram_1113, MEM_stage_inst_dmem_ram_1114, MEM_stage_inst_dmem_ram_1115, MEM_stage_inst_dmem_ram_1116, MEM_stage_inst_dmem_ram_1117, MEM_stage_inst_dmem_ram_1118, MEM_stage_inst_dmem_ram_1119, MEM_stage_inst_dmem_ram_1120, MEM_stage_inst_dmem_ram_1121, MEM_stage_inst_dmem_ram_1122, MEM_stage_inst_dmem_ram_1123, MEM_stage_inst_dmem_ram_1124, MEM_stage_inst_dmem_ram_1125, MEM_stage_inst_dmem_ram_1126, MEM_stage_inst_dmem_ram_1127, MEM_stage_inst_dmem_ram_1128, MEM_stage_inst_dmem_ram_1129, MEM_stage_inst_dmem_ram_1130, MEM_stage_inst_dmem_ram_1131, MEM_stage_inst_dmem_ram_1132, MEM_stage_inst_dmem_ram_1133, MEM_stage_inst_dmem_ram_1134, MEM_stage_inst_dmem_ram_1135, MEM_stage_inst_dmem_ram_1136, MEM_stage_inst_dmem_ram_1137, MEM_stage_inst_dmem_ram_1138, MEM_stage_inst_dmem_ram_1139, MEM_stage_inst_dmem_ram_1140, MEM_stage_inst_dmem_ram_1141, MEM_stage_inst_dmem_ram_1142, MEM_stage_inst_dmem_ram_1143, MEM_stage_inst_dmem_ram_1144, MEM_stage_inst_dmem_ram_1145, MEM_stage_inst_dmem_ram_1146, MEM_stage_inst_dmem_ram_1147, MEM_stage_inst_dmem_ram_1148, MEM_stage_inst_dmem_ram_1149, MEM_stage_inst_dmem_ram_1150, MEM_stage_inst_dmem_ram_1151, MEM_stage_inst_dmem_ram_1152, MEM_stage_inst_dmem_ram_1153, MEM_stage_inst_dmem_ram_1154, MEM_stage_inst_dmem_ram_1155, MEM_stage_inst_dmem_ram_1156, MEM_stage_inst_dmem_ram_1157, MEM_stage_inst_dmem_ram_1158, MEM_stage_inst_dmem_ram_1159, MEM_stage_inst_dmem_ram_1160, MEM_stage_inst_dmem_ram_1161, MEM_stage_inst_dmem_ram_1162, MEM_stage_inst_dmem_ram_1163, MEM_stage_inst_dmem_ram_1164, MEM_stage_inst_dmem_ram_1165, MEM_stage_inst_dmem_ram_1166, MEM_stage_inst_dmem_ram_1167, MEM_stage_inst_dmem_ram_1168, MEM_stage_inst_dmem_ram_1169, MEM_stage_inst_dmem_ram_1170, MEM_stage_inst_dmem_ram_1171, MEM_stage_inst_dmem_ram_1172, MEM_stage_inst_dmem_ram_1173, MEM_stage_inst_dmem_ram_1174, MEM_stage_inst_dmem_ram_1175, MEM_stage_inst_dmem_ram_1176, MEM_stage_inst_dmem_ram_1177, MEM_stage_inst_dmem_ram_1178, MEM_stage_inst_dmem_ram_1179, MEM_stage_inst_dmem_ram_1180, MEM_stage_inst_dmem_ram_1181, MEM_stage_inst_dmem_ram_1182, MEM_stage_inst_dmem_ram_1183, MEM_stage_inst_dmem_ram_1184, MEM_stage_inst_dmem_ram_1185, MEM_stage_inst_dmem_ram_1186, MEM_stage_inst_dmem_ram_1187, MEM_stage_inst_dmem_ram_1188, MEM_stage_inst_dmem_ram_1189, MEM_stage_inst_dmem_ram_1190, MEM_stage_inst_dmem_ram_1191, MEM_stage_inst_dmem_ram_1192, MEM_stage_inst_dmem_ram_1193, MEM_stage_inst_dmem_ram_1194, MEM_stage_inst_dmem_ram_1195, MEM_stage_inst_dmem_ram_1196, MEM_stage_inst_dmem_ram_1197, MEM_stage_inst_dmem_ram_1198, MEM_stage_inst_dmem_ram_1199, MEM_stage_inst_dmem_ram_1200, MEM_stage_inst_dmem_ram_1201, MEM_stage_inst_dmem_ram_1202, MEM_stage_inst_dmem_ram_1203, MEM_stage_inst_dmem_ram_1204, MEM_stage_inst_dmem_ram_1205, MEM_stage_inst_dmem_ram_1206, MEM_stage_inst_dmem_ram_1207, MEM_stage_inst_dmem_ram_1208, MEM_stage_inst_dmem_ram_1209, MEM_stage_inst_dmem_ram_1210, MEM_stage_inst_dmem_ram_1211, MEM_stage_inst_dmem_ram_1212, MEM_stage_inst_dmem_ram_1213, MEM_stage_inst_dmem_ram_1214, MEM_stage_inst_dmem_ram_1215, MEM_stage_inst_dmem_ram_1216, MEM_stage_inst_dmem_ram_1217, MEM_stage_inst_dmem_ram_1218, MEM_stage_inst_dmem_ram_1219, MEM_stage_inst_dmem_ram_1220, MEM_stage_inst_dmem_ram_1221, MEM_stage_inst_dmem_ram_1222, MEM_stage_inst_dmem_ram_1223, MEM_stage_inst_dmem_ram_1224, MEM_stage_inst_dmem_ram_1225, MEM_stage_inst_dmem_ram_1226, MEM_stage_inst_dmem_ram_1227, MEM_stage_inst_dmem_ram_1228, MEM_stage_inst_dmem_ram_1229, MEM_stage_inst_dmem_ram_1230, MEM_stage_inst_dmem_ram_1231, MEM_stage_inst_dmem_ram_1232, MEM_stage_inst_dmem_ram_1233, MEM_stage_inst_dmem_ram_1234, MEM_stage_inst_dmem_ram_1235, MEM_stage_inst_dmem_ram_1236, MEM_stage_inst_dmem_ram_1237, MEM_stage_inst_dmem_ram_1238, MEM_stage_inst_dmem_ram_1239, MEM_stage_inst_dmem_ram_1240, MEM_stage_inst_dmem_ram_1241, MEM_stage_inst_dmem_ram_1242, MEM_stage_inst_dmem_ram_1243, MEM_stage_inst_dmem_ram_1244, MEM_stage_inst_dmem_ram_1245, MEM_stage_inst_dmem_ram_1246, MEM_stage_inst_dmem_ram_1247, MEM_stage_inst_dmem_ram_1248, MEM_stage_inst_dmem_ram_1249, MEM_stage_inst_dmem_ram_1250, MEM_stage_inst_dmem_ram_1251, MEM_stage_inst_dmem_ram_1252, MEM_stage_inst_dmem_ram_1253, MEM_stage_inst_dmem_ram_1254, MEM_stage_inst_dmem_ram_1255, MEM_stage_inst_dmem_ram_1256, MEM_stage_inst_dmem_ram_1257, MEM_stage_inst_dmem_ram_1258, MEM_stage_inst_dmem_ram_1259, MEM_stage_inst_dmem_ram_1260, MEM_stage_inst_dmem_ram_1261, MEM_stage_inst_dmem_ram_1262, MEM_stage_inst_dmem_ram_1263, MEM_stage_inst_dmem_ram_1264, MEM_stage_inst_dmem_ram_1265, MEM_stage_inst_dmem_ram_1266, MEM_stage_inst_dmem_ram_1267, MEM_stage_inst_dmem_ram_1268, MEM_stage_inst_dmem_ram_1269, MEM_stage_inst_dmem_ram_1270, MEM_stage_inst_dmem_ram_1271, MEM_stage_inst_dmem_ram_1272, MEM_stage_inst_dmem_ram_1273, MEM_stage_inst_dmem_ram_1274, MEM_stage_inst_dmem_ram_1275, MEM_stage_inst_dmem_ram_1276, MEM_stage_inst_dmem_ram_1277, MEM_stage_inst_dmem_ram_1278, MEM_stage_inst_dmem_ram_1279, MEM_stage_inst_dmem_ram_1280, MEM_stage_inst_dmem_ram_1281, MEM_stage_inst_dmem_ram_1282, MEM_stage_inst_dmem_ram_1283, MEM_stage_inst_dmem_ram_1284, MEM_stage_inst_dmem_ram_1285, MEM_stage_inst_dmem_ram_1286, MEM_stage_inst_dmem_ram_1287, MEM_stage_inst_dmem_ram_1288, MEM_stage_inst_dmem_ram_1289, MEM_stage_inst_dmem_ram_1290, MEM_stage_inst_dmem_ram_1291, MEM_stage_inst_dmem_ram_1292, MEM_stage_inst_dmem_ram_1293, MEM_stage_inst_dmem_ram_1294, MEM_stage_inst_dmem_ram_1295, MEM_stage_inst_dmem_ram_1296, MEM_stage_inst_dmem_ram_1297, MEM_stage_inst_dmem_ram_1298, MEM_stage_inst_dmem_ram_1299, MEM_stage_inst_dmem_ram_1300, MEM_stage_inst_dmem_ram_1301, MEM_stage_inst_dmem_ram_1302, MEM_stage_inst_dmem_ram_1303, MEM_stage_inst_dmem_ram_1304, MEM_stage_inst_dmem_ram_1305, MEM_stage_inst_dmem_ram_1306, MEM_stage_inst_dmem_ram_1307, MEM_stage_inst_dmem_ram_1308, MEM_stage_inst_dmem_ram_1309, MEM_stage_inst_dmem_ram_1310, MEM_stage_inst_dmem_ram_1311, MEM_stage_inst_dmem_ram_1312, MEM_stage_inst_dmem_ram_1313, MEM_stage_inst_dmem_ram_1314, MEM_stage_inst_dmem_ram_1315, MEM_stage_inst_dmem_ram_1316, MEM_stage_inst_dmem_ram_1317, MEM_stage_inst_dmem_ram_1318, MEM_stage_inst_dmem_ram_1319, MEM_stage_inst_dmem_ram_1320, MEM_stage_inst_dmem_ram_1321, MEM_stage_inst_dmem_ram_1322, MEM_stage_inst_dmem_ram_1323, MEM_stage_inst_dmem_ram_1324, MEM_stage_inst_dmem_ram_1325, MEM_stage_inst_dmem_ram_1326, MEM_stage_inst_dmem_ram_1327, MEM_stage_inst_dmem_ram_1328, MEM_stage_inst_dmem_ram_1329, MEM_stage_inst_dmem_ram_1330, MEM_stage_inst_dmem_ram_1331, MEM_stage_inst_dmem_ram_1332, MEM_stage_inst_dmem_ram_1333, MEM_stage_inst_dmem_ram_1334, MEM_stage_inst_dmem_ram_1335, MEM_stage_inst_dmem_ram_1336, MEM_stage_inst_dmem_ram_1337, MEM_stage_inst_dmem_ram_1338, MEM_stage_inst_dmem_ram_1339, MEM_stage_inst_dmem_ram_1340, MEM_stage_inst_dmem_ram_1341, MEM_stage_inst_dmem_ram_1342, MEM_stage_inst_dmem_ram_1343, MEM_stage_inst_dmem_ram_1344, MEM_stage_inst_dmem_ram_1345, MEM_stage_inst_dmem_ram_1346, MEM_stage_inst_dmem_ram_1347, MEM_stage_inst_dmem_ram_1348, MEM_stage_inst_dmem_ram_1349, MEM_stage_inst_dmem_ram_1350, MEM_stage_inst_dmem_ram_1351, MEM_stage_inst_dmem_ram_1352, MEM_stage_inst_dmem_ram_1353, MEM_stage_inst_dmem_ram_1354, MEM_stage_inst_dmem_ram_1355, MEM_stage_inst_dmem_ram_1356, MEM_stage_inst_dmem_ram_1357, MEM_stage_inst_dmem_ram_1358, MEM_stage_inst_dmem_ram_1359, MEM_stage_inst_dmem_ram_1360, MEM_stage_inst_dmem_ram_1361, MEM_stage_inst_dmem_ram_1362, MEM_stage_inst_dmem_ram_1363, MEM_stage_inst_dmem_ram_1364, MEM_stage_inst_dmem_ram_1365, MEM_stage_inst_dmem_ram_1366, MEM_stage_inst_dmem_ram_1367, MEM_stage_inst_dmem_ram_1368, MEM_stage_inst_dmem_ram_1369, MEM_stage_inst_dmem_ram_1370, MEM_stage_inst_dmem_ram_1371, MEM_stage_inst_dmem_ram_1372, MEM_stage_inst_dmem_ram_1373, MEM_stage_inst_dmem_ram_1374, MEM_stage_inst_dmem_ram_1375, MEM_stage_inst_dmem_ram_1376, MEM_stage_inst_dmem_ram_1377, MEM_stage_inst_dmem_ram_1378, MEM_stage_inst_dmem_ram_1379, MEM_stage_inst_dmem_ram_1380, MEM_stage_inst_dmem_ram_1381, MEM_stage_inst_dmem_ram_1382, MEM_stage_inst_dmem_ram_1383, MEM_stage_inst_dmem_ram_1384, MEM_stage_inst_dmem_ram_1385, MEM_stage_inst_dmem_ram_1386, MEM_stage_inst_dmem_ram_1387, MEM_stage_inst_dmem_ram_1388, MEM_stage_inst_dmem_ram_1389, MEM_stage_inst_dmem_ram_1390, MEM_stage_inst_dmem_ram_1391, MEM_stage_inst_dmem_ram_1392, MEM_stage_inst_dmem_ram_1393, MEM_stage_inst_dmem_ram_1394, MEM_stage_inst_dmem_ram_1395, MEM_stage_inst_dmem_ram_1396, MEM_stage_inst_dmem_ram_1397, MEM_stage_inst_dmem_ram_1398, MEM_stage_inst_dmem_ram_1399, MEM_stage_inst_dmem_ram_1400, MEM_stage_inst_dmem_ram_1401, MEM_stage_inst_dmem_ram_1402, MEM_stage_inst_dmem_ram_1403, MEM_stage_inst_dmem_ram_1404, MEM_stage_inst_dmem_ram_1405, MEM_stage_inst_dmem_ram_1406, MEM_stage_inst_dmem_ram_1407, MEM_stage_inst_dmem_ram_1408, MEM_stage_inst_dmem_ram_1409, MEM_stage_inst_dmem_ram_1410, MEM_stage_inst_dmem_ram_1411, MEM_stage_inst_dmem_ram_1412, MEM_stage_inst_dmem_ram_1413, MEM_stage_inst_dmem_ram_1414, MEM_stage_inst_dmem_ram_1415, MEM_stage_inst_dmem_ram_1416, MEM_stage_inst_dmem_ram_1417, MEM_stage_inst_dmem_ram_1418, MEM_stage_inst_dmem_ram_1419, MEM_stage_inst_dmem_ram_1420, MEM_stage_inst_dmem_ram_1421, MEM_stage_inst_dmem_ram_1422, MEM_stage_inst_dmem_ram_1423, MEM_stage_inst_dmem_ram_1424, MEM_stage_inst_dmem_ram_1425, MEM_stage_inst_dmem_ram_1426, MEM_stage_inst_dmem_ram_1427, MEM_stage_inst_dmem_ram_1428, MEM_stage_inst_dmem_ram_1429, MEM_stage_inst_dmem_ram_1430, MEM_stage_inst_dmem_ram_1431, MEM_stage_inst_dmem_ram_1432, MEM_stage_inst_dmem_ram_1433, MEM_stage_inst_dmem_ram_1434, MEM_stage_inst_dmem_ram_1435, MEM_stage_inst_dmem_ram_1436, MEM_stage_inst_dmem_ram_1437, MEM_stage_inst_dmem_ram_1438, MEM_stage_inst_dmem_ram_1439, MEM_stage_inst_dmem_ram_1440, MEM_stage_inst_dmem_ram_1441, MEM_stage_inst_dmem_ram_1442, MEM_stage_inst_dmem_ram_1443, MEM_stage_inst_dmem_ram_1444, MEM_stage_inst_dmem_ram_1445, MEM_stage_inst_dmem_ram_1446, MEM_stage_inst_dmem_ram_1447, MEM_stage_inst_dmem_ram_1448, MEM_stage_inst_dmem_ram_1449, MEM_stage_inst_dmem_ram_1450, MEM_stage_inst_dmem_ram_1451, MEM_stage_inst_dmem_ram_1452, MEM_stage_inst_dmem_ram_1453, MEM_stage_inst_dmem_ram_1454, MEM_stage_inst_dmem_ram_1455, MEM_stage_inst_dmem_ram_1456, MEM_stage_inst_dmem_ram_1457, MEM_stage_inst_dmem_ram_1458, MEM_stage_inst_dmem_ram_1459, MEM_stage_inst_dmem_ram_1460, MEM_stage_inst_dmem_ram_1461, MEM_stage_inst_dmem_ram_1462, MEM_stage_inst_dmem_ram_1463, MEM_stage_inst_dmem_ram_1464, MEM_stage_inst_dmem_ram_1465, MEM_stage_inst_dmem_ram_1466, MEM_stage_inst_dmem_ram_1467, MEM_stage_inst_dmem_ram_1468, MEM_stage_inst_dmem_ram_1469, MEM_stage_inst_dmem_ram_1470, MEM_stage_inst_dmem_ram_1471, MEM_stage_inst_dmem_ram_1472, MEM_stage_inst_dmem_ram_1473, MEM_stage_inst_dmem_ram_1474, MEM_stage_inst_dmem_ram_1475, MEM_stage_inst_dmem_ram_1476, MEM_stage_inst_dmem_ram_1477, MEM_stage_inst_dmem_ram_1478, MEM_stage_inst_dmem_ram_1479, MEM_stage_inst_dmem_ram_1480, MEM_stage_inst_dmem_ram_1481, MEM_stage_inst_dmem_ram_1482, MEM_stage_inst_dmem_ram_1483, MEM_stage_inst_dmem_ram_1484, MEM_stage_inst_dmem_ram_1485, MEM_stage_inst_dmem_ram_1486, MEM_stage_inst_dmem_ram_1487, MEM_stage_inst_dmem_ram_1488, MEM_stage_inst_dmem_ram_1489, MEM_stage_inst_dmem_ram_1490, MEM_stage_inst_dmem_ram_1491, MEM_stage_inst_dmem_ram_1492, MEM_stage_inst_dmem_ram_1493, MEM_stage_inst_dmem_ram_1494, MEM_stage_inst_dmem_ram_1495, MEM_stage_inst_dmem_ram_1496, MEM_stage_inst_dmem_ram_1497, MEM_stage_inst_dmem_ram_1498, MEM_stage_inst_dmem_ram_1499, MEM_stage_inst_dmem_ram_1500, MEM_stage_inst_dmem_ram_1501, MEM_stage_inst_dmem_ram_1502, MEM_stage_inst_dmem_ram_1503, MEM_stage_inst_dmem_ram_1504, MEM_stage_inst_dmem_ram_1505, MEM_stage_inst_dmem_ram_1506, MEM_stage_inst_dmem_ram_1507, MEM_stage_inst_dmem_ram_1508, MEM_stage_inst_dmem_ram_1509, MEM_stage_inst_dmem_ram_1510, MEM_stage_inst_dmem_ram_1511, MEM_stage_inst_dmem_ram_1512, MEM_stage_inst_dmem_ram_1513, MEM_stage_inst_dmem_ram_1514, MEM_stage_inst_dmem_ram_1515, MEM_stage_inst_dmem_ram_1516, MEM_stage_inst_dmem_ram_1517, MEM_stage_inst_dmem_ram_1518, MEM_stage_inst_dmem_ram_1519, MEM_stage_inst_dmem_ram_1520, MEM_stage_inst_dmem_ram_1521, MEM_stage_inst_dmem_ram_1522, MEM_stage_inst_dmem_ram_1523, MEM_stage_inst_dmem_ram_1524, MEM_stage_inst_dmem_ram_1525, MEM_stage_inst_dmem_ram_1526, MEM_stage_inst_dmem_ram_1527, MEM_stage_inst_dmem_ram_1528, MEM_stage_inst_dmem_ram_1529, MEM_stage_inst_dmem_ram_1530, MEM_stage_inst_dmem_ram_1531, MEM_stage_inst_dmem_ram_1532, MEM_stage_inst_dmem_ram_1533, MEM_stage_inst_dmem_ram_1534, MEM_stage_inst_dmem_ram_1535, MEM_stage_inst_dmem_ram_512, MEM_stage_inst_dmem_ram_513, MEM_stage_inst_dmem_ram_514, MEM_stage_inst_dmem_ram_515, MEM_stage_inst_dmem_ram_516, MEM_stage_inst_dmem_ram_517, MEM_stage_inst_dmem_ram_518, MEM_stage_inst_dmem_ram_519, MEM_stage_inst_dmem_ram_520, MEM_stage_inst_dmem_ram_521, MEM_stage_inst_dmem_ram_522, MEM_stage_inst_dmem_ram_523, MEM_stage_inst_dmem_ram_524, MEM_stage_inst_dmem_ram_525, MEM_stage_inst_dmem_ram_526, MEM_stage_inst_dmem_ram_527, MEM_stage_inst_dmem_ram_528, MEM_stage_inst_dmem_ram_529, MEM_stage_inst_dmem_ram_530, MEM_stage_inst_dmem_ram_531, MEM_stage_inst_dmem_ram_532, MEM_stage_inst_dmem_ram_533, MEM_stage_inst_dmem_ram_534, MEM_stage_inst_dmem_ram_535, MEM_stage_inst_dmem_ram_536, MEM_stage_inst_dmem_ram_537, MEM_stage_inst_dmem_ram_538, MEM_stage_inst_dmem_ram_539, MEM_stage_inst_dmem_ram_540, MEM_stage_inst_dmem_ram_541, MEM_stage_inst_dmem_ram_542, MEM_stage_inst_dmem_ram_543, MEM_stage_inst_dmem_ram_544, MEM_stage_inst_dmem_ram_545, MEM_stage_inst_dmem_ram_546, MEM_stage_inst_dmem_ram_547, MEM_stage_inst_dmem_ram_548, MEM_stage_inst_dmem_ram_549, MEM_stage_inst_dmem_ram_550, MEM_stage_inst_dmem_ram_551, MEM_stage_inst_dmem_ram_552, MEM_stage_inst_dmem_ram_553, MEM_stage_inst_dmem_ram_554, MEM_stage_inst_dmem_ram_555, MEM_stage_inst_dmem_ram_556, MEM_stage_inst_dmem_ram_557, MEM_stage_inst_dmem_ram_558, MEM_stage_inst_dmem_ram_559, MEM_stage_inst_dmem_ram_560, MEM_stage_inst_dmem_ram_561, MEM_stage_inst_dmem_ram_562, MEM_stage_inst_dmem_ram_563, MEM_stage_inst_dmem_ram_564, MEM_stage_inst_dmem_ram_565, MEM_stage_inst_dmem_ram_566, MEM_stage_inst_dmem_ram_567, MEM_stage_inst_dmem_ram_568, MEM_stage_inst_dmem_ram_569, MEM_stage_inst_dmem_ram_570, MEM_stage_inst_dmem_ram_571, MEM_stage_inst_dmem_ram_572, MEM_stage_inst_dmem_ram_573, MEM_stage_inst_dmem_ram_574, MEM_stage_inst_dmem_ram_575, MEM_stage_inst_dmem_ram_576, MEM_stage_inst_dmem_ram_577, MEM_stage_inst_dmem_ram_578, MEM_stage_inst_dmem_ram_579, MEM_stage_inst_dmem_ram_580, MEM_stage_inst_dmem_ram_581, MEM_stage_inst_dmem_ram_582, MEM_stage_inst_dmem_ram_583, MEM_stage_inst_dmem_ram_584, MEM_stage_inst_dmem_ram_585, MEM_stage_inst_dmem_ram_586, MEM_stage_inst_dmem_ram_587, MEM_stage_inst_dmem_ram_588, MEM_stage_inst_dmem_ram_589, MEM_stage_inst_dmem_ram_590, MEM_stage_inst_dmem_ram_591, MEM_stage_inst_dmem_ram_592, MEM_stage_inst_dmem_ram_593, MEM_stage_inst_dmem_ram_594, MEM_stage_inst_dmem_ram_595, MEM_stage_inst_dmem_ram_596, MEM_stage_inst_dmem_ram_597, MEM_stage_inst_dmem_ram_598, MEM_stage_inst_dmem_ram_599, MEM_stage_inst_dmem_ram_600, MEM_stage_inst_dmem_ram_601, MEM_stage_inst_dmem_ram_602, MEM_stage_inst_dmem_ram_603, MEM_stage_inst_dmem_ram_604, MEM_stage_inst_dmem_ram_605, MEM_stage_inst_dmem_ram_606, MEM_stage_inst_dmem_ram_607, MEM_stage_inst_dmem_ram_608, MEM_stage_inst_dmem_ram_609, MEM_stage_inst_dmem_ram_610, MEM_stage_inst_dmem_ram_611, MEM_stage_inst_dmem_ram_612, MEM_stage_inst_dmem_ram_613, MEM_stage_inst_dmem_ram_614, MEM_stage_inst_dmem_ram_615, MEM_stage_inst_dmem_ram_616, MEM_stage_inst_dmem_ram_617, MEM_stage_inst_dmem_ram_618, MEM_stage_inst_dmem_ram_619, MEM_stage_inst_dmem_ram_620, MEM_stage_inst_dmem_ram_621, MEM_stage_inst_dmem_ram_622, MEM_stage_inst_dmem_ram_623, MEM_stage_inst_dmem_ram_624, MEM_stage_inst_dmem_ram_625, MEM_stage_inst_dmem_ram_626, MEM_stage_inst_dmem_ram_627, MEM_stage_inst_dmem_ram_628, MEM_stage_inst_dmem_ram_629, MEM_stage_inst_dmem_ram_630, MEM_stage_inst_dmem_ram_631, MEM_stage_inst_dmem_ram_632, MEM_stage_inst_dmem_ram_633, MEM_stage_inst_dmem_ram_634, MEM_stage_inst_dmem_ram_635, MEM_stage_inst_dmem_ram_636, MEM_stage_inst_dmem_ram_637, MEM_stage_inst_dmem_ram_638, MEM_stage_inst_dmem_ram_639, MEM_stage_inst_dmem_ram_640, MEM_stage_inst_dmem_ram_641, MEM_stage_inst_dmem_ram_642, MEM_stage_inst_dmem_ram_643, MEM_stage_inst_dmem_ram_644, MEM_stage_inst_dmem_ram_645, MEM_stage_inst_dmem_ram_646, MEM_stage_inst_dmem_ram_647, MEM_stage_inst_dmem_ram_648, MEM_stage_inst_dmem_ram_649, MEM_stage_inst_dmem_ram_650, MEM_stage_inst_dmem_ram_651, MEM_stage_inst_dmem_ram_652, MEM_stage_inst_dmem_ram_653, MEM_stage_inst_dmem_ram_654, MEM_stage_inst_dmem_ram_655, MEM_stage_inst_dmem_ram_656, MEM_stage_inst_dmem_ram_657, MEM_stage_inst_dmem_ram_658, MEM_stage_inst_dmem_ram_659, MEM_stage_inst_dmem_ram_660, MEM_stage_inst_dmem_ram_661, MEM_stage_inst_dmem_ram_662, MEM_stage_inst_dmem_ram_663, MEM_stage_inst_dmem_ram_664, MEM_stage_inst_dmem_ram_665, MEM_stage_inst_dmem_ram_666, MEM_stage_inst_dmem_ram_667, MEM_stage_inst_dmem_ram_668, MEM_stage_inst_dmem_ram_669, MEM_stage_inst_dmem_ram_670, MEM_stage_inst_dmem_ram_671, MEM_stage_inst_dmem_ram_672, MEM_stage_inst_dmem_ram_673, MEM_stage_inst_dmem_ram_674, MEM_stage_inst_dmem_ram_675, MEM_stage_inst_dmem_ram_676, MEM_stage_inst_dmem_ram_677, MEM_stage_inst_dmem_ram_678, MEM_stage_inst_dmem_ram_679, MEM_stage_inst_dmem_ram_680, MEM_stage_inst_dmem_ram_681, MEM_stage_inst_dmem_ram_682, MEM_stage_inst_dmem_ram_683, MEM_stage_inst_dmem_ram_684, MEM_stage_inst_dmem_ram_685, MEM_stage_inst_dmem_ram_686, MEM_stage_inst_dmem_ram_687, MEM_stage_inst_dmem_ram_688, MEM_stage_inst_dmem_ram_689, MEM_stage_inst_dmem_ram_690, MEM_stage_inst_dmem_ram_691, MEM_stage_inst_dmem_ram_692, MEM_stage_inst_dmem_ram_693, MEM_stage_inst_dmem_ram_694, MEM_stage_inst_dmem_ram_695, MEM_stage_inst_dmem_ram_696, MEM_stage_inst_dmem_ram_697, MEM_stage_inst_dmem_ram_698, MEM_stage_inst_dmem_ram_699, MEM_stage_inst_dmem_ram_700, MEM_stage_inst_dmem_ram_701, MEM_stage_inst_dmem_ram_702, MEM_stage_inst_dmem_ram_703, MEM_stage_inst_dmem_ram_704, MEM_stage_inst_dmem_ram_705, MEM_stage_inst_dmem_ram_706, MEM_stage_inst_dmem_ram_707, MEM_stage_inst_dmem_ram_708, MEM_stage_inst_dmem_ram_709, MEM_stage_inst_dmem_ram_710, MEM_stage_inst_dmem_ram_711, MEM_stage_inst_dmem_ram_712, MEM_stage_inst_dmem_ram_713, MEM_stage_inst_dmem_ram_714, MEM_stage_inst_dmem_ram_715, MEM_stage_inst_dmem_ram_716, MEM_stage_inst_dmem_ram_717, MEM_stage_inst_dmem_ram_718, MEM_stage_inst_dmem_ram_719, MEM_stage_inst_dmem_ram_720, MEM_stage_inst_dmem_ram_721, MEM_stage_inst_dmem_ram_722, MEM_stage_inst_dmem_ram_723, MEM_stage_inst_dmem_ram_724, MEM_stage_inst_dmem_ram_725, MEM_stage_inst_dmem_ram_726, MEM_stage_inst_dmem_ram_727, MEM_stage_inst_dmem_ram_728, MEM_stage_inst_dmem_ram_729, MEM_stage_inst_dmem_ram_730, MEM_stage_inst_dmem_ram_731, MEM_stage_inst_dmem_ram_732, MEM_stage_inst_dmem_ram_733, MEM_stage_inst_dmem_ram_734, MEM_stage_inst_dmem_ram_735, MEM_stage_inst_dmem_ram_736, MEM_stage_inst_dmem_ram_737, MEM_stage_inst_dmem_ram_738, MEM_stage_inst_dmem_ram_739, MEM_stage_inst_dmem_ram_740, MEM_stage_inst_dmem_ram_741, MEM_stage_inst_dmem_ram_742, MEM_stage_inst_dmem_ram_743, MEM_stage_inst_dmem_ram_744, MEM_stage_inst_dmem_ram_745, MEM_stage_inst_dmem_ram_746, MEM_stage_inst_dmem_ram_747, MEM_stage_inst_dmem_ram_748, MEM_stage_inst_dmem_ram_749, MEM_stage_inst_dmem_ram_750, MEM_stage_inst_dmem_ram_751, MEM_stage_inst_dmem_ram_752, MEM_stage_inst_dmem_ram_753, MEM_stage_inst_dmem_ram_754, MEM_stage_inst_dmem_ram_755, MEM_stage_inst_dmem_ram_756, MEM_stage_inst_dmem_ram_757, MEM_stage_inst_dmem_ram_758, MEM_stage_inst_dmem_ram_759, MEM_stage_inst_dmem_ram_760, MEM_stage_inst_dmem_ram_761, MEM_stage_inst_dmem_ram_762, MEM_stage_inst_dmem_ram_763, MEM_stage_inst_dmem_ram_764, MEM_stage_inst_dmem_ram_765, MEM_stage_inst_dmem_ram_766, MEM_stage_inst_dmem_ram_767, MEM_stage_inst_dmem_ram_768, MEM_stage_inst_dmem_ram_769, MEM_stage_inst_dmem_ram_770, MEM_stage_inst_dmem_ram_771, MEM_stage_inst_dmem_ram_772, MEM_stage_inst_dmem_ram_773, MEM_stage_inst_dmem_ram_774, MEM_stage_inst_dmem_ram_775, MEM_stage_inst_dmem_ram_776, MEM_stage_inst_dmem_ram_777, MEM_stage_inst_dmem_ram_778, MEM_stage_inst_dmem_ram_779, MEM_stage_inst_dmem_ram_780, MEM_stage_inst_dmem_ram_781, MEM_stage_inst_dmem_ram_782, MEM_stage_inst_dmem_ram_783, MEM_stage_inst_dmem_ram_784, MEM_stage_inst_dmem_ram_785, MEM_stage_inst_dmem_ram_786, MEM_stage_inst_dmem_ram_787, MEM_stage_inst_dmem_ram_788, MEM_stage_inst_dmem_ram_789, MEM_stage_inst_dmem_ram_790, MEM_stage_inst_dmem_ram_791, MEM_stage_inst_dmem_ram_792, MEM_stage_inst_dmem_ram_793, MEM_stage_inst_dmem_ram_794, MEM_stage_inst_dmem_ram_795, MEM_stage_inst_dmem_ram_796, MEM_stage_inst_dmem_ram_797, MEM_stage_inst_dmem_ram_798, MEM_stage_inst_dmem_ram_799, MEM_stage_inst_dmem_ram_800, MEM_stage_inst_dmem_ram_801, MEM_stage_inst_dmem_ram_802, MEM_stage_inst_dmem_ram_803, MEM_stage_inst_dmem_ram_804, MEM_stage_inst_dmem_ram_805, MEM_stage_inst_dmem_ram_806, MEM_stage_inst_dmem_ram_807, MEM_stage_inst_dmem_ram_808, MEM_stage_inst_dmem_ram_809, MEM_stage_inst_dmem_ram_810, MEM_stage_inst_dmem_ram_811, MEM_stage_inst_dmem_ram_812, MEM_stage_inst_dmem_ram_813, MEM_stage_inst_dmem_ram_814, MEM_stage_inst_dmem_ram_815, MEM_stage_inst_dmem_ram_816, MEM_stage_inst_dmem_ram_817, MEM_stage_inst_dmem_ram_818, MEM_stage_inst_dmem_ram_819, MEM_stage_inst_dmem_ram_820, MEM_stage_inst_dmem_ram_821, MEM_stage_inst_dmem_ram_822, MEM_stage_inst_dmem_ram_823, MEM_stage_inst_dmem_ram_824, MEM_stage_inst_dmem_ram_825, MEM_stage_inst_dmem_ram_826, MEM_stage_inst_dmem_ram_827, MEM_stage_inst_dmem_ram_828, MEM_stage_inst_dmem_ram_829, MEM_stage_inst_dmem_ram_830, MEM_stage_inst_dmem_ram_831, MEM_stage_inst_dmem_ram_832, MEM_stage_inst_dmem_ram_833, MEM_stage_inst_dmem_ram_834, MEM_stage_inst_dmem_ram_835, MEM_stage_inst_dmem_ram_836, MEM_stage_inst_dmem_ram_837, MEM_stage_inst_dmem_ram_838, MEM_stage_inst_dmem_ram_839, MEM_stage_inst_dmem_ram_840, MEM_stage_inst_dmem_ram_841, MEM_stage_inst_dmem_ram_842, MEM_stage_inst_dmem_ram_843, MEM_stage_inst_dmem_ram_844, MEM_stage_inst_dmem_ram_845, MEM_stage_inst_dmem_ram_846, MEM_stage_inst_dmem_ram_847, MEM_stage_inst_dmem_ram_848, MEM_stage_inst_dmem_ram_849, MEM_stage_inst_dmem_ram_850, MEM_stage_inst_dmem_ram_851, MEM_stage_inst_dmem_ram_852, MEM_stage_inst_dmem_ram_853, MEM_stage_inst_dmem_ram_854, MEM_stage_inst_dmem_ram_855, MEM_stage_inst_dmem_ram_856, MEM_stage_inst_dmem_ram_857, MEM_stage_inst_dmem_ram_858, MEM_stage_inst_dmem_ram_859, MEM_stage_inst_dmem_ram_860, MEM_stage_inst_dmem_ram_861, MEM_stage_inst_dmem_ram_862, MEM_stage_inst_dmem_ram_863, MEM_stage_inst_dmem_ram_864, MEM_stage_inst_dmem_ram_865, MEM_stage_inst_dmem_ram_866, MEM_stage_inst_dmem_ram_867, MEM_stage_inst_dmem_ram_868, MEM_stage_inst_dmem_ram_869, MEM_stage_inst_dmem_ram_870, MEM_stage_inst_dmem_ram_871, MEM_stage_inst_dmem_ram_872, MEM_stage_inst_dmem_ram_873, MEM_stage_inst_dmem_ram_874, MEM_stage_inst_dmem_ram_875, MEM_stage_inst_dmem_ram_876, MEM_stage_inst_dmem_ram_877, MEM_stage_inst_dmem_ram_878, MEM_stage_inst_dmem_ram_879, MEM_stage_inst_dmem_ram_880, MEM_stage_inst_dmem_ram_881, MEM_stage_inst_dmem_ram_882, MEM_stage_inst_dmem_ram_883, MEM_stage_inst_dmem_ram_884, MEM_stage_inst_dmem_ram_885, MEM_stage_inst_dmem_ram_886, MEM_stage_inst_dmem_ram_887, MEM_stage_inst_dmem_ram_888, MEM_stage_inst_dmem_ram_889, MEM_stage_inst_dmem_ram_890, MEM_stage_inst_dmem_ram_891, MEM_stage_inst_dmem_ram_892, MEM_stage_inst_dmem_ram_893, MEM_stage_inst_dmem_ram_894, MEM_stage_inst_dmem_ram_895, MEM_stage_inst_dmem_ram_896, MEM_stage_inst_dmem_ram_897, MEM_stage_inst_dmem_ram_898, MEM_stage_inst_dmem_ram_899, MEM_stage_inst_dmem_ram_900, MEM_stage_inst_dmem_ram_901, MEM_stage_inst_dmem_ram_902, MEM_stage_inst_dmem_ram_903, MEM_stage_inst_dmem_ram_904, MEM_stage_inst_dmem_ram_905, MEM_stage_inst_dmem_ram_906, MEM_stage_inst_dmem_ram_907, MEM_stage_inst_dmem_ram_908, MEM_stage_inst_dmem_ram_909, MEM_stage_inst_dmem_ram_910, MEM_stage_inst_dmem_ram_911, MEM_stage_inst_dmem_ram_912, MEM_stage_inst_dmem_ram_913, MEM_stage_inst_dmem_ram_914, MEM_stage_inst_dmem_ram_915, MEM_stage_inst_dmem_ram_916, MEM_stage_inst_dmem_ram_917, MEM_stage_inst_dmem_ram_918, MEM_stage_inst_dmem_ram_919, MEM_stage_inst_dmem_ram_920, MEM_stage_inst_dmem_ram_921, MEM_stage_inst_dmem_ram_922, MEM_stage_inst_dmem_ram_923, MEM_stage_inst_dmem_ram_924, MEM_stage_inst_dmem_ram_925, MEM_stage_inst_dmem_ram_926, MEM_stage_inst_dmem_ram_927, MEM_stage_inst_dmem_ram_928, MEM_stage_inst_dmem_ram_929, MEM_stage_inst_dmem_ram_930, MEM_stage_inst_dmem_ram_931, MEM_stage_inst_dmem_ram_932, MEM_stage_inst_dmem_ram_933, MEM_stage_inst_dmem_ram_934, MEM_stage_inst_dmem_ram_935, MEM_stage_inst_dmem_ram_936, MEM_stage_inst_dmem_ram_937, MEM_stage_inst_dmem_ram_938, MEM_stage_inst_dmem_ram_939, MEM_stage_inst_dmem_ram_940, MEM_stage_inst_dmem_ram_941, MEM_stage_inst_dmem_ram_942, MEM_stage_inst_dmem_ram_943, MEM_stage_inst_dmem_ram_944, MEM_stage_inst_dmem_ram_945, MEM_stage_inst_dmem_ram_946, MEM_stage_inst_dmem_ram_947, MEM_stage_inst_dmem_ram_948, MEM_stage_inst_dmem_ram_949, MEM_stage_inst_dmem_ram_950, MEM_stage_inst_dmem_ram_951, MEM_stage_inst_dmem_ram_952, MEM_stage_inst_dmem_ram_953, MEM_stage_inst_dmem_ram_954, MEM_stage_inst_dmem_ram_955, MEM_stage_inst_dmem_ram_956, MEM_stage_inst_dmem_ram_957, MEM_stage_inst_dmem_ram_958, MEM_stage_inst_dmem_ram_959, MEM_stage_inst_dmem_ram_960, MEM_stage_inst_dmem_ram_961, MEM_stage_inst_dmem_ram_962, MEM_stage_inst_dmem_ram_963, MEM_stage_inst_dmem_ram_964, MEM_stage_inst_dmem_ram_965, MEM_stage_inst_dmem_ram_966, MEM_stage_inst_dmem_ram_967, MEM_stage_inst_dmem_ram_968, MEM_stage_inst_dmem_ram_969, MEM_stage_inst_dmem_ram_970, MEM_stage_inst_dmem_ram_971, MEM_stage_inst_dmem_ram_972, MEM_stage_inst_dmem_ram_973, MEM_stage_inst_dmem_ram_974, MEM_stage_inst_dmem_ram_975, MEM_stage_inst_dmem_ram_976, MEM_stage_inst_dmem_ram_977, MEM_stage_inst_dmem_ram_978, MEM_stage_inst_dmem_ram_979, MEM_stage_inst_dmem_ram_980, MEM_stage_inst_dmem_ram_981, MEM_stage_inst_dmem_ram_982, MEM_stage_inst_dmem_ram_983, MEM_stage_inst_dmem_ram_984, MEM_stage_inst_dmem_ram_985, MEM_stage_inst_dmem_ram_986, MEM_stage_inst_dmem_ram_987, MEM_stage_inst_dmem_ram_988, MEM_stage_inst_dmem_ram_989, MEM_stage_inst_dmem_ram_990, MEM_stage_inst_dmem_ram_991, MEM_stage_inst_dmem_ram_992, MEM_stage_inst_dmem_ram_993, MEM_stage_inst_dmem_ram_994, MEM_stage_inst_dmem_ram_995, MEM_stage_inst_dmem_ram_996, MEM_stage_inst_dmem_ram_997, MEM_stage_inst_dmem_ram_998, MEM_stage_inst_dmem_ram_999, MEM_stage_inst_dmem_ram_1000, MEM_stage_inst_dmem_ram_1001, MEM_stage_inst_dmem_ram_1002, MEM_stage_inst_dmem_ram_1003, MEM_stage_inst_dmem_ram_1004, MEM_stage_inst_dmem_ram_1005, MEM_stage_inst_dmem_ram_1006, MEM_stage_inst_dmem_ram_1007, MEM_stage_inst_dmem_ram_1008, MEM_stage_inst_dmem_ram_1009, MEM_stage_inst_dmem_ram_1010, MEM_stage_inst_dmem_ram_1011, MEM_stage_inst_dmem_ram_1012, MEM_stage_inst_dmem_ram_1013, MEM_stage_inst_dmem_ram_1014, MEM_stage_inst_dmem_ram_1015, MEM_stage_inst_dmem_ram_1016, MEM_stage_inst_dmem_ram_1017, MEM_stage_inst_dmem_ram_1018, MEM_stage_inst_dmem_ram_1019, MEM_stage_inst_dmem_ram_1020, MEM_stage_inst_dmem_ram_1021, MEM_stage_inst_dmem_ram_1022, MEM_stage_inst_dmem_ram_1023, MEM_stage_inst_dmem_ram_1, MEM_stage_inst_dmem_ram_2, MEM_stage_inst_dmem_ram_3, MEM_stage_inst_dmem_ram_4, MEM_stage_inst_dmem_ram_5, MEM_stage_inst_dmem_ram_6, MEM_stage_inst_dmem_ram_7, MEM_stage_inst_dmem_ram_8, MEM_stage_inst_dmem_ram_9, MEM_stage_inst_dmem_ram_10, MEM_stage_inst_dmem_ram_11, MEM_stage_inst_dmem_ram_12, MEM_stage_inst_dmem_ram_13, MEM_stage_inst_dmem_ram_14, MEM_stage_inst_dmem_ram_15, MEM_stage_inst_dmem_ram_16, MEM_stage_inst_dmem_ram_17, MEM_stage_inst_dmem_ram_18, MEM_stage_inst_dmem_ram_19, MEM_stage_inst_dmem_ram_20, MEM_stage_inst_dmem_ram_21, MEM_stage_inst_dmem_ram_22, MEM_stage_inst_dmem_ram_23, MEM_stage_inst_dmem_ram_24, MEM_stage_inst_dmem_ram_25, MEM_stage_inst_dmem_ram_26, MEM_stage_inst_dmem_ram_27, MEM_stage_inst_dmem_ram_28, MEM_stage_inst_dmem_ram_29, MEM_stage_inst_dmem_ram_30, MEM_stage_inst_dmem_ram_31, MEM_stage_inst_dmem_ram_32, MEM_stage_inst_dmem_ram_33, MEM_stage_inst_dmem_ram_34, MEM_stage_inst_dmem_ram_35, MEM_stage_inst_dmem_ram_36, MEM_stage_inst_dmem_ram_37, MEM_stage_inst_dmem_ram_38, MEM_stage_inst_dmem_ram_39, MEM_stage_inst_dmem_ram_40, MEM_stage_inst_dmem_ram_41, MEM_stage_inst_dmem_ram_42, MEM_stage_inst_dmem_ram_43, MEM_stage_inst_dmem_ram_44, MEM_stage_inst_dmem_ram_45, MEM_stage_inst_dmem_ram_46, MEM_stage_inst_dmem_ram_47, MEM_stage_inst_dmem_ram_48, MEM_stage_inst_dmem_ram_49, MEM_stage_inst_dmem_ram_50, MEM_stage_inst_dmem_ram_51, MEM_stage_inst_dmem_ram_52, MEM_stage_inst_dmem_ram_53, MEM_stage_inst_dmem_ram_54, MEM_stage_inst_dmem_ram_55, MEM_stage_inst_dmem_ram_56, MEM_stage_inst_dmem_ram_57, MEM_stage_inst_dmem_ram_58, MEM_stage_inst_dmem_ram_59, MEM_stage_inst_dmem_ram_60, MEM_stage_inst_dmem_ram_61, MEM_stage_inst_dmem_ram_62, MEM_stage_inst_dmem_ram_63, MEM_stage_inst_dmem_ram_64, MEM_stage_inst_dmem_ram_65, MEM_stage_inst_dmem_ram_66, MEM_stage_inst_dmem_ram_67, MEM_stage_inst_dmem_ram_68, MEM_stage_inst_dmem_ram_69, MEM_stage_inst_dmem_ram_70, MEM_stage_inst_dmem_ram_71, MEM_stage_inst_dmem_ram_72, MEM_stage_inst_dmem_ram_73, MEM_stage_inst_dmem_ram_74, MEM_stage_inst_dmem_ram_75, MEM_stage_inst_dmem_ram_76, MEM_stage_inst_dmem_ram_77, MEM_stage_inst_dmem_ram_78, MEM_stage_inst_dmem_ram_79, MEM_stage_inst_dmem_ram_80, MEM_stage_inst_dmem_ram_81, MEM_stage_inst_dmem_ram_82, MEM_stage_inst_dmem_ram_83, MEM_stage_inst_dmem_ram_84, MEM_stage_inst_dmem_ram_85, MEM_stage_inst_dmem_ram_86, MEM_stage_inst_dmem_ram_87, MEM_stage_inst_dmem_ram_88, MEM_stage_inst_dmem_ram_89, MEM_stage_inst_dmem_ram_90, MEM_stage_inst_dmem_ram_91, MEM_stage_inst_dmem_ram_92, MEM_stage_inst_dmem_ram_93, MEM_stage_inst_dmem_ram_94, MEM_stage_inst_dmem_ram_95, MEM_stage_inst_dmem_ram_96, MEM_stage_inst_dmem_ram_97, MEM_stage_inst_dmem_ram_98, MEM_stage_inst_dmem_ram_99, MEM_stage_inst_dmem_ram_100, MEM_stage_inst_dmem_ram_101, MEM_stage_inst_dmem_ram_102, MEM_stage_inst_dmem_ram_103, MEM_stage_inst_dmem_ram_104, MEM_stage_inst_dmem_ram_105, MEM_stage_inst_dmem_ram_106, MEM_stage_inst_dmem_ram_107, MEM_stage_inst_dmem_ram_108, MEM_stage_inst_dmem_ram_109, MEM_stage_inst_dmem_ram_110, MEM_stage_inst_dmem_ram_111, MEM_stage_inst_dmem_ram_112, MEM_stage_inst_dmem_ram_113, MEM_stage_inst_dmem_ram_114, MEM_stage_inst_dmem_ram_115, MEM_stage_inst_dmem_ram_116, MEM_stage_inst_dmem_ram_117, MEM_stage_inst_dmem_ram_118, MEM_stage_inst_dmem_ram_119, MEM_stage_inst_dmem_ram_120, MEM_stage_inst_dmem_ram_121, MEM_stage_inst_dmem_ram_122, MEM_stage_inst_dmem_ram_123, MEM_stage_inst_dmem_ram_124, MEM_stage_inst_dmem_ram_125, MEM_stage_inst_dmem_ram_126, MEM_stage_inst_dmem_ram_127, MEM_stage_inst_dmem_ram_128, MEM_stage_inst_dmem_ram_129, MEM_stage_inst_dmem_ram_130, MEM_stage_inst_dmem_ram_131, MEM_stage_inst_dmem_ram_132, MEM_stage_inst_dmem_ram_133, MEM_stage_inst_dmem_ram_134, MEM_stage_inst_dmem_ram_135, MEM_stage_inst_dmem_ram_136, MEM_stage_inst_dmem_ram_137, MEM_stage_inst_dmem_ram_138, MEM_stage_inst_dmem_ram_139, MEM_stage_inst_dmem_ram_140, MEM_stage_inst_dmem_ram_141, MEM_stage_inst_dmem_ram_142, MEM_stage_inst_dmem_ram_143, MEM_stage_inst_dmem_ram_144, MEM_stage_inst_dmem_ram_145, MEM_stage_inst_dmem_ram_146, MEM_stage_inst_dmem_ram_147, MEM_stage_inst_dmem_ram_148, MEM_stage_inst_dmem_ram_149, MEM_stage_inst_dmem_ram_150, MEM_stage_inst_dmem_ram_151, MEM_stage_inst_dmem_ram_152, MEM_stage_inst_dmem_ram_153, MEM_stage_inst_dmem_ram_154, MEM_stage_inst_dmem_ram_155, MEM_stage_inst_dmem_ram_156, MEM_stage_inst_dmem_ram_157, MEM_stage_inst_dmem_ram_158, MEM_stage_inst_dmem_ram_159, MEM_stage_inst_dmem_ram_160, MEM_stage_inst_dmem_ram_161, MEM_stage_inst_dmem_ram_162, MEM_stage_inst_dmem_ram_163, MEM_stage_inst_dmem_ram_164, MEM_stage_inst_dmem_ram_165, MEM_stage_inst_dmem_ram_166, MEM_stage_inst_dmem_ram_167, MEM_stage_inst_dmem_ram_168, MEM_stage_inst_dmem_ram_169, MEM_stage_inst_dmem_ram_170, MEM_stage_inst_dmem_ram_171, MEM_stage_inst_dmem_ram_172, MEM_stage_inst_dmem_ram_173, MEM_stage_inst_dmem_ram_174, MEM_stage_inst_dmem_ram_175, MEM_stage_inst_dmem_ram_176, MEM_stage_inst_dmem_ram_177, MEM_stage_inst_dmem_ram_178, MEM_stage_inst_dmem_ram_179, MEM_stage_inst_dmem_ram_180, MEM_stage_inst_dmem_ram_181, MEM_stage_inst_dmem_ram_182, MEM_stage_inst_dmem_ram_183, MEM_stage_inst_dmem_ram_184, MEM_stage_inst_dmem_ram_185, MEM_stage_inst_dmem_ram_186, MEM_stage_inst_dmem_ram_187, MEM_stage_inst_dmem_ram_188, MEM_stage_inst_dmem_ram_189, MEM_stage_inst_dmem_ram_190, MEM_stage_inst_dmem_ram_191, MEM_stage_inst_dmem_ram_192, MEM_stage_inst_dmem_ram_193, MEM_stage_inst_dmem_ram_194, MEM_stage_inst_dmem_ram_195, MEM_stage_inst_dmem_ram_196, MEM_stage_inst_dmem_ram_197, MEM_stage_inst_dmem_ram_198, MEM_stage_inst_dmem_ram_199, MEM_stage_inst_dmem_ram_200, MEM_stage_inst_dmem_ram_201, MEM_stage_inst_dmem_ram_202, MEM_stage_inst_dmem_ram_203, MEM_stage_inst_dmem_ram_204, MEM_stage_inst_dmem_ram_205, MEM_stage_inst_dmem_ram_206, MEM_stage_inst_dmem_ram_207, MEM_stage_inst_dmem_ram_208, MEM_stage_inst_dmem_ram_209, MEM_stage_inst_dmem_ram_210, MEM_stage_inst_dmem_ram_211, MEM_stage_inst_dmem_ram_212, MEM_stage_inst_dmem_ram_213, MEM_stage_inst_dmem_ram_214, MEM_stage_inst_dmem_ram_215, MEM_stage_inst_dmem_ram_216, MEM_stage_inst_dmem_ram_217, MEM_stage_inst_dmem_ram_218, MEM_stage_inst_dmem_ram_219, MEM_stage_inst_dmem_ram_220, MEM_stage_inst_dmem_ram_221, MEM_stage_inst_dmem_ram_222, MEM_stage_inst_dmem_ram_223, MEM_stage_inst_dmem_ram_224, MEM_stage_inst_dmem_ram_225, MEM_stage_inst_dmem_ram_226, MEM_stage_inst_dmem_ram_227, MEM_stage_inst_dmem_ram_228, MEM_stage_inst_dmem_ram_229, MEM_stage_inst_dmem_ram_230, MEM_stage_inst_dmem_ram_231, MEM_stage_inst_dmem_ram_232, MEM_stage_inst_dmem_ram_233, MEM_stage_inst_dmem_ram_234, MEM_stage_inst_dmem_ram_235, MEM_stage_inst_dmem_ram_236, MEM_stage_inst_dmem_ram_237, MEM_stage_inst_dmem_ram_238, MEM_stage_inst_dmem_ram_239, MEM_stage_inst_dmem_ram_240, MEM_stage_inst_dmem_ram_241, MEM_stage_inst_dmem_ram_242, MEM_stage_inst_dmem_ram_243, MEM_stage_inst_dmem_ram_244, MEM_stage_inst_dmem_ram_245, MEM_stage_inst_dmem_ram_246, MEM_stage_inst_dmem_ram_247, MEM_stage_inst_dmem_ram_248, MEM_stage_inst_dmem_ram_249, MEM_stage_inst_dmem_ram_250, MEM_stage_inst_dmem_ram_251, MEM_stage_inst_dmem_ram_252, MEM_stage_inst_dmem_ram_253, MEM_stage_inst_dmem_ram_254, MEM_stage_inst_dmem_ram_255, MEM_stage_inst_dmem_ram_256, MEM_stage_inst_dmem_ram_257, MEM_stage_inst_dmem_ram_258, MEM_stage_inst_dmem_ram_259, MEM_stage_inst_dmem_ram_260, MEM_stage_inst_dmem_ram_261, MEM_stage_inst_dmem_ram_262, MEM_stage_inst_dmem_ram_263, MEM_stage_inst_dmem_ram_264, MEM_stage_inst_dmem_ram_265, MEM_stage_inst_dmem_ram_266, MEM_stage_inst_dmem_ram_267, MEM_stage_inst_dmem_ram_268, MEM_stage_inst_dmem_ram_269, MEM_stage_inst_dmem_ram_270, MEM_stage_inst_dmem_ram_271, MEM_stage_inst_dmem_ram_272, MEM_stage_inst_dmem_ram_273, MEM_stage_inst_dmem_ram_274, MEM_stage_inst_dmem_ram_275, MEM_stage_inst_dmem_ram_276, MEM_stage_inst_dmem_ram_277, MEM_stage_inst_dmem_ram_278, MEM_stage_inst_dmem_ram_279, MEM_stage_inst_dmem_ram_280, MEM_stage_inst_dmem_ram_281, MEM_stage_inst_dmem_ram_282, MEM_stage_inst_dmem_ram_283, MEM_stage_inst_dmem_ram_284, MEM_stage_inst_dmem_ram_285, MEM_stage_inst_dmem_ram_286, MEM_stage_inst_dmem_ram_287, MEM_stage_inst_dmem_ram_288, MEM_stage_inst_dmem_ram_289, MEM_stage_inst_dmem_ram_290, MEM_stage_inst_dmem_ram_291, MEM_stage_inst_dmem_ram_292, MEM_stage_inst_dmem_ram_293, MEM_stage_inst_dmem_ram_294, MEM_stage_inst_dmem_ram_295, MEM_stage_inst_dmem_ram_296, MEM_stage_inst_dmem_ram_297, MEM_stage_inst_dmem_ram_298, MEM_stage_inst_dmem_ram_299, MEM_stage_inst_dmem_ram_300, MEM_stage_inst_dmem_ram_301, MEM_stage_inst_dmem_ram_302, MEM_stage_inst_dmem_ram_303, MEM_stage_inst_dmem_ram_304, MEM_stage_inst_dmem_ram_305, MEM_stage_inst_dmem_ram_306, MEM_stage_inst_dmem_ram_307, MEM_stage_inst_dmem_ram_308, MEM_stage_inst_dmem_ram_309, MEM_stage_inst_dmem_ram_310, MEM_stage_inst_dmem_ram_311, MEM_stage_inst_dmem_ram_312, MEM_stage_inst_dmem_ram_313, MEM_stage_inst_dmem_ram_314, MEM_stage_inst_dmem_ram_315, MEM_stage_inst_dmem_ram_316, MEM_stage_inst_dmem_ram_317, MEM_stage_inst_dmem_ram_318, MEM_stage_inst_dmem_ram_319, MEM_stage_inst_dmem_ram_320, MEM_stage_inst_dmem_ram_321, MEM_stage_inst_dmem_ram_322, MEM_stage_inst_dmem_ram_323, MEM_stage_inst_dmem_ram_324, MEM_stage_inst_dmem_ram_325, MEM_stage_inst_dmem_ram_326, MEM_stage_inst_dmem_ram_327, MEM_stage_inst_dmem_ram_328, MEM_stage_inst_dmem_ram_329, MEM_stage_inst_dmem_ram_330, MEM_stage_inst_dmem_ram_331, MEM_stage_inst_dmem_ram_332, MEM_stage_inst_dmem_ram_333, MEM_stage_inst_dmem_ram_334, MEM_stage_inst_dmem_ram_335, MEM_stage_inst_dmem_ram_336, MEM_stage_inst_dmem_ram_337, MEM_stage_inst_dmem_ram_338, MEM_stage_inst_dmem_ram_339, MEM_stage_inst_dmem_ram_340, MEM_stage_inst_dmem_ram_341, MEM_stage_inst_dmem_ram_342, MEM_stage_inst_dmem_ram_343, MEM_stage_inst_dmem_ram_344, MEM_stage_inst_dmem_ram_345, MEM_stage_inst_dmem_ram_346, MEM_stage_inst_dmem_ram_347, MEM_stage_inst_dmem_ram_348, MEM_stage_inst_dmem_ram_349, MEM_stage_inst_dmem_ram_350, MEM_stage_inst_dmem_ram_351, MEM_stage_inst_dmem_ram_352, MEM_stage_inst_dmem_ram_353, MEM_stage_inst_dmem_ram_354, MEM_stage_inst_dmem_ram_355, MEM_stage_inst_dmem_ram_356, MEM_stage_inst_dmem_ram_357, MEM_stage_inst_dmem_ram_358, MEM_stage_inst_dmem_ram_359, MEM_stage_inst_dmem_ram_360, MEM_stage_inst_dmem_ram_361, MEM_stage_inst_dmem_ram_362, MEM_stage_inst_dmem_ram_363, MEM_stage_inst_dmem_ram_364, MEM_stage_inst_dmem_ram_365, MEM_stage_inst_dmem_ram_366, MEM_stage_inst_dmem_ram_367, MEM_stage_inst_dmem_ram_368, MEM_stage_inst_dmem_ram_369, MEM_stage_inst_dmem_ram_370, MEM_stage_inst_dmem_ram_371, MEM_stage_inst_dmem_ram_372, MEM_stage_inst_dmem_ram_373, MEM_stage_inst_dmem_ram_374, MEM_stage_inst_dmem_ram_375, MEM_stage_inst_dmem_ram_376, MEM_stage_inst_dmem_ram_377, MEM_stage_inst_dmem_ram_378, MEM_stage_inst_dmem_ram_379, MEM_stage_inst_dmem_ram_380, MEM_stage_inst_dmem_ram_381, MEM_stage_inst_dmem_ram_382, MEM_stage_inst_dmem_ram_383, MEM_stage_inst_dmem_ram_384, MEM_stage_inst_dmem_ram_385, MEM_stage_inst_dmem_ram_386, MEM_stage_inst_dmem_ram_387, MEM_stage_inst_dmem_ram_388, MEM_stage_inst_dmem_ram_389, MEM_stage_inst_dmem_ram_390, MEM_stage_inst_dmem_ram_391, MEM_stage_inst_dmem_ram_392, MEM_stage_inst_dmem_ram_393, MEM_stage_inst_dmem_ram_394, MEM_stage_inst_dmem_ram_395, MEM_stage_inst_dmem_ram_396, MEM_stage_inst_dmem_ram_397, MEM_stage_inst_dmem_ram_398, MEM_stage_inst_dmem_ram_399, MEM_stage_inst_dmem_ram_400, MEM_stage_inst_dmem_ram_401, MEM_stage_inst_dmem_ram_402, MEM_stage_inst_dmem_ram_403, MEM_stage_inst_dmem_ram_404, MEM_stage_inst_dmem_ram_405, MEM_stage_inst_dmem_ram_406, MEM_stage_inst_dmem_ram_407, MEM_stage_inst_dmem_ram_408, MEM_stage_inst_dmem_ram_409, MEM_stage_inst_dmem_ram_410, MEM_stage_inst_dmem_ram_411, MEM_stage_inst_dmem_ram_412, MEM_stage_inst_dmem_ram_413, MEM_stage_inst_dmem_ram_414, MEM_stage_inst_dmem_ram_415, MEM_stage_inst_dmem_ram_416, MEM_stage_inst_dmem_ram_417, MEM_stage_inst_dmem_ram_418, MEM_stage_inst_dmem_ram_419, MEM_stage_inst_dmem_ram_420, MEM_stage_inst_dmem_ram_421, MEM_stage_inst_dmem_ram_422, MEM_stage_inst_dmem_ram_423, MEM_stage_inst_dmem_ram_424, MEM_stage_inst_dmem_ram_425, MEM_stage_inst_dmem_ram_426, MEM_stage_inst_dmem_ram_427, MEM_stage_inst_dmem_ram_428, MEM_stage_inst_dmem_ram_429, MEM_stage_inst_dmem_ram_430, MEM_stage_inst_dmem_ram_431, MEM_stage_inst_dmem_ram_432, MEM_stage_inst_dmem_ram_433, MEM_stage_inst_dmem_ram_434, MEM_stage_inst_dmem_ram_435, MEM_stage_inst_dmem_ram_436, MEM_stage_inst_dmem_ram_437, MEM_stage_inst_dmem_ram_438, MEM_stage_inst_dmem_ram_439, MEM_stage_inst_dmem_ram_440, MEM_stage_inst_dmem_ram_441, MEM_stage_inst_dmem_ram_442, MEM_stage_inst_dmem_ram_443, MEM_stage_inst_dmem_ram_444, MEM_stage_inst_dmem_ram_445, MEM_stage_inst_dmem_ram_446, MEM_stage_inst_dmem_ram_447, MEM_stage_inst_dmem_ram_448, MEM_stage_inst_dmem_ram_449, MEM_stage_inst_dmem_ram_450, MEM_stage_inst_dmem_ram_451, MEM_stage_inst_dmem_ram_452, MEM_stage_inst_dmem_ram_453, MEM_stage_inst_dmem_ram_454, MEM_stage_inst_dmem_ram_455, MEM_stage_inst_dmem_ram_456, MEM_stage_inst_dmem_ram_457, MEM_stage_inst_dmem_ram_458, MEM_stage_inst_dmem_ram_459, MEM_stage_inst_dmem_ram_460, MEM_stage_inst_dmem_ram_461, MEM_stage_inst_dmem_ram_462, MEM_stage_inst_dmem_ram_463, MEM_stage_inst_dmem_ram_464, MEM_stage_inst_dmem_ram_465, MEM_stage_inst_dmem_ram_466, MEM_stage_inst_dmem_ram_467, MEM_stage_inst_dmem_ram_468, MEM_stage_inst_dmem_ram_469, MEM_stage_inst_dmem_ram_470, MEM_stage_inst_dmem_ram_471, MEM_stage_inst_dmem_ram_472, MEM_stage_inst_dmem_ram_473, MEM_stage_inst_dmem_ram_474, MEM_stage_inst_dmem_ram_475, MEM_stage_inst_dmem_ram_476, MEM_stage_inst_dmem_ram_477, MEM_stage_inst_dmem_ram_478, MEM_stage_inst_dmem_ram_479, MEM_stage_inst_dmem_ram_480, MEM_stage_inst_dmem_ram_481, MEM_stage_inst_dmem_ram_482, MEM_stage_inst_dmem_ram_483, MEM_stage_inst_dmem_ram_484, MEM_stage_inst_dmem_ram_485, MEM_stage_inst_dmem_ram_486, MEM_stage_inst_dmem_ram_487, MEM_stage_inst_dmem_ram_488, MEM_stage_inst_dmem_ram_489, MEM_stage_inst_dmem_ram_490, MEM_stage_inst_dmem_ram_491, MEM_stage_inst_dmem_ram_492, MEM_stage_inst_dmem_ram_493, MEM_stage_inst_dmem_ram_494, MEM_stage_inst_dmem_ram_495, MEM_stage_inst_dmem_ram_496, MEM_stage_inst_dmem_ram_497, MEM_stage_inst_dmem_ram_498, MEM_stage_inst_dmem_ram_499, MEM_stage_inst_dmem_ram_500, MEM_stage_inst_dmem_ram_501, MEM_stage_inst_dmem_ram_502, MEM_stage_inst_dmem_ram_503, MEM_stage_inst_dmem_ram_504, MEM_stage_inst_dmem_ram_505, MEM_stage_inst_dmem_ram_506, MEM_stage_inst_dmem_ram_507, MEM_stage_inst_dmem_ram_508, MEM_stage_inst_dmem_ram_509, MEM_stage_inst_dmem_ram_510, MEM_stage_inst_dmem_ram_511, MEM_stage_inst_dmem_ram_0 );
input clk, rst, reg_write_dest_2, n3475, mem_op_dest_0, reg_write_dest_0, mem_op_dest_1, reg_write_dest_1, n3484, mem_op_dest_2, EX_pipeline_reg_out_0, EX_pipeline_reg_out_4, n3522, reg_write_en, n3516, EX_pipeline_reg_out_37, MEM_pipeline_reg_out_36, EX_pipeline_reg_out_20, EX_pipeline_reg_out_22, MEM_pipeline_reg_out_21, EX_pipeline_reg_out_5, EX_pipeline_reg_out_30, MEM_pipeline_reg_out_29, EX_pipeline_reg_out_13, EX_pipeline_reg_out_32, MEM_pipeline_reg_out_31, EX_pipeline_reg_out_15, EX_pipeline_reg_out_34, MEM_pipeline_reg_out_33, EX_pipeline_reg_out_17, EX_pipeline_reg_out_36, MEM_pipeline_reg_out_35, EX_pipeline_reg_out_19, EX_pipeline_reg_out_26, MEM_pipeline_reg_out_25, EX_pipeline_reg_out_9, EX_pipeline_reg_out_28, MEM_pipeline_reg_out_27, EX_pipeline_reg_out_11, EX_pipeline_reg_out_33, MEM_pipeline_reg_out_32, EX_pipeline_reg_out_16, EX_pipeline_reg_out_35, MEM_pipeline_reg_out_34, EX_pipeline_reg_out_18, EX_pipeline_reg_out_24, MEM_pipeline_reg_out_23, EX_pipeline_reg_out_7, EX_pipeline_reg_out_25, MEM_pipeline_reg_out_24, EX_pipeline_reg_out_8, EX_pipeline_reg_out_23, MEM_pipeline_reg_out_22, EX_pipeline_reg_out_6, EX_pipeline_reg_out_27, MEM_pipeline_reg_out_26, EX_pipeline_reg_out_10, EX_pipeline_reg_out_31, MEM_pipeline_reg_out_30, EX_pipeline_reg_out_14, EX_pipeline_reg_out_29, MEM_pipeline_reg_out_28, EX_pipeline_reg_out_12, MEM_pipeline_reg_out_5, MEM_pipeline_reg_out_6, MEM_pipeline_reg_out_7, MEM_pipeline_reg_out_8, MEM_pipeline_reg_out_9, MEM_pipeline_reg_out_10, MEM_pipeline_reg_out_11, MEM_pipeline_reg_out_12, MEM_pipeline_reg_out_13, MEM_pipeline_reg_out_14, MEM_pipeline_reg_out_15, MEM_pipeline_reg_out_16, MEM_pipeline_reg_out_17, MEM_pipeline_reg_out_18, MEM_pipeline_reg_out_19, MEM_pipeline_reg_out_20, n3511, branch_offset_imm_3, n3513, branch_offset_imm_5, n3509, branch_offset_imm_1, n3514, branch_offset_imm_4, n3512, ID_stage_inst_instruction_reg_14, n3510, ID_stage_inst_instruction_reg_13, branch_offset_imm_0, reg_read_addr_1_0, reg_read_addr_1_1, n3480, reg_read_addr_1_2, n3479, ID_stage_inst_instruction_reg_9, ex_op_dest_0, ID_stage_inst_instruction_reg_10, n3515, ex_op_dest_1, ID_stage_inst_instruction_reg_11, ex_op_dest_2, ID_stage_inst_instruction_reg_12, n3487, ID_stage_inst_instruction_reg_15, ID_pipeline_reg_out_55, ID_pipeline_reg_out_54, n3473, ID_pipeline_reg_out_56, n3488, ID_pipeline_reg_out_0, ID_pipeline_reg_out_4, ID_pipeline_reg_out_21, register_file_inst_reg_array_111, ID_pipeline_reg_out_53, n3485, register_file_inst_reg_array_95, register_file_inst_reg_array_79, register_file_inst_reg_array_63, n3492, register_file_inst_reg_array_47, register_file_inst_reg_array_31, register_file_inst_reg_array_15, ID_pipeline_reg_out_20, ID_pipeline_reg_out_37, register_file_inst_reg_array_96, register_file_inst_reg_array_80, register_file_inst_reg_array_64, register_file_inst_reg_array_48, n3491, register_file_inst_reg_array_32, register_file_inst_reg_array_16, register_file_inst_reg_array_0, ID_pipeline_reg_out_5, ID_pipeline_reg_out_38, n3486, register_file_inst_reg_array_104, register_file_inst_reg_array_88, register_file_inst_reg_array_72, register_file_inst_reg_array_56, n3500, register_file_inst_reg_array_40, register_file_inst_reg_array_24, register_file_inst_reg_array_8, ID_pipeline_reg_out_13, ID_pipeline_reg_out_30, ID_pipeline_reg_out_46, register_file_inst_reg_array_106, register_file_inst_reg_array_90, register_file_inst_reg_array_74, register_file_inst_reg_array_58, n3504, register_file_inst_reg_array_42, register_file_inst_reg_array_26, register_file_inst_reg_array_10, ID_pipeline_reg_out_15, ID_pipeline_reg_out_32, ID_pipeline_reg_out_48, register_file_inst_reg_array_108, register_file_inst_reg_array_92, register_file_inst_reg_array_76, register_file_inst_reg_array_60, n3495, register_file_inst_reg_array_44, register_file_inst_reg_array_28, register_file_inst_reg_array_12, ID_pipeline_reg_out_17, ID_pipeline_reg_out_34, ID_pipeline_reg_out_50, register_file_inst_reg_array_110, register_file_inst_reg_array_94, register_file_inst_reg_array_78, register_file_inst_reg_array_62, n3501, register_file_inst_reg_array_46, register_file_inst_reg_array_30, register_file_inst_reg_array_14, ID_pipeline_reg_out_19, ID_pipeline_reg_out_36, ID_pipeline_reg_out_52, register_file_inst_reg_array_100, register_file_inst_reg_array_84, register_file_inst_reg_array_68, register_file_inst_reg_array_52, n3496, register_file_inst_reg_array_36, register_file_inst_reg_array_20, register_file_inst_reg_array_4, ID_pipeline_reg_out_9, ID_pipeline_reg_out_26, n3474, ID_pipeline_reg_out_42, register_file_inst_reg_array_102, register_file_inst_reg_array_86, register_file_inst_reg_array_70, register_file_inst_reg_array_54, n3503, register_file_inst_reg_array_38, register_file_inst_reg_array_22, register_file_inst_reg_array_6, ID_pipeline_reg_out_11, ID_pipeline_reg_out_28, ID_pipeline_reg_out_44, register_file_inst_reg_array_107, register_file_inst_reg_array_91, register_file_inst_reg_array_75, register_file_inst_reg_array_59, n3498, register_file_inst_reg_array_43, register_file_inst_reg_array_27, register_file_inst_reg_array_11, ID_pipeline_reg_out_16, ID_pipeline_reg_out_33, ID_pipeline_reg_out_49, register_file_inst_reg_array_109, register_file_inst_reg_array_93, register_file_inst_reg_array_77, register_file_inst_reg_array_61, n3502, register_file_inst_reg_array_45, register_file_inst_reg_array_29, register_file_inst_reg_array_13, ID_pipeline_reg_out_18, ID_pipeline_reg_out_35, ID_pipeline_reg_out_51, n3483, register_file_inst_reg_array_98, register_file_inst_reg_array_82, register_file_inst_reg_array_66, register_file_inst_reg_array_50, n3494, register_file_inst_reg_array_34, register_file_inst_reg_array_18, register_file_inst_reg_array_2, ID_pipeline_reg_out_7, ID_pipeline_reg_out_40, n3508, register_file_inst_reg_array_99, register_file_inst_reg_array_83, register_file_inst_reg_array_67, register_file_inst_reg_array_51, n3506, register_file_inst_reg_array_35, register_file_inst_reg_array_19, register_file_inst_reg_array_3, ID_pipeline_reg_out_8, ID_pipeline_reg_out_41, n3482, register_file_inst_reg_array_97, register_file_inst_reg_array_81, register_file_inst_reg_array_65, register_file_inst_reg_array_49, n3499, register_file_inst_reg_array_33, register_file_inst_reg_array_17, register_file_inst_reg_array_1, ID_pipeline_reg_out_6, ID_pipeline_reg_out_39, register_file_inst_reg_array_101, register_file_inst_reg_array_85, register_file_inst_reg_array_69, register_file_inst_reg_array_53, n3497, register_file_inst_reg_array_37, register_file_inst_reg_array_21, register_file_inst_reg_array_5, ID_pipeline_reg_out_10, ID_pipeline_reg_out_27, ID_pipeline_reg_out_43, n3489, register_file_inst_reg_array_105, register_file_inst_reg_array_89, register_file_inst_reg_array_73, register_file_inst_reg_array_57, n3493, register_file_inst_reg_array_41, register_file_inst_reg_array_25, register_file_inst_reg_array_9, ID_pipeline_reg_out_14, ID_pipeline_reg_out_31, ID_pipeline_reg_out_47, n3490, register_file_inst_reg_array_103, register_file_inst_reg_array_87, register_file_inst_reg_array_71, register_file_inst_reg_array_55, n3505, register_file_inst_reg_array_39, register_file_inst_reg_array_23, register_file_inst_reg_array_7, ID_pipeline_reg_out_12, ID_pipeline_reg_out_29, ID_pipeline_reg_out_45, n3507, n3481, ID_pipeline_reg_out_23, n3478, MEM_pipeline_reg_out_0, n3477, ID_pipeline_reg_out_24, n3476, ID_pipeline_reg_out_22, n3472, ID_pipeline_reg_out_25, n3471, MEM_stage_inst_dmem_ram_3584, MEM_stage_inst_dmem_ram_3585, MEM_stage_inst_dmem_ram_3586, MEM_stage_inst_dmem_ram_3587, MEM_stage_inst_dmem_ram_3588, MEM_stage_inst_dmem_ram_3589, MEM_stage_inst_dmem_ram_3590, MEM_stage_inst_dmem_ram_3591, MEM_stage_inst_dmem_ram_3592, MEM_stage_inst_dmem_ram_3593, MEM_stage_inst_dmem_ram_3594, MEM_stage_inst_dmem_ram_3595, MEM_stage_inst_dmem_ram_3596, MEM_stage_inst_dmem_ram_3597, MEM_stage_inst_dmem_ram_3598, MEM_stage_inst_dmem_ram_3599, MEM_stage_inst_dmem_ram_3600, MEM_stage_inst_dmem_ram_3601, MEM_stage_inst_dmem_ram_3602, MEM_stage_inst_dmem_ram_3603, MEM_stage_inst_dmem_ram_3604, MEM_stage_inst_dmem_ram_3605, MEM_stage_inst_dmem_ram_3606, MEM_stage_inst_dmem_ram_3607, MEM_stage_inst_dmem_ram_3608, MEM_stage_inst_dmem_ram_3609, MEM_stage_inst_dmem_ram_3610, MEM_stage_inst_dmem_ram_3611, MEM_stage_inst_dmem_ram_3612, MEM_stage_inst_dmem_ram_3613, MEM_stage_inst_dmem_ram_3614, MEM_stage_inst_dmem_ram_3615, MEM_stage_inst_dmem_ram_3616, MEM_stage_inst_dmem_ram_3617, MEM_stage_inst_dmem_ram_3618, MEM_stage_inst_dmem_ram_3619, MEM_stage_inst_dmem_ram_3620, MEM_stage_inst_dmem_ram_3621, MEM_stage_inst_dmem_ram_3622, MEM_stage_inst_dmem_ram_3623, MEM_stage_inst_dmem_ram_3624, MEM_stage_inst_dmem_ram_3625, MEM_stage_inst_dmem_ram_3626, MEM_stage_inst_dmem_ram_3627, MEM_stage_inst_dmem_ram_3628, MEM_stage_inst_dmem_ram_3629, MEM_stage_inst_dmem_ram_3630, MEM_stage_inst_dmem_ram_3631, MEM_stage_inst_dmem_ram_3632, MEM_stage_inst_dmem_ram_3633, MEM_stage_inst_dmem_ram_3634, MEM_stage_inst_dmem_ram_3635, MEM_stage_inst_dmem_ram_3636, MEM_stage_inst_dmem_ram_3637, MEM_stage_inst_dmem_ram_3638, MEM_stage_inst_dmem_ram_3639, MEM_stage_inst_dmem_ram_3640, MEM_stage_inst_dmem_ram_3641, MEM_stage_inst_dmem_ram_3642, MEM_stage_inst_dmem_ram_3643, MEM_stage_inst_dmem_ram_3644, MEM_stage_inst_dmem_ram_3645, MEM_stage_inst_dmem_ram_3646, MEM_stage_inst_dmem_ram_3647, MEM_stage_inst_dmem_ram_3648, MEM_stage_inst_dmem_ram_3649, MEM_stage_inst_dmem_ram_3650, MEM_stage_inst_dmem_ram_3651, MEM_stage_inst_dmem_ram_3652, MEM_stage_inst_dmem_ram_3653, MEM_stage_inst_dmem_ram_3654, MEM_stage_inst_dmem_ram_3655, MEM_stage_inst_dmem_ram_3656, MEM_stage_inst_dmem_ram_3657, MEM_stage_inst_dmem_ram_3658, MEM_stage_inst_dmem_ram_3659, MEM_stage_inst_dmem_ram_3660, MEM_stage_inst_dmem_ram_3661, MEM_stage_inst_dmem_ram_3662, MEM_stage_inst_dmem_ram_3663, MEM_stage_inst_dmem_ram_3664, MEM_stage_inst_dmem_ram_3665, MEM_stage_inst_dmem_ram_3666, MEM_stage_inst_dmem_ram_3667, MEM_stage_inst_dmem_ram_3668, MEM_stage_inst_dmem_ram_3669, MEM_stage_inst_dmem_ram_3670, MEM_stage_inst_dmem_ram_3671, MEM_stage_inst_dmem_ram_3672, MEM_stage_inst_dmem_ram_3673, MEM_stage_inst_dmem_ram_3674, MEM_stage_inst_dmem_ram_3675, MEM_stage_inst_dmem_ram_3676, MEM_stage_inst_dmem_ram_3677, MEM_stage_inst_dmem_ram_3678, MEM_stage_inst_dmem_ram_3679, MEM_stage_inst_dmem_ram_3680, MEM_stage_inst_dmem_ram_3681, MEM_stage_inst_dmem_ram_3682, MEM_stage_inst_dmem_ram_3683, MEM_stage_inst_dmem_ram_3684, MEM_stage_inst_dmem_ram_3685, MEM_stage_inst_dmem_ram_3686, MEM_stage_inst_dmem_ram_3687, MEM_stage_inst_dmem_ram_3688, MEM_stage_inst_dmem_ram_3689, MEM_stage_inst_dmem_ram_3690, MEM_stage_inst_dmem_ram_3691, MEM_stage_inst_dmem_ram_3692, MEM_stage_inst_dmem_ram_3693, MEM_stage_inst_dmem_ram_3694, MEM_stage_inst_dmem_ram_3695, MEM_stage_inst_dmem_ram_3696, MEM_stage_inst_dmem_ram_3697, MEM_stage_inst_dmem_ram_3698, MEM_stage_inst_dmem_ram_3699, MEM_stage_inst_dmem_ram_3700, MEM_stage_inst_dmem_ram_3701, MEM_stage_inst_dmem_ram_3702, MEM_stage_inst_dmem_ram_3703, MEM_stage_inst_dmem_ram_3704, MEM_stage_inst_dmem_ram_3705, MEM_stage_inst_dmem_ram_3706, MEM_stage_inst_dmem_ram_3707, MEM_stage_inst_dmem_ram_3708, MEM_stage_inst_dmem_ram_3709, MEM_stage_inst_dmem_ram_3710, MEM_stage_inst_dmem_ram_3711, MEM_stage_inst_dmem_ram_3712, MEM_stage_inst_dmem_ram_3713, MEM_stage_inst_dmem_ram_3714, MEM_stage_inst_dmem_ram_3715, MEM_stage_inst_dmem_ram_3716, MEM_stage_inst_dmem_ram_3717, MEM_stage_inst_dmem_ram_3718, MEM_stage_inst_dmem_ram_3719, MEM_stage_inst_dmem_ram_3720, MEM_stage_inst_dmem_ram_3721, MEM_stage_inst_dmem_ram_3722, MEM_stage_inst_dmem_ram_3723, MEM_stage_inst_dmem_ram_3724, MEM_stage_inst_dmem_ram_3725, MEM_stage_inst_dmem_ram_3726, MEM_stage_inst_dmem_ram_3727, MEM_stage_inst_dmem_ram_3728, MEM_stage_inst_dmem_ram_3729, MEM_stage_inst_dmem_ram_3730, MEM_stage_inst_dmem_ram_3731, MEM_stage_inst_dmem_ram_3732, MEM_stage_inst_dmem_ram_3733, MEM_stage_inst_dmem_ram_3734, MEM_stage_inst_dmem_ram_3735, MEM_stage_inst_dmem_ram_3736, MEM_stage_inst_dmem_ram_3737, MEM_stage_inst_dmem_ram_3738, MEM_stage_inst_dmem_ram_3739, MEM_stage_inst_dmem_ram_3740, MEM_stage_inst_dmem_ram_3741, MEM_stage_inst_dmem_ram_3742, MEM_stage_inst_dmem_ram_3743, MEM_stage_inst_dmem_ram_3744, MEM_stage_inst_dmem_ram_3745, MEM_stage_inst_dmem_ram_3746, MEM_stage_inst_dmem_ram_3747, MEM_stage_inst_dmem_ram_3748, MEM_stage_inst_dmem_ram_3749, MEM_stage_inst_dmem_ram_3750, MEM_stage_inst_dmem_ram_3751, MEM_stage_inst_dmem_ram_3752, MEM_stage_inst_dmem_ram_3753, MEM_stage_inst_dmem_ram_3754, MEM_stage_inst_dmem_ram_3755, MEM_stage_inst_dmem_ram_3756, MEM_stage_inst_dmem_ram_3757, MEM_stage_inst_dmem_ram_3758, MEM_stage_inst_dmem_ram_3759, MEM_stage_inst_dmem_ram_3760, MEM_stage_inst_dmem_ram_3761, MEM_stage_inst_dmem_ram_3762, MEM_stage_inst_dmem_ram_3763, MEM_stage_inst_dmem_ram_3764, MEM_stage_inst_dmem_ram_3765, MEM_stage_inst_dmem_ram_3766, MEM_stage_inst_dmem_ram_3767, MEM_stage_inst_dmem_ram_3768, MEM_stage_inst_dmem_ram_3769, MEM_stage_inst_dmem_ram_3770, MEM_stage_inst_dmem_ram_3771, MEM_stage_inst_dmem_ram_3772, MEM_stage_inst_dmem_ram_3773, MEM_stage_inst_dmem_ram_3774, MEM_stage_inst_dmem_ram_3775, MEM_stage_inst_dmem_ram_3776, MEM_stage_inst_dmem_ram_3777, MEM_stage_inst_dmem_ram_3778, MEM_stage_inst_dmem_ram_3779, MEM_stage_inst_dmem_ram_3780, MEM_stage_inst_dmem_ram_3781, MEM_stage_inst_dmem_ram_3782, MEM_stage_inst_dmem_ram_3783, MEM_stage_inst_dmem_ram_3784, MEM_stage_inst_dmem_ram_3785, MEM_stage_inst_dmem_ram_3786, MEM_stage_inst_dmem_ram_3787, MEM_stage_inst_dmem_ram_3788, MEM_stage_inst_dmem_ram_3789, MEM_stage_inst_dmem_ram_3790, MEM_stage_inst_dmem_ram_3791, MEM_stage_inst_dmem_ram_3792, MEM_stage_inst_dmem_ram_3793, MEM_stage_inst_dmem_ram_3794, MEM_stage_inst_dmem_ram_3795, MEM_stage_inst_dmem_ram_3796, MEM_stage_inst_dmem_ram_3797, MEM_stage_inst_dmem_ram_3798, MEM_stage_inst_dmem_ram_3799, MEM_stage_inst_dmem_ram_3800, MEM_stage_inst_dmem_ram_3801, MEM_stage_inst_dmem_ram_3802, MEM_stage_inst_dmem_ram_3803, MEM_stage_inst_dmem_ram_3804, MEM_stage_inst_dmem_ram_3805, MEM_stage_inst_dmem_ram_3806, MEM_stage_inst_dmem_ram_3807, MEM_stage_inst_dmem_ram_3808, MEM_stage_inst_dmem_ram_3809, MEM_stage_inst_dmem_ram_3810, MEM_stage_inst_dmem_ram_3811, MEM_stage_inst_dmem_ram_3812, MEM_stage_inst_dmem_ram_3813, MEM_stage_inst_dmem_ram_3814, MEM_stage_inst_dmem_ram_3815, MEM_stage_inst_dmem_ram_3816, MEM_stage_inst_dmem_ram_3817, MEM_stage_inst_dmem_ram_3818, MEM_stage_inst_dmem_ram_3819, MEM_stage_inst_dmem_ram_3820, MEM_stage_inst_dmem_ram_3821, MEM_stage_inst_dmem_ram_3822, MEM_stage_inst_dmem_ram_3823, MEM_stage_inst_dmem_ram_3824, MEM_stage_inst_dmem_ram_3825, MEM_stage_inst_dmem_ram_3826, MEM_stage_inst_dmem_ram_3827, MEM_stage_inst_dmem_ram_3828, MEM_stage_inst_dmem_ram_3829, MEM_stage_inst_dmem_ram_3830, MEM_stage_inst_dmem_ram_3831, MEM_stage_inst_dmem_ram_3832, MEM_stage_inst_dmem_ram_3833, MEM_stage_inst_dmem_ram_3834, MEM_stage_inst_dmem_ram_3835, MEM_stage_inst_dmem_ram_3836, MEM_stage_inst_dmem_ram_3837, MEM_stage_inst_dmem_ram_3838, MEM_stage_inst_dmem_ram_3839, MEM_stage_inst_dmem_ram_3840, MEM_stage_inst_dmem_ram_3841, MEM_stage_inst_dmem_ram_3842, MEM_stage_inst_dmem_ram_3843, MEM_stage_inst_dmem_ram_3844, MEM_stage_inst_dmem_ram_3845, MEM_stage_inst_dmem_ram_3846, MEM_stage_inst_dmem_ram_3847, MEM_stage_inst_dmem_ram_3848, MEM_stage_inst_dmem_ram_3849, MEM_stage_inst_dmem_ram_3850, MEM_stage_inst_dmem_ram_3851, MEM_stage_inst_dmem_ram_3852, MEM_stage_inst_dmem_ram_3853, MEM_stage_inst_dmem_ram_3854, MEM_stage_inst_dmem_ram_3855, MEM_stage_inst_dmem_ram_3856, MEM_stage_inst_dmem_ram_3857, MEM_stage_inst_dmem_ram_3858, MEM_stage_inst_dmem_ram_3859, MEM_stage_inst_dmem_ram_3860, MEM_stage_inst_dmem_ram_3861, MEM_stage_inst_dmem_ram_3862, MEM_stage_inst_dmem_ram_3863, MEM_stage_inst_dmem_ram_3864, MEM_stage_inst_dmem_ram_3865, MEM_stage_inst_dmem_ram_3866, MEM_stage_inst_dmem_ram_3867, MEM_stage_inst_dmem_ram_3868, MEM_stage_inst_dmem_ram_3869, MEM_stage_inst_dmem_ram_3870, MEM_stage_inst_dmem_ram_3871, MEM_stage_inst_dmem_ram_3872, MEM_stage_inst_dmem_ram_3873, MEM_stage_inst_dmem_ram_3874, MEM_stage_inst_dmem_ram_3875, MEM_stage_inst_dmem_ram_3876, MEM_stage_inst_dmem_ram_3877, MEM_stage_inst_dmem_ram_3878, MEM_stage_inst_dmem_ram_3879, MEM_stage_inst_dmem_ram_3880, MEM_stage_inst_dmem_ram_3881, MEM_stage_inst_dmem_ram_3882, MEM_stage_inst_dmem_ram_3883, MEM_stage_inst_dmem_ram_3884, MEM_stage_inst_dmem_ram_3885, MEM_stage_inst_dmem_ram_3886, MEM_stage_inst_dmem_ram_3887, MEM_stage_inst_dmem_ram_3888, MEM_stage_inst_dmem_ram_3889, MEM_stage_inst_dmem_ram_3890, MEM_stage_inst_dmem_ram_3891, MEM_stage_inst_dmem_ram_3892, MEM_stage_inst_dmem_ram_3893, MEM_stage_inst_dmem_ram_3894, MEM_stage_inst_dmem_ram_3895, MEM_stage_inst_dmem_ram_3896, MEM_stage_inst_dmem_ram_3897, MEM_stage_inst_dmem_ram_3898, MEM_stage_inst_dmem_ram_3899, MEM_stage_inst_dmem_ram_3900, MEM_stage_inst_dmem_ram_3901, MEM_stage_inst_dmem_ram_3902, MEM_stage_inst_dmem_ram_3903, MEM_stage_inst_dmem_ram_3904, MEM_stage_inst_dmem_ram_3905, MEM_stage_inst_dmem_ram_3906, MEM_stage_inst_dmem_ram_3907, MEM_stage_inst_dmem_ram_3908, MEM_stage_inst_dmem_ram_3909, MEM_stage_inst_dmem_ram_3910, MEM_stage_inst_dmem_ram_3911, MEM_stage_inst_dmem_ram_3912, MEM_stage_inst_dmem_ram_3913, MEM_stage_inst_dmem_ram_3914, MEM_stage_inst_dmem_ram_3915, MEM_stage_inst_dmem_ram_3916, MEM_stage_inst_dmem_ram_3917, MEM_stage_inst_dmem_ram_3918, MEM_stage_inst_dmem_ram_3919, MEM_stage_inst_dmem_ram_3920, MEM_stage_inst_dmem_ram_3921, MEM_stage_inst_dmem_ram_3922, MEM_stage_inst_dmem_ram_3923, MEM_stage_inst_dmem_ram_3924, MEM_stage_inst_dmem_ram_3925, MEM_stage_inst_dmem_ram_3926, MEM_stage_inst_dmem_ram_3927, MEM_stage_inst_dmem_ram_3928, MEM_stage_inst_dmem_ram_3929, MEM_stage_inst_dmem_ram_3930, MEM_stage_inst_dmem_ram_3931, MEM_stage_inst_dmem_ram_3932, MEM_stage_inst_dmem_ram_3933, MEM_stage_inst_dmem_ram_3934, MEM_stage_inst_dmem_ram_3935, MEM_stage_inst_dmem_ram_3936, MEM_stage_inst_dmem_ram_3937, MEM_stage_inst_dmem_ram_3938, MEM_stage_inst_dmem_ram_3939, MEM_stage_inst_dmem_ram_3940, MEM_stage_inst_dmem_ram_3941, MEM_stage_inst_dmem_ram_3942, MEM_stage_inst_dmem_ram_3943, MEM_stage_inst_dmem_ram_3944, MEM_stage_inst_dmem_ram_3945, MEM_stage_inst_dmem_ram_3946, MEM_stage_inst_dmem_ram_3947, MEM_stage_inst_dmem_ram_3948, MEM_stage_inst_dmem_ram_3949, MEM_stage_inst_dmem_ram_3950, MEM_stage_inst_dmem_ram_3951, MEM_stage_inst_dmem_ram_3952, MEM_stage_inst_dmem_ram_3953, MEM_stage_inst_dmem_ram_3954, MEM_stage_inst_dmem_ram_3955, MEM_stage_inst_dmem_ram_3956, MEM_stage_inst_dmem_ram_3957, MEM_stage_inst_dmem_ram_3958, MEM_stage_inst_dmem_ram_3959, MEM_stage_inst_dmem_ram_3960, MEM_stage_inst_dmem_ram_3961, MEM_stage_inst_dmem_ram_3962, MEM_stage_inst_dmem_ram_3963, MEM_stage_inst_dmem_ram_3964, MEM_stage_inst_dmem_ram_3965, MEM_stage_inst_dmem_ram_3966, MEM_stage_inst_dmem_ram_3967, MEM_stage_inst_dmem_ram_3968, MEM_stage_inst_dmem_ram_3969, MEM_stage_inst_dmem_ram_3970, MEM_stage_inst_dmem_ram_3971, MEM_stage_inst_dmem_ram_3972, MEM_stage_inst_dmem_ram_3973, MEM_stage_inst_dmem_ram_3974, MEM_stage_inst_dmem_ram_3975, MEM_stage_inst_dmem_ram_3976, MEM_stage_inst_dmem_ram_3977, MEM_stage_inst_dmem_ram_3978, MEM_stage_inst_dmem_ram_3979, MEM_stage_inst_dmem_ram_3980, MEM_stage_inst_dmem_ram_3981, MEM_stage_inst_dmem_ram_3982, MEM_stage_inst_dmem_ram_3983, MEM_stage_inst_dmem_ram_3984, MEM_stage_inst_dmem_ram_3985, MEM_stage_inst_dmem_ram_3986, MEM_stage_inst_dmem_ram_3987, MEM_stage_inst_dmem_ram_3988, MEM_stage_inst_dmem_ram_3989, MEM_stage_inst_dmem_ram_3990, MEM_stage_inst_dmem_ram_3991, MEM_stage_inst_dmem_ram_3992, MEM_stage_inst_dmem_ram_3993, MEM_stage_inst_dmem_ram_3994, MEM_stage_inst_dmem_ram_3995, MEM_stage_inst_dmem_ram_3996, MEM_stage_inst_dmem_ram_3997, MEM_stage_inst_dmem_ram_3998, MEM_stage_inst_dmem_ram_3999, MEM_stage_inst_dmem_ram_4000, MEM_stage_inst_dmem_ram_4001, MEM_stage_inst_dmem_ram_4002, MEM_stage_inst_dmem_ram_4003, MEM_stage_inst_dmem_ram_4004, MEM_stage_inst_dmem_ram_4005, MEM_stage_inst_dmem_ram_4006, MEM_stage_inst_dmem_ram_4007, MEM_stage_inst_dmem_ram_4008, MEM_stage_inst_dmem_ram_4009, MEM_stage_inst_dmem_ram_4010, MEM_stage_inst_dmem_ram_4011, MEM_stage_inst_dmem_ram_4012, MEM_stage_inst_dmem_ram_4013, MEM_stage_inst_dmem_ram_4014, MEM_stage_inst_dmem_ram_4015, MEM_stage_inst_dmem_ram_4016, MEM_stage_inst_dmem_ram_4017, MEM_stage_inst_dmem_ram_4018, MEM_stage_inst_dmem_ram_4019, MEM_stage_inst_dmem_ram_4020, MEM_stage_inst_dmem_ram_4021, MEM_stage_inst_dmem_ram_4022, MEM_stage_inst_dmem_ram_4023, MEM_stage_inst_dmem_ram_4024, MEM_stage_inst_dmem_ram_4025, MEM_stage_inst_dmem_ram_4026, MEM_stage_inst_dmem_ram_4027, MEM_stage_inst_dmem_ram_4028, MEM_stage_inst_dmem_ram_4029, MEM_stage_inst_dmem_ram_4030, MEM_stage_inst_dmem_ram_4031, MEM_stage_inst_dmem_ram_4032, MEM_stage_inst_dmem_ram_4033, MEM_stage_inst_dmem_ram_4034, MEM_stage_inst_dmem_ram_4035, MEM_stage_inst_dmem_ram_4036, MEM_stage_inst_dmem_ram_4037, MEM_stage_inst_dmem_ram_4038, MEM_stage_inst_dmem_ram_4039, MEM_stage_inst_dmem_ram_4040, MEM_stage_inst_dmem_ram_4041, MEM_stage_inst_dmem_ram_4042, MEM_stage_inst_dmem_ram_4043, MEM_stage_inst_dmem_ram_4044, MEM_stage_inst_dmem_ram_4045, MEM_stage_inst_dmem_ram_4046, MEM_stage_inst_dmem_ram_4047, MEM_stage_inst_dmem_ram_4048, MEM_stage_inst_dmem_ram_4049, MEM_stage_inst_dmem_ram_4050, MEM_stage_inst_dmem_ram_4051, MEM_stage_inst_dmem_ram_4052, MEM_stage_inst_dmem_ram_4053, MEM_stage_inst_dmem_ram_4054, MEM_stage_inst_dmem_ram_4055, MEM_stage_inst_dmem_ram_4056, MEM_stage_inst_dmem_ram_4057, MEM_stage_inst_dmem_ram_4058, MEM_stage_inst_dmem_ram_4059, MEM_stage_inst_dmem_ram_4060, MEM_stage_inst_dmem_ram_4061, MEM_stage_inst_dmem_ram_4062, MEM_stage_inst_dmem_ram_4063, MEM_stage_inst_dmem_ram_4064, MEM_stage_inst_dmem_ram_4065, MEM_stage_inst_dmem_ram_4066, MEM_stage_inst_dmem_ram_4067, MEM_stage_inst_dmem_ram_4068, MEM_stage_inst_dmem_ram_4069, MEM_stage_inst_dmem_ram_4070, MEM_stage_inst_dmem_ram_4071, MEM_stage_inst_dmem_ram_4072, MEM_stage_inst_dmem_ram_4073, MEM_stage_inst_dmem_ram_4074, MEM_stage_inst_dmem_ram_4075, MEM_stage_inst_dmem_ram_4076, MEM_stage_inst_dmem_ram_4077, MEM_stage_inst_dmem_ram_4078, MEM_stage_inst_dmem_ram_4079, MEM_stage_inst_dmem_ram_4080, MEM_stage_inst_dmem_ram_4081, MEM_stage_inst_dmem_ram_4082, MEM_stage_inst_dmem_ram_4083, MEM_stage_inst_dmem_ram_4084, MEM_stage_inst_dmem_ram_4085, MEM_stage_inst_dmem_ram_4086, MEM_stage_inst_dmem_ram_4087, MEM_stage_inst_dmem_ram_4088, MEM_stage_inst_dmem_ram_4089, MEM_stage_inst_dmem_ram_4090, MEM_stage_inst_dmem_ram_4091, MEM_stage_inst_dmem_ram_4092, MEM_stage_inst_dmem_ram_4093, MEM_stage_inst_dmem_ram_4094, MEM_stage_inst_dmem_ram_4095, MEM_stage_inst_dmem_ram_3072, MEM_stage_inst_dmem_ram_3073, MEM_stage_inst_dmem_ram_3074, MEM_stage_inst_dmem_ram_3075, MEM_stage_inst_dmem_ram_3076, MEM_stage_inst_dmem_ram_3077, MEM_stage_inst_dmem_ram_3078, MEM_stage_inst_dmem_ram_3079, MEM_stage_inst_dmem_ram_3080, MEM_stage_inst_dmem_ram_3081, MEM_stage_inst_dmem_ram_3082, MEM_stage_inst_dmem_ram_3083, MEM_stage_inst_dmem_ram_3084, MEM_stage_inst_dmem_ram_3085, MEM_stage_inst_dmem_ram_3086, MEM_stage_inst_dmem_ram_3087, MEM_stage_inst_dmem_ram_3088, MEM_stage_inst_dmem_ram_3089, MEM_stage_inst_dmem_ram_3090, MEM_stage_inst_dmem_ram_3091, MEM_stage_inst_dmem_ram_3092, MEM_stage_inst_dmem_ram_3093, MEM_stage_inst_dmem_ram_3094, MEM_stage_inst_dmem_ram_3095, MEM_stage_inst_dmem_ram_3096, MEM_stage_inst_dmem_ram_3097, MEM_stage_inst_dmem_ram_3098, MEM_stage_inst_dmem_ram_3099, MEM_stage_inst_dmem_ram_3100, MEM_stage_inst_dmem_ram_3101, MEM_stage_inst_dmem_ram_3102, MEM_stage_inst_dmem_ram_3103, MEM_stage_inst_dmem_ram_3104, MEM_stage_inst_dmem_ram_3105, MEM_stage_inst_dmem_ram_3106, MEM_stage_inst_dmem_ram_3107, MEM_stage_inst_dmem_ram_3108, MEM_stage_inst_dmem_ram_3109, MEM_stage_inst_dmem_ram_3110, MEM_stage_inst_dmem_ram_3111, MEM_stage_inst_dmem_ram_3112, MEM_stage_inst_dmem_ram_3113, MEM_stage_inst_dmem_ram_3114, MEM_stage_inst_dmem_ram_3115, MEM_stage_inst_dmem_ram_3116, MEM_stage_inst_dmem_ram_3117, MEM_stage_inst_dmem_ram_3118, MEM_stage_inst_dmem_ram_3119, MEM_stage_inst_dmem_ram_3120, MEM_stage_inst_dmem_ram_3121, MEM_stage_inst_dmem_ram_3122, MEM_stage_inst_dmem_ram_3123, MEM_stage_inst_dmem_ram_3124, MEM_stage_inst_dmem_ram_3125, MEM_stage_inst_dmem_ram_3126, MEM_stage_inst_dmem_ram_3127, MEM_stage_inst_dmem_ram_3128, MEM_stage_inst_dmem_ram_3129, MEM_stage_inst_dmem_ram_3130, MEM_stage_inst_dmem_ram_3131, MEM_stage_inst_dmem_ram_3132, MEM_stage_inst_dmem_ram_3133, MEM_stage_inst_dmem_ram_3134, MEM_stage_inst_dmem_ram_3135, MEM_stage_inst_dmem_ram_3136, MEM_stage_inst_dmem_ram_3137, MEM_stage_inst_dmem_ram_3138, MEM_stage_inst_dmem_ram_3139, MEM_stage_inst_dmem_ram_3140, MEM_stage_inst_dmem_ram_3141, MEM_stage_inst_dmem_ram_3142, MEM_stage_inst_dmem_ram_3143, MEM_stage_inst_dmem_ram_3144, MEM_stage_inst_dmem_ram_3145, MEM_stage_inst_dmem_ram_3146, MEM_stage_inst_dmem_ram_3147, MEM_stage_inst_dmem_ram_3148, MEM_stage_inst_dmem_ram_3149, MEM_stage_inst_dmem_ram_3150, MEM_stage_inst_dmem_ram_3151, MEM_stage_inst_dmem_ram_3152, MEM_stage_inst_dmem_ram_3153, MEM_stage_inst_dmem_ram_3154, MEM_stage_inst_dmem_ram_3155, MEM_stage_inst_dmem_ram_3156, MEM_stage_inst_dmem_ram_3157, MEM_stage_inst_dmem_ram_3158, MEM_stage_inst_dmem_ram_3159, MEM_stage_inst_dmem_ram_3160, MEM_stage_inst_dmem_ram_3161, MEM_stage_inst_dmem_ram_3162, MEM_stage_inst_dmem_ram_3163, MEM_stage_inst_dmem_ram_3164, MEM_stage_inst_dmem_ram_3165, MEM_stage_inst_dmem_ram_3166, MEM_stage_inst_dmem_ram_3167, MEM_stage_inst_dmem_ram_3168, MEM_stage_inst_dmem_ram_3169, MEM_stage_inst_dmem_ram_3170, MEM_stage_inst_dmem_ram_3171, MEM_stage_inst_dmem_ram_3172, MEM_stage_inst_dmem_ram_3173, MEM_stage_inst_dmem_ram_3174, MEM_stage_inst_dmem_ram_3175, MEM_stage_inst_dmem_ram_3176, MEM_stage_inst_dmem_ram_3177, MEM_stage_inst_dmem_ram_3178, MEM_stage_inst_dmem_ram_3179, MEM_stage_inst_dmem_ram_3180, MEM_stage_inst_dmem_ram_3181, MEM_stage_inst_dmem_ram_3182, MEM_stage_inst_dmem_ram_3183, MEM_stage_inst_dmem_ram_3184, MEM_stage_inst_dmem_ram_3185, MEM_stage_inst_dmem_ram_3186, MEM_stage_inst_dmem_ram_3187, MEM_stage_inst_dmem_ram_3188, MEM_stage_inst_dmem_ram_3189, MEM_stage_inst_dmem_ram_3190, MEM_stage_inst_dmem_ram_3191, MEM_stage_inst_dmem_ram_3192, MEM_stage_inst_dmem_ram_3193, MEM_stage_inst_dmem_ram_3194, MEM_stage_inst_dmem_ram_3195, MEM_stage_inst_dmem_ram_3196, MEM_stage_inst_dmem_ram_3197, MEM_stage_inst_dmem_ram_3198, MEM_stage_inst_dmem_ram_3199, MEM_stage_inst_dmem_ram_3200, MEM_stage_inst_dmem_ram_3201, MEM_stage_inst_dmem_ram_3202, MEM_stage_inst_dmem_ram_3203, MEM_stage_inst_dmem_ram_3204, MEM_stage_inst_dmem_ram_3205, MEM_stage_inst_dmem_ram_3206, MEM_stage_inst_dmem_ram_3207, MEM_stage_inst_dmem_ram_3208, MEM_stage_inst_dmem_ram_3209, MEM_stage_inst_dmem_ram_3210, MEM_stage_inst_dmem_ram_3211, MEM_stage_inst_dmem_ram_3212, MEM_stage_inst_dmem_ram_3213, MEM_stage_inst_dmem_ram_3214, MEM_stage_inst_dmem_ram_3215, MEM_stage_inst_dmem_ram_3216, MEM_stage_inst_dmem_ram_3217, MEM_stage_inst_dmem_ram_3218, MEM_stage_inst_dmem_ram_3219, MEM_stage_inst_dmem_ram_3220, MEM_stage_inst_dmem_ram_3221, MEM_stage_inst_dmem_ram_3222, MEM_stage_inst_dmem_ram_3223, MEM_stage_inst_dmem_ram_3224, MEM_stage_inst_dmem_ram_3225, MEM_stage_inst_dmem_ram_3226, MEM_stage_inst_dmem_ram_3227, MEM_stage_inst_dmem_ram_3228, MEM_stage_inst_dmem_ram_3229, MEM_stage_inst_dmem_ram_3230, MEM_stage_inst_dmem_ram_3231, MEM_stage_inst_dmem_ram_3232, MEM_stage_inst_dmem_ram_3233, MEM_stage_inst_dmem_ram_3234, MEM_stage_inst_dmem_ram_3235, MEM_stage_inst_dmem_ram_3236, MEM_stage_inst_dmem_ram_3237, MEM_stage_inst_dmem_ram_3238, MEM_stage_inst_dmem_ram_3239, MEM_stage_inst_dmem_ram_3240, MEM_stage_inst_dmem_ram_3241, MEM_stage_inst_dmem_ram_3242, MEM_stage_inst_dmem_ram_3243, MEM_stage_inst_dmem_ram_3244, MEM_stage_inst_dmem_ram_3245, MEM_stage_inst_dmem_ram_3246, MEM_stage_inst_dmem_ram_3247, MEM_stage_inst_dmem_ram_3248, MEM_stage_inst_dmem_ram_3249, MEM_stage_inst_dmem_ram_3250, MEM_stage_inst_dmem_ram_3251, MEM_stage_inst_dmem_ram_3252, MEM_stage_inst_dmem_ram_3253, MEM_stage_inst_dmem_ram_3254, MEM_stage_inst_dmem_ram_3255, MEM_stage_inst_dmem_ram_3256, MEM_stage_inst_dmem_ram_3257, MEM_stage_inst_dmem_ram_3258, MEM_stage_inst_dmem_ram_3259, MEM_stage_inst_dmem_ram_3260, MEM_stage_inst_dmem_ram_3261, MEM_stage_inst_dmem_ram_3262, MEM_stage_inst_dmem_ram_3263, MEM_stage_inst_dmem_ram_3264, MEM_stage_inst_dmem_ram_3265, MEM_stage_inst_dmem_ram_3266, MEM_stage_inst_dmem_ram_3267, MEM_stage_inst_dmem_ram_3268, MEM_stage_inst_dmem_ram_3269, MEM_stage_inst_dmem_ram_3270, MEM_stage_inst_dmem_ram_3271, MEM_stage_inst_dmem_ram_3272, MEM_stage_inst_dmem_ram_3273, MEM_stage_inst_dmem_ram_3274, MEM_stage_inst_dmem_ram_3275, MEM_stage_inst_dmem_ram_3276, MEM_stage_inst_dmem_ram_3277, MEM_stage_inst_dmem_ram_3278, MEM_stage_inst_dmem_ram_3279, MEM_stage_inst_dmem_ram_3280, MEM_stage_inst_dmem_ram_3281, MEM_stage_inst_dmem_ram_3282, MEM_stage_inst_dmem_ram_3283, MEM_stage_inst_dmem_ram_3284, MEM_stage_inst_dmem_ram_3285, MEM_stage_inst_dmem_ram_3286, MEM_stage_inst_dmem_ram_3287, MEM_stage_inst_dmem_ram_3288, MEM_stage_inst_dmem_ram_3289, MEM_stage_inst_dmem_ram_3290, MEM_stage_inst_dmem_ram_3291, MEM_stage_inst_dmem_ram_3292, MEM_stage_inst_dmem_ram_3293, MEM_stage_inst_dmem_ram_3294, MEM_stage_inst_dmem_ram_3295, MEM_stage_inst_dmem_ram_3296, MEM_stage_inst_dmem_ram_3297, MEM_stage_inst_dmem_ram_3298, MEM_stage_inst_dmem_ram_3299, MEM_stage_inst_dmem_ram_3300, MEM_stage_inst_dmem_ram_3301, MEM_stage_inst_dmem_ram_3302, MEM_stage_inst_dmem_ram_3303, MEM_stage_inst_dmem_ram_3304, MEM_stage_inst_dmem_ram_3305, MEM_stage_inst_dmem_ram_3306, MEM_stage_inst_dmem_ram_3307, MEM_stage_inst_dmem_ram_3308, MEM_stage_inst_dmem_ram_3309, MEM_stage_inst_dmem_ram_3310, MEM_stage_inst_dmem_ram_3311, MEM_stage_inst_dmem_ram_3312, MEM_stage_inst_dmem_ram_3313, MEM_stage_inst_dmem_ram_3314, MEM_stage_inst_dmem_ram_3315, MEM_stage_inst_dmem_ram_3316, MEM_stage_inst_dmem_ram_3317, MEM_stage_inst_dmem_ram_3318, MEM_stage_inst_dmem_ram_3319, MEM_stage_inst_dmem_ram_3320, MEM_stage_inst_dmem_ram_3321, MEM_stage_inst_dmem_ram_3322, MEM_stage_inst_dmem_ram_3323, MEM_stage_inst_dmem_ram_3324, MEM_stage_inst_dmem_ram_3325, MEM_stage_inst_dmem_ram_3326, MEM_stage_inst_dmem_ram_3327, MEM_stage_inst_dmem_ram_3328, MEM_stage_inst_dmem_ram_3329, MEM_stage_inst_dmem_ram_3330, MEM_stage_inst_dmem_ram_3331, MEM_stage_inst_dmem_ram_3332, MEM_stage_inst_dmem_ram_3333, MEM_stage_inst_dmem_ram_3334, MEM_stage_inst_dmem_ram_3335, MEM_stage_inst_dmem_ram_3336, MEM_stage_inst_dmem_ram_3337, MEM_stage_inst_dmem_ram_3338, MEM_stage_inst_dmem_ram_3339, MEM_stage_inst_dmem_ram_3340, MEM_stage_inst_dmem_ram_3341, MEM_stage_inst_dmem_ram_3342, MEM_stage_inst_dmem_ram_3343, MEM_stage_inst_dmem_ram_3344, MEM_stage_inst_dmem_ram_3345, MEM_stage_inst_dmem_ram_3346, MEM_stage_inst_dmem_ram_3347, MEM_stage_inst_dmem_ram_3348, MEM_stage_inst_dmem_ram_3349, MEM_stage_inst_dmem_ram_3350, MEM_stage_inst_dmem_ram_3351, MEM_stage_inst_dmem_ram_3352, MEM_stage_inst_dmem_ram_3353, MEM_stage_inst_dmem_ram_3354, MEM_stage_inst_dmem_ram_3355, MEM_stage_inst_dmem_ram_3356, MEM_stage_inst_dmem_ram_3357, MEM_stage_inst_dmem_ram_3358, MEM_stage_inst_dmem_ram_3359, MEM_stage_inst_dmem_ram_3360, MEM_stage_inst_dmem_ram_3361, MEM_stage_inst_dmem_ram_3362, MEM_stage_inst_dmem_ram_3363, MEM_stage_inst_dmem_ram_3364, MEM_stage_inst_dmem_ram_3365, MEM_stage_inst_dmem_ram_3366, MEM_stage_inst_dmem_ram_3367, MEM_stage_inst_dmem_ram_3368, MEM_stage_inst_dmem_ram_3369, MEM_stage_inst_dmem_ram_3370, MEM_stage_inst_dmem_ram_3371, MEM_stage_inst_dmem_ram_3372, MEM_stage_inst_dmem_ram_3373, MEM_stage_inst_dmem_ram_3374, MEM_stage_inst_dmem_ram_3375, MEM_stage_inst_dmem_ram_3376, MEM_stage_inst_dmem_ram_3377, MEM_stage_inst_dmem_ram_3378, MEM_stage_inst_dmem_ram_3379, MEM_stage_inst_dmem_ram_3380, MEM_stage_inst_dmem_ram_3381, MEM_stage_inst_dmem_ram_3382, MEM_stage_inst_dmem_ram_3383, MEM_stage_inst_dmem_ram_3384, MEM_stage_inst_dmem_ram_3385, MEM_stage_inst_dmem_ram_3386, MEM_stage_inst_dmem_ram_3387, MEM_stage_inst_dmem_ram_3388, MEM_stage_inst_dmem_ram_3389, MEM_stage_inst_dmem_ram_3390, MEM_stage_inst_dmem_ram_3391, MEM_stage_inst_dmem_ram_3392, MEM_stage_inst_dmem_ram_3393, MEM_stage_inst_dmem_ram_3394, MEM_stage_inst_dmem_ram_3395, MEM_stage_inst_dmem_ram_3396, MEM_stage_inst_dmem_ram_3397, MEM_stage_inst_dmem_ram_3398, MEM_stage_inst_dmem_ram_3399, MEM_stage_inst_dmem_ram_3400, MEM_stage_inst_dmem_ram_3401, MEM_stage_inst_dmem_ram_3402, MEM_stage_inst_dmem_ram_3403, MEM_stage_inst_dmem_ram_3404, MEM_stage_inst_dmem_ram_3405, MEM_stage_inst_dmem_ram_3406, MEM_stage_inst_dmem_ram_3407, MEM_stage_inst_dmem_ram_3408, MEM_stage_inst_dmem_ram_3409, MEM_stage_inst_dmem_ram_3410, MEM_stage_inst_dmem_ram_3411, MEM_stage_inst_dmem_ram_3412, MEM_stage_inst_dmem_ram_3413, MEM_stage_inst_dmem_ram_3414, MEM_stage_inst_dmem_ram_3415, MEM_stage_inst_dmem_ram_3416, MEM_stage_inst_dmem_ram_3417, MEM_stage_inst_dmem_ram_3418, MEM_stage_inst_dmem_ram_3419, MEM_stage_inst_dmem_ram_3420, MEM_stage_inst_dmem_ram_3421, MEM_stage_inst_dmem_ram_3422, MEM_stage_inst_dmem_ram_3423, MEM_stage_inst_dmem_ram_3424, MEM_stage_inst_dmem_ram_3425, MEM_stage_inst_dmem_ram_3426, MEM_stage_inst_dmem_ram_3427, MEM_stage_inst_dmem_ram_3428, MEM_stage_inst_dmem_ram_3429, MEM_stage_inst_dmem_ram_3430, MEM_stage_inst_dmem_ram_3431, MEM_stage_inst_dmem_ram_3432, MEM_stage_inst_dmem_ram_3433, MEM_stage_inst_dmem_ram_3434, MEM_stage_inst_dmem_ram_3435, MEM_stage_inst_dmem_ram_3436, MEM_stage_inst_dmem_ram_3437, MEM_stage_inst_dmem_ram_3438, MEM_stage_inst_dmem_ram_3439, MEM_stage_inst_dmem_ram_3440, MEM_stage_inst_dmem_ram_3441, MEM_stage_inst_dmem_ram_3442, MEM_stage_inst_dmem_ram_3443, MEM_stage_inst_dmem_ram_3444, MEM_stage_inst_dmem_ram_3445, MEM_stage_inst_dmem_ram_3446, MEM_stage_inst_dmem_ram_3447, MEM_stage_inst_dmem_ram_3448, MEM_stage_inst_dmem_ram_3449, MEM_stage_inst_dmem_ram_3450, MEM_stage_inst_dmem_ram_3451, MEM_stage_inst_dmem_ram_3452, MEM_stage_inst_dmem_ram_3453, MEM_stage_inst_dmem_ram_3454, MEM_stage_inst_dmem_ram_3455, MEM_stage_inst_dmem_ram_3456, MEM_stage_inst_dmem_ram_3457, MEM_stage_inst_dmem_ram_3458, MEM_stage_inst_dmem_ram_3459, MEM_stage_inst_dmem_ram_3460, MEM_stage_inst_dmem_ram_3461, MEM_stage_inst_dmem_ram_3462, MEM_stage_inst_dmem_ram_3463, MEM_stage_inst_dmem_ram_3464, MEM_stage_inst_dmem_ram_3465, MEM_stage_inst_dmem_ram_3466, MEM_stage_inst_dmem_ram_3467, MEM_stage_inst_dmem_ram_3468, MEM_stage_inst_dmem_ram_3469, MEM_stage_inst_dmem_ram_3470, MEM_stage_inst_dmem_ram_3471, MEM_stage_inst_dmem_ram_3472, MEM_stage_inst_dmem_ram_3473, MEM_stage_inst_dmem_ram_3474, MEM_stage_inst_dmem_ram_3475, MEM_stage_inst_dmem_ram_3476, MEM_stage_inst_dmem_ram_3477, MEM_stage_inst_dmem_ram_3478, MEM_stage_inst_dmem_ram_3479, MEM_stage_inst_dmem_ram_3480, MEM_stage_inst_dmem_ram_3481, MEM_stage_inst_dmem_ram_3482, MEM_stage_inst_dmem_ram_3483, MEM_stage_inst_dmem_ram_3484, MEM_stage_inst_dmem_ram_3485, MEM_stage_inst_dmem_ram_3486, MEM_stage_inst_dmem_ram_3487, MEM_stage_inst_dmem_ram_3488, MEM_stage_inst_dmem_ram_3489, MEM_stage_inst_dmem_ram_3490, MEM_stage_inst_dmem_ram_3491, MEM_stage_inst_dmem_ram_3492, MEM_stage_inst_dmem_ram_3493, MEM_stage_inst_dmem_ram_3494, MEM_stage_inst_dmem_ram_3495, MEM_stage_inst_dmem_ram_3496, MEM_stage_inst_dmem_ram_3497, MEM_stage_inst_dmem_ram_3498, MEM_stage_inst_dmem_ram_3499, MEM_stage_inst_dmem_ram_3500, MEM_stage_inst_dmem_ram_3501, MEM_stage_inst_dmem_ram_3502, MEM_stage_inst_dmem_ram_3503, MEM_stage_inst_dmem_ram_3504, MEM_stage_inst_dmem_ram_3505, MEM_stage_inst_dmem_ram_3506, MEM_stage_inst_dmem_ram_3507, MEM_stage_inst_dmem_ram_3508, MEM_stage_inst_dmem_ram_3509, MEM_stage_inst_dmem_ram_3510, MEM_stage_inst_dmem_ram_3511, MEM_stage_inst_dmem_ram_3512, MEM_stage_inst_dmem_ram_3513, MEM_stage_inst_dmem_ram_3514, MEM_stage_inst_dmem_ram_3515, MEM_stage_inst_dmem_ram_3516, MEM_stage_inst_dmem_ram_3517, MEM_stage_inst_dmem_ram_3518, MEM_stage_inst_dmem_ram_3519, MEM_stage_inst_dmem_ram_3520, MEM_stage_inst_dmem_ram_3521, MEM_stage_inst_dmem_ram_3522, MEM_stage_inst_dmem_ram_3523, MEM_stage_inst_dmem_ram_3524, MEM_stage_inst_dmem_ram_3525, MEM_stage_inst_dmem_ram_3526, MEM_stage_inst_dmem_ram_3527, MEM_stage_inst_dmem_ram_3528, MEM_stage_inst_dmem_ram_3529, MEM_stage_inst_dmem_ram_3530, MEM_stage_inst_dmem_ram_3531, MEM_stage_inst_dmem_ram_3532, MEM_stage_inst_dmem_ram_3533, MEM_stage_inst_dmem_ram_3534, MEM_stage_inst_dmem_ram_3535, MEM_stage_inst_dmem_ram_3536, MEM_stage_inst_dmem_ram_3537, MEM_stage_inst_dmem_ram_3538, MEM_stage_inst_dmem_ram_3539, MEM_stage_inst_dmem_ram_3540, MEM_stage_inst_dmem_ram_3541, MEM_stage_inst_dmem_ram_3542, MEM_stage_inst_dmem_ram_3543, MEM_stage_inst_dmem_ram_3544, MEM_stage_inst_dmem_ram_3545, MEM_stage_inst_dmem_ram_3546, MEM_stage_inst_dmem_ram_3547, MEM_stage_inst_dmem_ram_3548, MEM_stage_inst_dmem_ram_3549, MEM_stage_inst_dmem_ram_3550, MEM_stage_inst_dmem_ram_3551, MEM_stage_inst_dmem_ram_3552, MEM_stage_inst_dmem_ram_3553, MEM_stage_inst_dmem_ram_3554, MEM_stage_inst_dmem_ram_3555, MEM_stage_inst_dmem_ram_3556, MEM_stage_inst_dmem_ram_3557, MEM_stage_inst_dmem_ram_3558, MEM_stage_inst_dmem_ram_3559, MEM_stage_inst_dmem_ram_3560, MEM_stage_inst_dmem_ram_3561, MEM_stage_inst_dmem_ram_3562, MEM_stage_inst_dmem_ram_3563, MEM_stage_inst_dmem_ram_3564, MEM_stage_inst_dmem_ram_3565, MEM_stage_inst_dmem_ram_3566, MEM_stage_inst_dmem_ram_3567, MEM_stage_inst_dmem_ram_3568, MEM_stage_inst_dmem_ram_3569, MEM_stage_inst_dmem_ram_3570, MEM_stage_inst_dmem_ram_3571, MEM_stage_inst_dmem_ram_3572, MEM_stage_inst_dmem_ram_3573, MEM_stage_inst_dmem_ram_3574, MEM_stage_inst_dmem_ram_3575, MEM_stage_inst_dmem_ram_3576, MEM_stage_inst_dmem_ram_3577, MEM_stage_inst_dmem_ram_3578, MEM_stage_inst_dmem_ram_3579, MEM_stage_inst_dmem_ram_3580, MEM_stage_inst_dmem_ram_3581, MEM_stage_inst_dmem_ram_3582, MEM_stage_inst_dmem_ram_3583, MEM_stage_inst_dmem_ram_2560, MEM_stage_inst_dmem_ram_2561, MEM_stage_inst_dmem_ram_2562, MEM_stage_inst_dmem_ram_2563, MEM_stage_inst_dmem_ram_2564, MEM_stage_inst_dmem_ram_2565, MEM_stage_inst_dmem_ram_2566, MEM_stage_inst_dmem_ram_2567, MEM_stage_inst_dmem_ram_2568, MEM_stage_inst_dmem_ram_2569, MEM_stage_inst_dmem_ram_2570, MEM_stage_inst_dmem_ram_2571, MEM_stage_inst_dmem_ram_2572, MEM_stage_inst_dmem_ram_2573, MEM_stage_inst_dmem_ram_2574, MEM_stage_inst_dmem_ram_2575, MEM_stage_inst_dmem_ram_2576, MEM_stage_inst_dmem_ram_2577, MEM_stage_inst_dmem_ram_2578, MEM_stage_inst_dmem_ram_2579, MEM_stage_inst_dmem_ram_2580, MEM_stage_inst_dmem_ram_2581, MEM_stage_inst_dmem_ram_2582, MEM_stage_inst_dmem_ram_2583, MEM_stage_inst_dmem_ram_2584, MEM_stage_inst_dmem_ram_2585, MEM_stage_inst_dmem_ram_2586, MEM_stage_inst_dmem_ram_2587, MEM_stage_inst_dmem_ram_2588, MEM_stage_inst_dmem_ram_2589, MEM_stage_inst_dmem_ram_2590, MEM_stage_inst_dmem_ram_2591, MEM_stage_inst_dmem_ram_2592, MEM_stage_inst_dmem_ram_2593, MEM_stage_inst_dmem_ram_2594, MEM_stage_inst_dmem_ram_2595, MEM_stage_inst_dmem_ram_2596, MEM_stage_inst_dmem_ram_2597, MEM_stage_inst_dmem_ram_2598, MEM_stage_inst_dmem_ram_2599, MEM_stage_inst_dmem_ram_2600, MEM_stage_inst_dmem_ram_2601, MEM_stage_inst_dmem_ram_2602, MEM_stage_inst_dmem_ram_2603, MEM_stage_inst_dmem_ram_2604, MEM_stage_inst_dmem_ram_2605, MEM_stage_inst_dmem_ram_2606, MEM_stage_inst_dmem_ram_2607, MEM_stage_inst_dmem_ram_2608, MEM_stage_inst_dmem_ram_2609, MEM_stage_inst_dmem_ram_2610, MEM_stage_inst_dmem_ram_2611, MEM_stage_inst_dmem_ram_2612, MEM_stage_inst_dmem_ram_2613, MEM_stage_inst_dmem_ram_2614, MEM_stage_inst_dmem_ram_2615, MEM_stage_inst_dmem_ram_2616, MEM_stage_inst_dmem_ram_2617, MEM_stage_inst_dmem_ram_2618, MEM_stage_inst_dmem_ram_2619, MEM_stage_inst_dmem_ram_2620, MEM_stage_inst_dmem_ram_2621, MEM_stage_inst_dmem_ram_2622, MEM_stage_inst_dmem_ram_2623, MEM_stage_inst_dmem_ram_2624, MEM_stage_inst_dmem_ram_2625, MEM_stage_inst_dmem_ram_2626, MEM_stage_inst_dmem_ram_2627, MEM_stage_inst_dmem_ram_2628, MEM_stage_inst_dmem_ram_2629, MEM_stage_inst_dmem_ram_2630, MEM_stage_inst_dmem_ram_2631, MEM_stage_inst_dmem_ram_2632, MEM_stage_inst_dmem_ram_2633, MEM_stage_inst_dmem_ram_2634, MEM_stage_inst_dmem_ram_2635, MEM_stage_inst_dmem_ram_2636, MEM_stage_inst_dmem_ram_2637, MEM_stage_inst_dmem_ram_2638, MEM_stage_inst_dmem_ram_2639, MEM_stage_inst_dmem_ram_2640, MEM_stage_inst_dmem_ram_2641, MEM_stage_inst_dmem_ram_2642, MEM_stage_inst_dmem_ram_2643, MEM_stage_inst_dmem_ram_2644, MEM_stage_inst_dmem_ram_2645, MEM_stage_inst_dmem_ram_2646, MEM_stage_inst_dmem_ram_2647, MEM_stage_inst_dmem_ram_2648, MEM_stage_inst_dmem_ram_2649, MEM_stage_inst_dmem_ram_2650, MEM_stage_inst_dmem_ram_2651, MEM_stage_inst_dmem_ram_2652, MEM_stage_inst_dmem_ram_2653, MEM_stage_inst_dmem_ram_2654, MEM_stage_inst_dmem_ram_2655, MEM_stage_inst_dmem_ram_2656, MEM_stage_inst_dmem_ram_2657, MEM_stage_inst_dmem_ram_2658, MEM_stage_inst_dmem_ram_2659, MEM_stage_inst_dmem_ram_2660, MEM_stage_inst_dmem_ram_2661, MEM_stage_inst_dmem_ram_2662, MEM_stage_inst_dmem_ram_2663, MEM_stage_inst_dmem_ram_2664, MEM_stage_inst_dmem_ram_2665, MEM_stage_inst_dmem_ram_2666, MEM_stage_inst_dmem_ram_2667, MEM_stage_inst_dmem_ram_2668, MEM_stage_inst_dmem_ram_2669, MEM_stage_inst_dmem_ram_2670, MEM_stage_inst_dmem_ram_2671, MEM_stage_inst_dmem_ram_2672, MEM_stage_inst_dmem_ram_2673, MEM_stage_inst_dmem_ram_2674, MEM_stage_inst_dmem_ram_2675, MEM_stage_inst_dmem_ram_2676, MEM_stage_inst_dmem_ram_2677, MEM_stage_inst_dmem_ram_2678, MEM_stage_inst_dmem_ram_2679, MEM_stage_inst_dmem_ram_2680, MEM_stage_inst_dmem_ram_2681, MEM_stage_inst_dmem_ram_2682, MEM_stage_inst_dmem_ram_2683, MEM_stage_inst_dmem_ram_2684, MEM_stage_inst_dmem_ram_2685, MEM_stage_inst_dmem_ram_2686, MEM_stage_inst_dmem_ram_2687, MEM_stage_inst_dmem_ram_2688, MEM_stage_inst_dmem_ram_2689, MEM_stage_inst_dmem_ram_2690, MEM_stage_inst_dmem_ram_2691, MEM_stage_inst_dmem_ram_2692, MEM_stage_inst_dmem_ram_2693, MEM_stage_inst_dmem_ram_2694, MEM_stage_inst_dmem_ram_2695, MEM_stage_inst_dmem_ram_2696, MEM_stage_inst_dmem_ram_2697, MEM_stage_inst_dmem_ram_2698, MEM_stage_inst_dmem_ram_2699, MEM_stage_inst_dmem_ram_2700, MEM_stage_inst_dmem_ram_2701, MEM_stage_inst_dmem_ram_2702, MEM_stage_inst_dmem_ram_2703, MEM_stage_inst_dmem_ram_2704, MEM_stage_inst_dmem_ram_2705, MEM_stage_inst_dmem_ram_2706, MEM_stage_inst_dmem_ram_2707, MEM_stage_inst_dmem_ram_2708, MEM_stage_inst_dmem_ram_2709, MEM_stage_inst_dmem_ram_2710, MEM_stage_inst_dmem_ram_2711, MEM_stage_inst_dmem_ram_2712, MEM_stage_inst_dmem_ram_2713, MEM_stage_inst_dmem_ram_2714, MEM_stage_inst_dmem_ram_2715, MEM_stage_inst_dmem_ram_2716, MEM_stage_inst_dmem_ram_2717, MEM_stage_inst_dmem_ram_2718, MEM_stage_inst_dmem_ram_2719, MEM_stage_inst_dmem_ram_2720, MEM_stage_inst_dmem_ram_2721, MEM_stage_inst_dmem_ram_2722, MEM_stage_inst_dmem_ram_2723, MEM_stage_inst_dmem_ram_2724, MEM_stage_inst_dmem_ram_2725, MEM_stage_inst_dmem_ram_2726, MEM_stage_inst_dmem_ram_2727, MEM_stage_inst_dmem_ram_2728, MEM_stage_inst_dmem_ram_2729, MEM_stage_inst_dmem_ram_2730, MEM_stage_inst_dmem_ram_2731, MEM_stage_inst_dmem_ram_2732, MEM_stage_inst_dmem_ram_2733, MEM_stage_inst_dmem_ram_2734, MEM_stage_inst_dmem_ram_2735, MEM_stage_inst_dmem_ram_2736, MEM_stage_inst_dmem_ram_2737, MEM_stage_inst_dmem_ram_2738, MEM_stage_inst_dmem_ram_2739, MEM_stage_inst_dmem_ram_2740, MEM_stage_inst_dmem_ram_2741, MEM_stage_inst_dmem_ram_2742, MEM_stage_inst_dmem_ram_2743, MEM_stage_inst_dmem_ram_2744, MEM_stage_inst_dmem_ram_2745, MEM_stage_inst_dmem_ram_2746, MEM_stage_inst_dmem_ram_2747, MEM_stage_inst_dmem_ram_2748, MEM_stage_inst_dmem_ram_2749, MEM_stage_inst_dmem_ram_2750, MEM_stage_inst_dmem_ram_2751, MEM_stage_inst_dmem_ram_2752, MEM_stage_inst_dmem_ram_2753, MEM_stage_inst_dmem_ram_2754, MEM_stage_inst_dmem_ram_2755, MEM_stage_inst_dmem_ram_2756, MEM_stage_inst_dmem_ram_2757, MEM_stage_inst_dmem_ram_2758, MEM_stage_inst_dmem_ram_2759, MEM_stage_inst_dmem_ram_2760, MEM_stage_inst_dmem_ram_2761, MEM_stage_inst_dmem_ram_2762, MEM_stage_inst_dmem_ram_2763, MEM_stage_inst_dmem_ram_2764, MEM_stage_inst_dmem_ram_2765, MEM_stage_inst_dmem_ram_2766, MEM_stage_inst_dmem_ram_2767, MEM_stage_inst_dmem_ram_2768, MEM_stage_inst_dmem_ram_2769, MEM_stage_inst_dmem_ram_2770, MEM_stage_inst_dmem_ram_2771, MEM_stage_inst_dmem_ram_2772, MEM_stage_inst_dmem_ram_2773, MEM_stage_inst_dmem_ram_2774, MEM_stage_inst_dmem_ram_2775, MEM_stage_inst_dmem_ram_2776, MEM_stage_inst_dmem_ram_2777, MEM_stage_inst_dmem_ram_2778, MEM_stage_inst_dmem_ram_2779, MEM_stage_inst_dmem_ram_2780, MEM_stage_inst_dmem_ram_2781, MEM_stage_inst_dmem_ram_2782, MEM_stage_inst_dmem_ram_2783, MEM_stage_inst_dmem_ram_2784, MEM_stage_inst_dmem_ram_2785, MEM_stage_inst_dmem_ram_2786, MEM_stage_inst_dmem_ram_2787, MEM_stage_inst_dmem_ram_2788, MEM_stage_inst_dmem_ram_2789, MEM_stage_inst_dmem_ram_2790, MEM_stage_inst_dmem_ram_2791, MEM_stage_inst_dmem_ram_2792, MEM_stage_inst_dmem_ram_2793, MEM_stage_inst_dmem_ram_2794, MEM_stage_inst_dmem_ram_2795, MEM_stage_inst_dmem_ram_2796, MEM_stage_inst_dmem_ram_2797, MEM_stage_inst_dmem_ram_2798, MEM_stage_inst_dmem_ram_2799, MEM_stage_inst_dmem_ram_2800, MEM_stage_inst_dmem_ram_2801, MEM_stage_inst_dmem_ram_2802, MEM_stage_inst_dmem_ram_2803, MEM_stage_inst_dmem_ram_2804, MEM_stage_inst_dmem_ram_2805, MEM_stage_inst_dmem_ram_2806, MEM_stage_inst_dmem_ram_2807, MEM_stage_inst_dmem_ram_2808, MEM_stage_inst_dmem_ram_2809, MEM_stage_inst_dmem_ram_2810, MEM_stage_inst_dmem_ram_2811, MEM_stage_inst_dmem_ram_2812, MEM_stage_inst_dmem_ram_2813, MEM_stage_inst_dmem_ram_2814, MEM_stage_inst_dmem_ram_2815, MEM_stage_inst_dmem_ram_2816, MEM_stage_inst_dmem_ram_2817, MEM_stage_inst_dmem_ram_2818, MEM_stage_inst_dmem_ram_2819, MEM_stage_inst_dmem_ram_2820, MEM_stage_inst_dmem_ram_2821, MEM_stage_inst_dmem_ram_2822, MEM_stage_inst_dmem_ram_2823, MEM_stage_inst_dmem_ram_2824, MEM_stage_inst_dmem_ram_2825, MEM_stage_inst_dmem_ram_2826, MEM_stage_inst_dmem_ram_2827, MEM_stage_inst_dmem_ram_2828, MEM_stage_inst_dmem_ram_2829, MEM_stage_inst_dmem_ram_2830, MEM_stage_inst_dmem_ram_2831, MEM_stage_inst_dmem_ram_2832, MEM_stage_inst_dmem_ram_2833, MEM_stage_inst_dmem_ram_2834, MEM_stage_inst_dmem_ram_2835, MEM_stage_inst_dmem_ram_2836, MEM_stage_inst_dmem_ram_2837, MEM_stage_inst_dmem_ram_2838, MEM_stage_inst_dmem_ram_2839, MEM_stage_inst_dmem_ram_2840, MEM_stage_inst_dmem_ram_2841, MEM_stage_inst_dmem_ram_2842, MEM_stage_inst_dmem_ram_2843, MEM_stage_inst_dmem_ram_2844, MEM_stage_inst_dmem_ram_2845, MEM_stage_inst_dmem_ram_2846, MEM_stage_inst_dmem_ram_2847, MEM_stage_inst_dmem_ram_2848, MEM_stage_inst_dmem_ram_2849, MEM_stage_inst_dmem_ram_2850, MEM_stage_inst_dmem_ram_2851, MEM_stage_inst_dmem_ram_2852, MEM_stage_inst_dmem_ram_2853, MEM_stage_inst_dmem_ram_2854, MEM_stage_inst_dmem_ram_2855, MEM_stage_inst_dmem_ram_2856, MEM_stage_inst_dmem_ram_2857, MEM_stage_inst_dmem_ram_2858, MEM_stage_inst_dmem_ram_2859, MEM_stage_inst_dmem_ram_2860, MEM_stage_inst_dmem_ram_2861, MEM_stage_inst_dmem_ram_2862, MEM_stage_inst_dmem_ram_2863, MEM_stage_inst_dmem_ram_2864, MEM_stage_inst_dmem_ram_2865, MEM_stage_inst_dmem_ram_2866, MEM_stage_inst_dmem_ram_2867, MEM_stage_inst_dmem_ram_2868, MEM_stage_inst_dmem_ram_2869, MEM_stage_inst_dmem_ram_2870, MEM_stage_inst_dmem_ram_2871, MEM_stage_inst_dmem_ram_2872, MEM_stage_inst_dmem_ram_2873, MEM_stage_inst_dmem_ram_2874, MEM_stage_inst_dmem_ram_2875, MEM_stage_inst_dmem_ram_2876, MEM_stage_inst_dmem_ram_2877, MEM_stage_inst_dmem_ram_2878, MEM_stage_inst_dmem_ram_2879, MEM_stage_inst_dmem_ram_2880, MEM_stage_inst_dmem_ram_2881, MEM_stage_inst_dmem_ram_2882, MEM_stage_inst_dmem_ram_2883, MEM_stage_inst_dmem_ram_2884, MEM_stage_inst_dmem_ram_2885, MEM_stage_inst_dmem_ram_2886, MEM_stage_inst_dmem_ram_2887, MEM_stage_inst_dmem_ram_2888, MEM_stage_inst_dmem_ram_2889, MEM_stage_inst_dmem_ram_2890, MEM_stage_inst_dmem_ram_2891, MEM_stage_inst_dmem_ram_2892, MEM_stage_inst_dmem_ram_2893, MEM_stage_inst_dmem_ram_2894, MEM_stage_inst_dmem_ram_2895, MEM_stage_inst_dmem_ram_2896, MEM_stage_inst_dmem_ram_2897, MEM_stage_inst_dmem_ram_2898, MEM_stage_inst_dmem_ram_2899, MEM_stage_inst_dmem_ram_2900, MEM_stage_inst_dmem_ram_2901, MEM_stage_inst_dmem_ram_2902, MEM_stage_inst_dmem_ram_2903, MEM_stage_inst_dmem_ram_2904, MEM_stage_inst_dmem_ram_2905, MEM_stage_inst_dmem_ram_2906, MEM_stage_inst_dmem_ram_2907, MEM_stage_inst_dmem_ram_2908, MEM_stage_inst_dmem_ram_2909, MEM_stage_inst_dmem_ram_2910, MEM_stage_inst_dmem_ram_2911, MEM_stage_inst_dmem_ram_2912, MEM_stage_inst_dmem_ram_2913, MEM_stage_inst_dmem_ram_2914, MEM_stage_inst_dmem_ram_2915, MEM_stage_inst_dmem_ram_2916, MEM_stage_inst_dmem_ram_2917, MEM_stage_inst_dmem_ram_2918, MEM_stage_inst_dmem_ram_2919, MEM_stage_inst_dmem_ram_2920, MEM_stage_inst_dmem_ram_2921, MEM_stage_inst_dmem_ram_2922, MEM_stage_inst_dmem_ram_2923, MEM_stage_inst_dmem_ram_2924, MEM_stage_inst_dmem_ram_2925, MEM_stage_inst_dmem_ram_2926, MEM_stage_inst_dmem_ram_2927, MEM_stage_inst_dmem_ram_2928, MEM_stage_inst_dmem_ram_2929, MEM_stage_inst_dmem_ram_2930, MEM_stage_inst_dmem_ram_2931, MEM_stage_inst_dmem_ram_2932, MEM_stage_inst_dmem_ram_2933, MEM_stage_inst_dmem_ram_2934, MEM_stage_inst_dmem_ram_2935, MEM_stage_inst_dmem_ram_2936, MEM_stage_inst_dmem_ram_2937, MEM_stage_inst_dmem_ram_2938, MEM_stage_inst_dmem_ram_2939, MEM_stage_inst_dmem_ram_2940, MEM_stage_inst_dmem_ram_2941, MEM_stage_inst_dmem_ram_2942, MEM_stage_inst_dmem_ram_2943, MEM_stage_inst_dmem_ram_2944, MEM_stage_inst_dmem_ram_2945, MEM_stage_inst_dmem_ram_2946, MEM_stage_inst_dmem_ram_2947, MEM_stage_inst_dmem_ram_2948, MEM_stage_inst_dmem_ram_2949, MEM_stage_inst_dmem_ram_2950, MEM_stage_inst_dmem_ram_2951, MEM_stage_inst_dmem_ram_2952, MEM_stage_inst_dmem_ram_2953, MEM_stage_inst_dmem_ram_2954, MEM_stage_inst_dmem_ram_2955, MEM_stage_inst_dmem_ram_2956, MEM_stage_inst_dmem_ram_2957, MEM_stage_inst_dmem_ram_2958, MEM_stage_inst_dmem_ram_2959, MEM_stage_inst_dmem_ram_2960, MEM_stage_inst_dmem_ram_2961, MEM_stage_inst_dmem_ram_2962, MEM_stage_inst_dmem_ram_2963, MEM_stage_inst_dmem_ram_2964, MEM_stage_inst_dmem_ram_2965, MEM_stage_inst_dmem_ram_2966, MEM_stage_inst_dmem_ram_2967, MEM_stage_inst_dmem_ram_2968, MEM_stage_inst_dmem_ram_2969, MEM_stage_inst_dmem_ram_2970, MEM_stage_inst_dmem_ram_2971, MEM_stage_inst_dmem_ram_2972, MEM_stage_inst_dmem_ram_2973, MEM_stage_inst_dmem_ram_2974, MEM_stage_inst_dmem_ram_2975, MEM_stage_inst_dmem_ram_2976, MEM_stage_inst_dmem_ram_2977, MEM_stage_inst_dmem_ram_2978, MEM_stage_inst_dmem_ram_2979, MEM_stage_inst_dmem_ram_2980, MEM_stage_inst_dmem_ram_2981, MEM_stage_inst_dmem_ram_2982, MEM_stage_inst_dmem_ram_2983, MEM_stage_inst_dmem_ram_2984, MEM_stage_inst_dmem_ram_2985, MEM_stage_inst_dmem_ram_2986, MEM_stage_inst_dmem_ram_2987, MEM_stage_inst_dmem_ram_2988, MEM_stage_inst_dmem_ram_2989, MEM_stage_inst_dmem_ram_2990, MEM_stage_inst_dmem_ram_2991, MEM_stage_inst_dmem_ram_2992, MEM_stage_inst_dmem_ram_2993, MEM_stage_inst_dmem_ram_2994, MEM_stage_inst_dmem_ram_2995, MEM_stage_inst_dmem_ram_2996, MEM_stage_inst_dmem_ram_2997, MEM_stage_inst_dmem_ram_2998, MEM_stage_inst_dmem_ram_2999, MEM_stage_inst_dmem_ram_3000, MEM_stage_inst_dmem_ram_3001, MEM_stage_inst_dmem_ram_3002, MEM_stage_inst_dmem_ram_3003, MEM_stage_inst_dmem_ram_3004, MEM_stage_inst_dmem_ram_3005, MEM_stage_inst_dmem_ram_3006, MEM_stage_inst_dmem_ram_3007, MEM_stage_inst_dmem_ram_3008, MEM_stage_inst_dmem_ram_3009, MEM_stage_inst_dmem_ram_3010, MEM_stage_inst_dmem_ram_3011, MEM_stage_inst_dmem_ram_3012, MEM_stage_inst_dmem_ram_3013, MEM_stage_inst_dmem_ram_3014, MEM_stage_inst_dmem_ram_3015, MEM_stage_inst_dmem_ram_3016, MEM_stage_inst_dmem_ram_3017, MEM_stage_inst_dmem_ram_3018, MEM_stage_inst_dmem_ram_3019, MEM_stage_inst_dmem_ram_3020, MEM_stage_inst_dmem_ram_3021, MEM_stage_inst_dmem_ram_3022, MEM_stage_inst_dmem_ram_3023, MEM_stage_inst_dmem_ram_3024, MEM_stage_inst_dmem_ram_3025, MEM_stage_inst_dmem_ram_3026, MEM_stage_inst_dmem_ram_3027, MEM_stage_inst_dmem_ram_3028, MEM_stage_inst_dmem_ram_3029, MEM_stage_inst_dmem_ram_3030, MEM_stage_inst_dmem_ram_3031, MEM_stage_inst_dmem_ram_3032, MEM_stage_inst_dmem_ram_3033, MEM_stage_inst_dmem_ram_3034, MEM_stage_inst_dmem_ram_3035, MEM_stage_inst_dmem_ram_3036, MEM_stage_inst_dmem_ram_3037, MEM_stage_inst_dmem_ram_3038, MEM_stage_inst_dmem_ram_3039, MEM_stage_inst_dmem_ram_3040, MEM_stage_inst_dmem_ram_3041, MEM_stage_inst_dmem_ram_3042, MEM_stage_inst_dmem_ram_3043, MEM_stage_inst_dmem_ram_3044, MEM_stage_inst_dmem_ram_3045, MEM_stage_inst_dmem_ram_3046, MEM_stage_inst_dmem_ram_3047, MEM_stage_inst_dmem_ram_3048, MEM_stage_inst_dmem_ram_3049, MEM_stage_inst_dmem_ram_3050, MEM_stage_inst_dmem_ram_3051, MEM_stage_inst_dmem_ram_3052, MEM_stage_inst_dmem_ram_3053, MEM_stage_inst_dmem_ram_3054, MEM_stage_inst_dmem_ram_3055, MEM_stage_inst_dmem_ram_3056, MEM_stage_inst_dmem_ram_3057, MEM_stage_inst_dmem_ram_3058, MEM_stage_inst_dmem_ram_3059, MEM_stage_inst_dmem_ram_3060, MEM_stage_inst_dmem_ram_3061, MEM_stage_inst_dmem_ram_3062, MEM_stage_inst_dmem_ram_3063, MEM_stage_inst_dmem_ram_3064, MEM_stage_inst_dmem_ram_3065, MEM_stage_inst_dmem_ram_3066, MEM_stage_inst_dmem_ram_3067, MEM_stage_inst_dmem_ram_3068, MEM_stage_inst_dmem_ram_3069, MEM_stage_inst_dmem_ram_3070, MEM_stage_inst_dmem_ram_3071, MEM_stage_inst_dmem_ram_2048, MEM_stage_inst_dmem_ram_2049, MEM_stage_inst_dmem_ram_2050, MEM_stage_inst_dmem_ram_2051, MEM_stage_inst_dmem_ram_2052, MEM_stage_inst_dmem_ram_2053, MEM_stage_inst_dmem_ram_2054, MEM_stage_inst_dmem_ram_2055, MEM_stage_inst_dmem_ram_2056, MEM_stage_inst_dmem_ram_2057, MEM_stage_inst_dmem_ram_2058, MEM_stage_inst_dmem_ram_2059, MEM_stage_inst_dmem_ram_2060, MEM_stage_inst_dmem_ram_2061, MEM_stage_inst_dmem_ram_2062, MEM_stage_inst_dmem_ram_2063, MEM_stage_inst_dmem_ram_2064, MEM_stage_inst_dmem_ram_2065, MEM_stage_inst_dmem_ram_2066, MEM_stage_inst_dmem_ram_2067, MEM_stage_inst_dmem_ram_2068, MEM_stage_inst_dmem_ram_2069, MEM_stage_inst_dmem_ram_2070, MEM_stage_inst_dmem_ram_2071, MEM_stage_inst_dmem_ram_2072, MEM_stage_inst_dmem_ram_2073, MEM_stage_inst_dmem_ram_2074, MEM_stage_inst_dmem_ram_2075, MEM_stage_inst_dmem_ram_2076, MEM_stage_inst_dmem_ram_2077, MEM_stage_inst_dmem_ram_2078, MEM_stage_inst_dmem_ram_2079, MEM_stage_inst_dmem_ram_2080, MEM_stage_inst_dmem_ram_2081, MEM_stage_inst_dmem_ram_2082, MEM_stage_inst_dmem_ram_2083, MEM_stage_inst_dmem_ram_2084, MEM_stage_inst_dmem_ram_2085, MEM_stage_inst_dmem_ram_2086, MEM_stage_inst_dmem_ram_2087, MEM_stage_inst_dmem_ram_2088, MEM_stage_inst_dmem_ram_2089, MEM_stage_inst_dmem_ram_2090, MEM_stage_inst_dmem_ram_2091, MEM_stage_inst_dmem_ram_2092, MEM_stage_inst_dmem_ram_2093, MEM_stage_inst_dmem_ram_2094, MEM_stage_inst_dmem_ram_2095, MEM_stage_inst_dmem_ram_2096, MEM_stage_inst_dmem_ram_2097, MEM_stage_inst_dmem_ram_2098, MEM_stage_inst_dmem_ram_2099, MEM_stage_inst_dmem_ram_2100, MEM_stage_inst_dmem_ram_2101, MEM_stage_inst_dmem_ram_2102, MEM_stage_inst_dmem_ram_2103, MEM_stage_inst_dmem_ram_2104, MEM_stage_inst_dmem_ram_2105, MEM_stage_inst_dmem_ram_2106, MEM_stage_inst_dmem_ram_2107, MEM_stage_inst_dmem_ram_2108, MEM_stage_inst_dmem_ram_2109, MEM_stage_inst_dmem_ram_2110, MEM_stage_inst_dmem_ram_2111, MEM_stage_inst_dmem_ram_2112, MEM_stage_inst_dmem_ram_2113, MEM_stage_inst_dmem_ram_2114, MEM_stage_inst_dmem_ram_2115, MEM_stage_inst_dmem_ram_2116, MEM_stage_inst_dmem_ram_2117, MEM_stage_inst_dmem_ram_2118, MEM_stage_inst_dmem_ram_2119, MEM_stage_inst_dmem_ram_2120, MEM_stage_inst_dmem_ram_2121, MEM_stage_inst_dmem_ram_2122, MEM_stage_inst_dmem_ram_2123, MEM_stage_inst_dmem_ram_2124, MEM_stage_inst_dmem_ram_2125, MEM_stage_inst_dmem_ram_2126, MEM_stage_inst_dmem_ram_2127, MEM_stage_inst_dmem_ram_2128, MEM_stage_inst_dmem_ram_2129, MEM_stage_inst_dmem_ram_2130, MEM_stage_inst_dmem_ram_2131, MEM_stage_inst_dmem_ram_2132, MEM_stage_inst_dmem_ram_2133, MEM_stage_inst_dmem_ram_2134, MEM_stage_inst_dmem_ram_2135, MEM_stage_inst_dmem_ram_2136, MEM_stage_inst_dmem_ram_2137, MEM_stage_inst_dmem_ram_2138, MEM_stage_inst_dmem_ram_2139, MEM_stage_inst_dmem_ram_2140, MEM_stage_inst_dmem_ram_2141, MEM_stage_inst_dmem_ram_2142, MEM_stage_inst_dmem_ram_2143, MEM_stage_inst_dmem_ram_2144, MEM_stage_inst_dmem_ram_2145, MEM_stage_inst_dmem_ram_2146, MEM_stage_inst_dmem_ram_2147, MEM_stage_inst_dmem_ram_2148, MEM_stage_inst_dmem_ram_2149, MEM_stage_inst_dmem_ram_2150, MEM_stage_inst_dmem_ram_2151, MEM_stage_inst_dmem_ram_2152, MEM_stage_inst_dmem_ram_2153, MEM_stage_inst_dmem_ram_2154, MEM_stage_inst_dmem_ram_2155, MEM_stage_inst_dmem_ram_2156, MEM_stage_inst_dmem_ram_2157, MEM_stage_inst_dmem_ram_2158, MEM_stage_inst_dmem_ram_2159, MEM_stage_inst_dmem_ram_2160, MEM_stage_inst_dmem_ram_2161, MEM_stage_inst_dmem_ram_2162, MEM_stage_inst_dmem_ram_2163, MEM_stage_inst_dmem_ram_2164, MEM_stage_inst_dmem_ram_2165, MEM_stage_inst_dmem_ram_2166, MEM_stage_inst_dmem_ram_2167, MEM_stage_inst_dmem_ram_2168, MEM_stage_inst_dmem_ram_2169, MEM_stage_inst_dmem_ram_2170, MEM_stage_inst_dmem_ram_2171, MEM_stage_inst_dmem_ram_2172, MEM_stage_inst_dmem_ram_2173, MEM_stage_inst_dmem_ram_2174, MEM_stage_inst_dmem_ram_2175, MEM_stage_inst_dmem_ram_2176, MEM_stage_inst_dmem_ram_2177, MEM_stage_inst_dmem_ram_2178, MEM_stage_inst_dmem_ram_2179, MEM_stage_inst_dmem_ram_2180, MEM_stage_inst_dmem_ram_2181, MEM_stage_inst_dmem_ram_2182, MEM_stage_inst_dmem_ram_2183, MEM_stage_inst_dmem_ram_2184, MEM_stage_inst_dmem_ram_2185, MEM_stage_inst_dmem_ram_2186, MEM_stage_inst_dmem_ram_2187, MEM_stage_inst_dmem_ram_2188, MEM_stage_inst_dmem_ram_2189, MEM_stage_inst_dmem_ram_2190, MEM_stage_inst_dmem_ram_2191, MEM_stage_inst_dmem_ram_2192, MEM_stage_inst_dmem_ram_2193, MEM_stage_inst_dmem_ram_2194, MEM_stage_inst_dmem_ram_2195, MEM_stage_inst_dmem_ram_2196, MEM_stage_inst_dmem_ram_2197, MEM_stage_inst_dmem_ram_2198, MEM_stage_inst_dmem_ram_2199, MEM_stage_inst_dmem_ram_2200, MEM_stage_inst_dmem_ram_2201, MEM_stage_inst_dmem_ram_2202, MEM_stage_inst_dmem_ram_2203, MEM_stage_inst_dmem_ram_2204, MEM_stage_inst_dmem_ram_2205, MEM_stage_inst_dmem_ram_2206, MEM_stage_inst_dmem_ram_2207, MEM_stage_inst_dmem_ram_2208, MEM_stage_inst_dmem_ram_2209, MEM_stage_inst_dmem_ram_2210, MEM_stage_inst_dmem_ram_2211, MEM_stage_inst_dmem_ram_2212, MEM_stage_inst_dmem_ram_2213, MEM_stage_inst_dmem_ram_2214, MEM_stage_inst_dmem_ram_2215, MEM_stage_inst_dmem_ram_2216, MEM_stage_inst_dmem_ram_2217, MEM_stage_inst_dmem_ram_2218, MEM_stage_inst_dmem_ram_2219, MEM_stage_inst_dmem_ram_2220, MEM_stage_inst_dmem_ram_2221, MEM_stage_inst_dmem_ram_2222, MEM_stage_inst_dmem_ram_2223, MEM_stage_inst_dmem_ram_2224, MEM_stage_inst_dmem_ram_2225, MEM_stage_inst_dmem_ram_2226, MEM_stage_inst_dmem_ram_2227, MEM_stage_inst_dmem_ram_2228, MEM_stage_inst_dmem_ram_2229, MEM_stage_inst_dmem_ram_2230, MEM_stage_inst_dmem_ram_2231, MEM_stage_inst_dmem_ram_2232, MEM_stage_inst_dmem_ram_2233, MEM_stage_inst_dmem_ram_2234, MEM_stage_inst_dmem_ram_2235, MEM_stage_inst_dmem_ram_2236, MEM_stage_inst_dmem_ram_2237, MEM_stage_inst_dmem_ram_2238, MEM_stage_inst_dmem_ram_2239, MEM_stage_inst_dmem_ram_2240, MEM_stage_inst_dmem_ram_2241, MEM_stage_inst_dmem_ram_2242, MEM_stage_inst_dmem_ram_2243, MEM_stage_inst_dmem_ram_2244, MEM_stage_inst_dmem_ram_2245, MEM_stage_inst_dmem_ram_2246, MEM_stage_inst_dmem_ram_2247, MEM_stage_inst_dmem_ram_2248, MEM_stage_inst_dmem_ram_2249, MEM_stage_inst_dmem_ram_2250, MEM_stage_inst_dmem_ram_2251, MEM_stage_inst_dmem_ram_2252, MEM_stage_inst_dmem_ram_2253, MEM_stage_inst_dmem_ram_2254, MEM_stage_inst_dmem_ram_2255, MEM_stage_inst_dmem_ram_2256, MEM_stage_inst_dmem_ram_2257, MEM_stage_inst_dmem_ram_2258, MEM_stage_inst_dmem_ram_2259, MEM_stage_inst_dmem_ram_2260, MEM_stage_inst_dmem_ram_2261, MEM_stage_inst_dmem_ram_2262, MEM_stage_inst_dmem_ram_2263, MEM_stage_inst_dmem_ram_2264, MEM_stage_inst_dmem_ram_2265, MEM_stage_inst_dmem_ram_2266, MEM_stage_inst_dmem_ram_2267, MEM_stage_inst_dmem_ram_2268, MEM_stage_inst_dmem_ram_2269, MEM_stage_inst_dmem_ram_2270, MEM_stage_inst_dmem_ram_2271, MEM_stage_inst_dmem_ram_2272, MEM_stage_inst_dmem_ram_2273, MEM_stage_inst_dmem_ram_2274, MEM_stage_inst_dmem_ram_2275, MEM_stage_inst_dmem_ram_2276, MEM_stage_inst_dmem_ram_2277, MEM_stage_inst_dmem_ram_2278, MEM_stage_inst_dmem_ram_2279, MEM_stage_inst_dmem_ram_2280, MEM_stage_inst_dmem_ram_2281, MEM_stage_inst_dmem_ram_2282, MEM_stage_inst_dmem_ram_2283, MEM_stage_inst_dmem_ram_2284, MEM_stage_inst_dmem_ram_2285, MEM_stage_inst_dmem_ram_2286, MEM_stage_inst_dmem_ram_2287, MEM_stage_inst_dmem_ram_2288, MEM_stage_inst_dmem_ram_2289, MEM_stage_inst_dmem_ram_2290, MEM_stage_inst_dmem_ram_2291, MEM_stage_inst_dmem_ram_2292, MEM_stage_inst_dmem_ram_2293, MEM_stage_inst_dmem_ram_2294, MEM_stage_inst_dmem_ram_2295, MEM_stage_inst_dmem_ram_2296, MEM_stage_inst_dmem_ram_2297, MEM_stage_inst_dmem_ram_2298, MEM_stage_inst_dmem_ram_2299, MEM_stage_inst_dmem_ram_2300, MEM_stage_inst_dmem_ram_2301, MEM_stage_inst_dmem_ram_2302, MEM_stage_inst_dmem_ram_2303, MEM_stage_inst_dmem_ram_2304, MEM_stage_inst_dmem_ram_2305, MEM_stage_inst_dmem_ram_2306, MEM_stage_inst_dmem_ram_2307, MEM_stage_inst_dmem_ram_2308, MEM_stage_inst_dmem_ram_2309, MEM_stage_inst_dmem_ram_2310, MEM_stage_inst_dmem_ram_2311, MEM_stage_inst_dmem_ram_2312, MEM_stage_inst_dmem_ram_2313, MEM_stage_inst_dmem_ram_2314, MEM_stage_inst_dmem_ram_2315, MEM_stage_inst_dmem_ram_2316, MEM_stage_inst_dmem_ram_2317, MEM_stage_inst_dmem_ram_2318, MEM_stage_inst_dmem_ram_2319, MEM_stage_inst_dmem_ram_2320, MEM_stage_inst_dmem_ram_2321, MEM_stage_inst_dmem_ram_2322, MEM_stage_inst_dmem_ram_2323, MEM_stage_inst_dmem_ram_2324, MEM_stage_inst_dmem_ram_2325, MEM_stage_inst_dmem_ram_2326, MEM_stage_inst_dmem_ram_2327, MEM_stage_inst_dmem_ram_2328, MEM_stage_inst_dmem_ram_2329, MEM_stage_inst_dmem_ram_2330, MEM_stage_inst_dmem_ram_2331, MEM_stage_inst_dmem_ram_2332, MEM_stage_inst_dmem_ram_2333, MEM_stage_inst_dmem_ram_2334, MEM_stage_inst_dmem_ram_2335, MEM_stage_inst_dmem_ram_2336, MEM_stage_inst_dmem_ram_2337, MEM_stage_inst_dmem_ram_2338, MEM_stage_inst_dmem_ram_2339, MEM_stage_inst_dmem_ram_2340, MEM_stage_inst_dmem_ram_2341, MEM_stage_inst_dmem_ram_2342, MEM_stage_inst_dmem_ram_2343, MEM_stage_inst_dmem_ram_2344, MEM_stage_inst_dmem_ram_2345, MEM_stage_inst_dmem_ram_2346, MEM_stage_inst_dmem_ram_2347, MEM_stage_inst_dmem_ram_2348, MEM_stage_inst_dmem_ram_2349, MEM_stage_inst_dmem_ram_2350, MEM_stage_inst_dmem_ram_2351, MEM_stage_inst_dmem_ram_2352, MEM_stage_inst_dmem_ram_2353, MEM_stage_inst_dmem_ram_2354, MEM_stage_inst_dmem_ram_2355, MEM_stage_inst_dmem_ram_2356, MEM_stage_inst_dmem_ram_2357, MEM_stage_inst_dmem_ram_2358, MEM_stage_inst_dmem_ram_2359, MEM_stage_inst_dmem_ram_2360, MEM_stage_inst_dmem_ram_2361, MEM_stage_inst_dmem_ram_2362, MEM_stage_inst_dmem_ram_2363, MEM_stage_inst_dmem_ram_2364, MEM_stage_inst_dmem_ram_2365, MEM_stage_inst_dmem_ram_2366, MEM_stage_inst_dmem_ram_2367, MEM_stage_inst_dmem_ram_2368, MEM_stage_inst_dmem_ram_2369, MEM_stage_inst_dmem_ram_2370, MEM_stage_inst_dmem_ram_2371, MEM_stage_inst_dmem_ram_2372, MEM_stage_inst_dmem_ram_2373, MEM_stage_inst_dmem_ram_2374, MEM_stage_inst_dmem_ram_2375, MEM_stage_inst_dmem_ram_2376, MEM_stage_inst_dmem_ram_2377, MEM_stage_inst_dmem_ram_2378, MEM_stage_inst_dmem_ram_2379, MEM_stage_inst_dmem_ram_2380, MEM_stage_inst_dmem_ram_2381, MEM_stage_inst_dmem_ram_2382, MEM_stage_inst_dmem_ram_2383, MEM_stage_inst_dmem_ram_2384, MEM_stage_inst_dmem_ram_2385, MEM_stage_inst_dmem_ram_2386, MEM_stage_inst_dmem_ram_2387, MEM_stage_inst_dmem_ram_2388, MEM_stage_inst_dmem_ram_2389, MEM_stage_inst_dmem_ram_2390, MEM_stage_inst_dmem_ram_2391, MEM_stage_inst_dmem_ram_2392, MEM_stage_inst_dmem_ram_2393, MEM_stage_inst_dmem_ram_2394, MEM_stage_inst_dmem_ram_2395, MEM_stage_inst_dmem_ram_2396, MEM_stage_inst_dmem_ram_2397, MEM_stage_inst_dmem_ram_2398, MEM_stage_inst_dmem_ram_2399, MEM_stage_inst_dmem_ram_2400, MEM_stage_inst_dmem_ram_2401, MEM_stage_inst_dmem_ram_2402, MEM_stage_inst_dmem_ram_2403, MEM_stage_inst_dmem_ram_2404, MEM_stage_inst_dmem_ram_2405, MEM_stage_inst_dmem_ram_2406, MEM_stage_inst_dmem_ram_2407, MEM_stage_inst_dmem_ram_2408, MEM_stage_inst_dmem_ram_2409, MEM_stage_inst_dmem_ram_2410, MEM_stage_inst_dmem_ram_2411, MEM_stage_inst_dmem_ram_2412, MEM_stage_inst_dmem_ram_2413, MEM_stage_inst_dmem_ram_2414, MEM_stage_inst_dmem_ram_2415, MEM_stage_inst_dmem_ram_2416, MEM_stage_inst_dmem_ram_2417, MEM_stage_inst_dmem_ram_2418, MEM_stage_inst_dmem_ram_2419, MEM_stage_inst_dmem_ram_2420, MEM_stage_inst_dmem_ram_2421, MEM_stage_inst_dmem_ram_2422, MEM_stage_inst_dmem_ram_2423, MEM_stage_inst_dmem_ram_2424, MEM_stage_inst_dmem_ram_2425, MEM_stage_inst_dmem_ram_2426, MEM_stage_inst_dmem_ram_2427, MEM_stage_inst_dmem_ram_2428, MEM_stage_inst_dmem_ram_2429, MEM_stage_inst_dmem_ram_2430, MEM_stage_inst_dmem_ram_2431, MEM_stage_inst_dmem_ram_2432, MEM_stage_inst_dmem_ram_2433, MEM_stage_inst_dmem_ram_2434, MEM_stage_inst_dmem_ram_2435, MEM_stage_inst_dmem_ram_2436, MEM_stage_inst_dmem_ram_2437, MEM_stage_inst_dmem_ram_2438, MEM_stage_inst_dmem_ram_2439, MEM_stage_inst_dmem_ram_2440, MEM_stage_inst_dmem_ram_2441, MEM_stage_inst_dmem_ram_2442, MEM_stage_inst_dmem_ram_2443, MEM_stage_inst_dmem_ram_2444, MEM_stage_inst_dmem_ram_2445, MEM_stage_inst_dmem_ram_2446, MEM_stage_inst_dmem_ram_2447, MEM_stage_inst_dmem_ram_2448, MEM_stage_inst_dmem_ram_2449, MEM_stage_inst_dmem_ram_2450, MEM_stage_inst_dmem_ram_2451, MEM_stage_inst_dmem_ram_2452, MEM_stage_inst_dmem_ram_2453, MEM_stage_inst_dmem_ram_2454, MEM_stage_inst_dmem_ram_2455, MEM_stage_inst_dmem_ram_2456, MEM_stage_inst_dmem_ram_2457, MEM_stage_inst_dmem_ram_2458, MEM_stage_inst_dmem_ram_2459, MEM_stage_inst_dmem_ram_2460, MEM_stage_inst_dmem_ram_2461, MEM_stage_inst_dmem_ram_2462, MEM_stage_inst_dmem_ram_2463, MEM_stage_inst_dmem_ram_2464, MEM_stage_inst_dmem_ram_2465, MEM_stage_inst_dmem_ram_2466, MEM_stage_inst_dmem_ram_2467, MEM_stage_inst_dmem_ram_2468, MEM_stage_inst_dmem_ram_2469, MEM_stage_inst_dmem_ram_2470, MEM_stage_inst_dmem_ram_2471, MEM_stage_inst_dmem_ram_2472, MEM_stage_inst_dmem_ram_2473, MEM_stage_inst_dmem_ram_2474, MEM_stage_inst_dmem_ram_2475, MEM_stage_inst_dmem_ram_2476, MEM_stage_inst_dmem_ram_2477, MEM_stage_inst_dmem_ram_2478, MEM_stage_inst_dmem_ram_2479, MEM_stage_inst_dmem_ram_2480, MEM_stage_inst_dmem_ram_2481, MEM_stage_inst_dmem_ram_2482, MEM_stage_inst_dmem_ram_2483, MEM_stage_inst_dmem_ram_2484, MEM_stage_inst_dmem_ram_2485, MEM_stage_inst_dmem_ram_2486, MEM_stage_inst_dmem_ram_2487, MEM_stage_inst_dmem_ram_2488, MEM_stage_inst_dmem_ram_2489, MEM_stage_inst_dmem_ram_2490, MEM_stage_inst_dmem_ram_2491, MEM_stage_inst_dmem_ram_2492, MEM_stage_inst_dmem_ram_2493, MEM_stage_inst_dmem_ram_2494, MEM_stage_inst_dmem_ram_2495, MEM_stage_inst_dmem_ram_2496, MEM_stage_inst_dmem_ram_2497, MEM_stage_inst_dmem_ram_2498, MEM_stage_inst_dmem_ram_2499, MEM_stage_inst_dmem_ram_2500, MEM_stage_inst_dmem_ram_2501, MEM_stage_inst_dmem_ram_2502, MEM_stage_inst_dmem_ram_2503, MEM_stage_inst_dmem_ram_2504, MEM_stage_inst_dmem_ram_2505, MEM_stage_inst_dmem_ram_2506, MEM_stage_inst_dmem_ram_2507, MEM_stage_inst_dmem_ram_2508, MEM_stage_inst_dmem_ram_2509, MEM_stage_inst_dmem_ram_2510, MEM_stage_inst_dmem_ram_2511, MEM_stage_inst_dmem_ram_2512, MEM_stage_inst_dmem_ram_2513, MEM_stage_inst_dmem_ram_2514, MEM_stage_inst_dmem_ram_2515, MEM_stage_inst_dmem_ram_2516, MEM_stage_inst_dmem_ram_2517, MEM_stage_inst_dmem_ram_2518, MEM_stage_inst_dmem_ram_2519, MEM_stage_inst_dmem_ram_2520, MEM_stage_inst_dmem_ram_2521, MEM_stage_inst_dmem_ram_2522, MEM_stage_inst_dmem_ram_2523, MEM_stage_inst_dmem_ram_2524, MEM_stage_inst_dmem_ram_2525, MEM_stage_inst_dmem_ram_2526, MEM_stage_inst_dmem_ram_2527, MEM_stage_inst_dmem_ram_2528, MEM_stage_inst_dmem_ram_2529, MEM_stage_inst_dmem_ram_2530, MEM_stage_inst_dmem_ram_2531, MEM_stage_inst_dmem_ram_2532, MEM_stage_inst_dmem_ram_2533, MEM_stage_inst_dmem_ram_2534, MEM_stage_inst_dmem_ram_2535, MEM_stage_inst_dmem_ram_2536, MEM_stage_inst_dmem_ram_2537, MEM_stage_inst_dmem_ram_2538, MEM_stage_inst_dmem_ram_2539, MEM_stage_inst_dmem_ram_2540, MEM_stage_inst_dmem_ram_2541, MEM_stage_inst_dmem_ram_2542, MEM_stage_inst_dmem_ram_2543, MEM_stage_inst_dmem_ram_2544, MEM_stage_inst_dmem_ram_2545, MEM_stage_inst_dmem_ram_2546, MEM_stage_inst_dmem_ram_2547, MEM_stage_inst_dmem_ram_2548, MEM_stage_inst_dmem_ram_2549, MEM_stage_inst_dmem_ram_2550, MEM_stage_inst_dmem_ram_2551, MEM_stage_inst_dmem_ram_2552, MEM_stage_inst_dmem_ram_2553, MEM_stage_inst_dmem_ram_2554, MEM_stage_inst_dmem_ram_2555, MEM_stage_inst_dmem_ram_2556, MEM_stage_inst_dmem_ram_2557, MEM_stage_inst_dmem_ram_2558, MEM_stage_inst_dmem_ram_2559, MEM_stage_inst_dmem_ram_1536, MEM_stage_inst_dmem_ram_1537, MEM_stage_inst_dmem_ram_1538, MEM_stage_inst_dmem_ram_1539, MEM_stage_inst_dmem_ram_1540, MEM_stage_inst_dmem_ram_1541, MEM_stage_inst_dmem_ram_1542, MEM_stage_inst_dmem_ram_1543, MEM_stage_inst_dmem_ram_1544, MEM_stage_inst_dmem_ram_1545, MEM_stage_inst_dmem_ram_1546, MEM_stage_inst_dmem_ram_1547, MEM_stage_inst_dmem_ram_1548, MEM_stage_inst_dmem_ram_1549, MEM_stage_inst_dmem_ram_1550, MEM_stage_inst_dmem_ram_1551, MEM_stage_inst_dmem_ram_1552, MEM_stage_inst_dmem_ram_1553, MEM_stage_inst_dmem_ram_1554, MEM_stage_inst_dmem_ram_1555, MEM_stage_inst_dmem_ram_1556, MEM_stage_inst_dmem_ram_1557, MEM_stage_inst_dmem_ram_1558, MEM_stage_inst_dmem_ram_1559, MEM_stage_inst_dmem_ram_1560, MEM_stage_inst_dmem_ram_1561, MEM_stage_inst_dmem_ram_1562, MEM_stage_inst_dmem_ram_1563, MEM_stage_inst_dmem_ram_1564, MEM_stage_inst_dmem_ram_1565, MEM_stage_inst_dmem_ram_1566, MEM_stage_inst_dmem_ram_1567, MEM_stage_inst_dmem_ram_1568, MEM_stage_inst_dmem_ram_1569, MEM_stage_inst_dmem_ram_1570, MEM_stage_inst_dmem_ram_1571, MEM_stage_inst_dmem_ram_1572, MEM_stage_inst_dmem_ram_1573, MEM_stage_inst_dmem_ram_1574, MEM_stage_inst_dmem_ram_1575, MEM_stage_inst_dmem_ram_1576, MEM_stage_inst_dmem_ram_1577, MEM_stage_inst_dmem_ram_1578, MEM_stage_inst_dmem_ram_1579, MEM_stage_inst_dmem_ram_1580, MEM_stage_inst_dmem_ram_1581, MEM_stage_inst_dmem_ram_1582, MEM_stage_inst_dmem_ram_1583, MEM_stage_inst_dmem_ram_1584, MEM_stage_inst_dmem_ram_1585, MEM_stage_inst_dmem_ram_1586, MEM_stage_inst_dmem_ram_1587, MEM_stage_inst_dmem_ram_1588, MEM_stage_inst_dmem_ram_1589, MEM_stage_inst_dmem_ram_1590, MEM_stage_inst_dmem_ram_1591, MEM_stage_inst_dmem_ram_1592, MEM_stage_inst_dmem_ram_1593, MEM_stage_inst_dmem_ram_1594, MEM_stage_inst_dmem_ram_1595, MEM_stage_inst_dmem_ram_1596, MEM_stage_inst_dmem_ram_1597, MEM_stage_inst_dmem_ram_1598, MEM_stage_inst_dmem_ram_1599, MEM_stage_inst_dmem_ram_1600, MEM_stage_inst_dmem_ram_1601, MEM_stage_inst_dmem_ram_1602, MEM_stage_inst_dmem_ram_1603, MEM_stage_inst_dmem_ram_1604, MEM_stage_inst_dmem_ram_1605, MEM_stage_inst_dmem_ram_1606, MEM_stage_inst_dmem_ram_1607, MEM_stage_inst_dmem_ram_1608, MEM_stage_inst_dmem_ram_1609, MEM_stage_inst_dmem_ram_1610, MEM_stage_inst_dmem_ram_1611, MEM_stage_inst_dmem_ram_1612, MEM_stage_inst_dmem_ram_1613, MEM_stage_inst_dmem_ram_1614, MEM_stage_inst_dmem_ram_1615, MEM_stage_inst_dmem_ram_1616, MEM_stage_inst_dmem_ram_1617, MEM_stage_inst_dmem_ram_1618, MEM_stage_inst_dmem_ram_1619, MEM_stage_inst_dmem_ram_1620, MEM_stage_inst_dmem_ram_1621, MEM_stage_inst_dmem_ram_1622, MEM_stage_inst_dmem_ram_1623, MEM_stage_inst_dmem_ram_1624, MEM_stage_inst_dmem_ram_1625, MEM_stage_inst_dmem_ram_1626, MEM_stage_inst_dmem_ram_1627, MEM_stage_inst_dmem_ram_1628, MEM_stage_inst_dmem_ram_1629, MEM_stage_inst_dmem_ram_1630, MEM_stage_inst_dmem_ram_1631, MEM_stage_inst_dmem_ram_1632, MEM_stage_inst_dmem_ram_1633, MEM_stage_inst_dmem_ram_1634, MEM_stage_inst_dmem_ram_1635, MEM_stage_inst_dmem_ram_1636, MEM_stage_inst_dmem_ram_1637, MEM_stage_inst_dmem_ram_1638, MEM_stage_inst_dmem_ram_1639, MEM_stage_inst_dmem_ram_1640, MEM_stage_inst_dmem_ram_1641, MEM_stage_inst_dmem_ram_1642, MEM_stage_inst_dmem_ram_1643, MEM_stage_inst_dmem_ram_1644, MEM_stage_inst_dmem_ram_1645, MEM_stage_inst_dmem_ram_1646, MEM_stage_inst_dmem_ram_1647, MEM_stage_inst_dmem_ram_1648, MEM_stage_inst_dmem_ram_1649, MEM_stage_inst_dmem_ram_1650, MEM_stage_inst_dmem_ram_1651, MEM_stage_inst_dmem_ram_1652, MEM_stage_inst_dmem_ram_1653, MEM_stage_inst_dmem_ram_1654, MEM_stage_inst_dmem_ram_1655, MEM_stage_inst_dmem_ram_1656, MEM_stage_inst_dmem_ram_1657, MEM_stage_inst_dmem_ram_1658, MEM_stage_inst_dmem_ram_1659, MEM_stage_inst_dmem_ram_1660, MEM_stage_inst_dmem_ram_1661, MEM_stage_inst_dmem_ram_1662, MEM_stage_inst_dmem_ram_1663, MEM_stage_inst_dmem_ram_1664, MEM_stage_inst_dmem_ram_1665, MEM_stage_inst_dmem_ram_1666, MEM_stage_inst_dmem_ram_1667, MEM_stage_inst_dmem_ram_1668, MEM_stage_inst_dmem_ram_1669, MEM_stage_inst_dmem_ram_1670, MEM_stage_inst_dmem_ram_1671, MEM_stage_inst_dmem_ram_1672, MEM_stage_inst_dmem_ram_1673, MEM_stage_inst_dmem_ram_1674, MEM_stage_inst_dmem_ram_1675, MEM_stage_inst_dmem_ram_1676, MEM_stage_inst_dmem_ram_1677, MEM_stage_inst_dmem_ram_1678, MEM_stage_inst_dmem_ram_1679, MEM_stage_inst_dmem_ram_1680, MEM_stage_inst_dmem_ram_1681, MEM_stage_inst_dmem_ram_1682, MEM_stage_inst_dmem_ram_1683, MEM_stage_inst_dmem_ram_1684, MEM_stage_inst_dmem_ram_1685, MEM_stage_inst_dmem_ram_1686, MEM_stage_inst_dmem_ram_1687, MEM_stage_inst_dmem_ram_1688, MEM_stage_inst_dmem_ram_1689, MEM_stage_inst_dmem_ram_1690, MEM_stage_inst_dmem_ram_1691, MEM_stage_inst_dmem_ram_1692, MEM_stage_inst_dmem_ram_1693, MEM_stage_inst_dmem_ram_1694, MEM_stage_inst_dmem_ram_1695, MEM_stage_inst_dmem_ram_1696, MEM_stage_inst_dmem_ram_1697, MEM_stage_inst_dmem_ram_1698, MEM_stage_inst_dmem_ram_1699, MEM_stage_inst_dmem_ram_1700, MEM_stage_inst_dmem_ram_1701, MEM_stage_inst_dmem_ram_1702, MEM_stage_inst_dmem_ram_1703, MEM_stage_inst_dmem_ram_1704, MEM_stage_inst_dmem_ram_1705, MEM_stage_inst_dmem_ram_1706, MEM_stage_inst_dmem_ram_1707, MEM_stage_inst_dmem_ram_1708, MEM_stage_inst_dmem_ram_1709, MEM_stage_inst_dmem_ram_1710, MEM_stage_inst_dmem_ram_1711, MEM_stage_inst_dmem_ram_1712, MEM_stage_inst_dmem_ram_1713, MEM_stage_inst_dmem_ram_1714, MEM_stage_inst_dmem_ram_1715, MEM_stage_inst_dmem_ram_1716, MEM_stage_inst_dmem_ram_1717, MEM_stage_inst_dmem_ram_1718, MEM_stage_inst_dmem_ram_1719, MEM_stage_inst_dmem_ram_1720, MEM_stage_inst_dmem_ram_1721, MEM_stage_inst_dmem_ram_1722, MEM_stage_inst_dmem_ram_1723, MEM_stage_inst_dmem_ram_1724, MEM_stage_inst_dmem_ram_1725, MEM_stage_inst_dmem_ram_1726, MEM_stage_inst_dmem_ram_1727, MEM_stage_inst_dmem_ram_1728, MEM_stage_inst_dmem_ram_1729, MEM_stage_inst_dmem_ram_1730, MEM_stage_inst_dmem_ram_1731, MEM_stage_inst_dmem_ram_1732, MEM_stage_inst_dmem_ram_1733, MEM_stage_inst_dmem_ram_1734, MEM_stage_inst_dmem_ram_1735, MEM_stage_inst_dmem_ram_1736, MEM_stage_inst_dmem_ram_1737, MEM_stage_inst_dmem_ram_1738, MEM_stage_inst_dmem_ram_1739, MEM_stage_inst_dmem_ram_1740, MEM_stage_inst_dmem_ram_1741, MEM_stage_inst_dmem_ram_1742, MEM_stage_inst_dmem_ram_1743, MEM_stage_inst_dmem_ram_1744, MEM_stage_inst_dmem_ram_1745, MEM_stage_inst_dmem_ram_1746, MEM_stage_inst_dmem_ram_1747, MEM_stage_inst_dmem_ram_1748, MEM_stage_inst_dmem_ram_1749, MEM_stage_inst_dmem_ram_1750, MEM_stage_inst_dmem_ram_1751, MEM_stage_inst_dmem_ram_1752, MEM_stage_inst_dmem_ram_1753, MEM_stage_inst_dmem_ram_1754, MEM_stage_inst_dmem_ram_1755, MEM_stage_inst_dmem_ram_1756, MEM_stage_inst_dmem_ram_1757, MEM_stage_inst_dmem_ram_1758, MEM_stage_inst_dmem_ram_1759, MEM_stage_inst_dmem_ram_1760, MEM_stage_inst_dmem_ram_1761, MEM_stage_inst_dmem_ram_1762, MEM_stage_inst_dmem_ram_1763, MEM_stage_inst_dmem_ram_1764, MEM_stage_inst_dmem_ram_1765, MEM_stage_inst_dmem_ram_1766, MEM_stage_inst_dmem_ram_1767, MEM_stage_inst_dmem_ram_1768, MEM_stage_inst_dmem_ram_1769, MEM_stage_inst_dmem_ram_1770, MEM_stage_inst_dmem_ram_1771, MEM_stage_inst_dmem_ram_1772, MEM_stage_inst_dmem_ram_1773, MEM_stage_inst_dmem_ram_1774, MEM_stage_inst_dmem_ram_1775, MEM_stage_inst_dmem_ram_1776, MEM_stage_inst_dmem_ram_1777, MEM_stage_inst_dmem_ram_1778, MEM_stage_inst_dmem_ram_1779, MEM_stage_inst_dmem_ram_1780, MEM_stage_inst_dmem_ram_1781, MEM_stage_inst_dmem_ram_1782, MEM_stage_inst_dmem_ram_1783, MEM_stage_inst_dmem_ram_1784, MEM_stage_inst_dmem_ram_1785, MEM_stage_inst_dmem_ram_1786, MEM_stage_inst_dmem_ram_1787, MEM_stage_inst_dmem_ram_1788, MEM_stage_inst_dmem_ram_1789, MEM_stage_inst_dmem_ram_1790, MEM_stage_inst_dmem_ram_1791, MEM_stage_inst_dmem_ram_1792, MEM_stage_inst_dmem_ram_1793, MEM_stage_inst_dmem_ram_1794, MEM_stage_inst_dmem_ram_1795, MEM_stage_inst_dmem_ram_1796, MEM_stage_inst_dmem_ram_1797, MEM_stage_inst_dmem_ram_1798, MEM_stage_inst_dmem_ram_1799, MEM_stage_inst_dmem_ram_1800, MEM_stage_inst_dmem_ram_1801, MEM_stage_inst_dmem_ram_1802, MEM_stage_inst_dmem_ram_1803, MEM_stage_inst_dmem_ram_1804, MEM_stage_inst_dmem_ram_1805, MEM_stage_inst_dmem_ram_1806, MEM_stage_inst_dmem_ram_1807, MEM_stage_inst_dmem_ram_1808, MEM_stage_inst_dmem_ram_1809, MEM_stage_inst_dmem_ram_1810, MEM_stage_inst_dmem_ram_1811, MEM_stage_inst_dmem_ram_1812, MEM_stage_inst_dmem_ram_1813, MEM_stage_inst_dmem_ram_1814, MEM_stage_inst_dmem_ram_1815, MEM_stage_inst_dmem_ram_1816, MEM_stage_inst_dmem_ram_1817, MEM_stage_inst_dmem_ram_1818, MEM_stage_inst_dmem_ram_1819, MEM_stage_inst_dmem_ram_1820, MEM_stage_inst_dmem_ram_1821, MEM_stage_inst_dmem_ram_1822, MEM_stage_inst_dmem_ram_1823, MEM_stage_inst_dmem_ram_1824, MEM_stage_inst_dmem_ram_1825, MEM_stage_inst_dmem_ram_1826, MEM_stage_inst_dmem_ram_1827, MEM_stage_inst_dmem_ram_1828, MEM_stage_inst_dmem_ram_1829, MEM_stage_inst_dmem_ram_1830, MEM_stage_inst_dmem_ram_1831, MEM_stage_inst_dmem_ram_1832, MEM_stage_inst_dmem_ram_1833, MEM_stage_inst_dmem_ram_1834, MEM_stage_inst_dmem_ram_1835, MEM_stage_inst_dmem_ram_1836, MEM_stage_inst_dmem_ram_1837, MEM_stage_inst_dmem_ram_1838, MEM_stage_inst_dmem_ram_1839, MEM_stage_inst_dmem_ram_1840, MEM_stage_inst_dmem_ram_1841, MEM_stage_inst_dmem_ram_1842, MEM_stage_inst_dmem_ram_1843, MEM_stage_inst_dmem_ram_1844, MEM_stage_inst_dmem_ram_1845, MEM_stage_inst_dmem_ram_1846, MEM_stage_inst_dmem_ram_1847, MEM_stage_inst_dmem_ram_1848, MEM_stage_inst_dmem_ram_1849, MEM_stage_inst_dmem_ram_1850, MEM_stage_inst_dmem_ram_1851, MEM_stage_inst_dmem_ram_1852, MEM_stage_inst_dmem_ram_1853, MEM_stage_inst_dmem_ram_1854, MEM_stage_inst_dmem_ram_1855, MEM_stage_inst_dmem_ram_1856, MEM_stage_inst_dmem_ram_1857, MEM_stage_inst_dmem_ram_1858, MEM_stage_inst_dmem_ram_1859, MEM_stage_inst_dmem_ram_1860, MEM_stage_inst_dmem_ram_1861, MEM_stage_inst_dmem_ram_1862, MEM_stage_inst_dmem_ram_1863, MEM_stage_inst_dmem_ram_1864, MEM_stage_inst_dmem_ram_1865, MEM_stage_inst_dmem_ram_1866, MEM_stage_inst_dmem_ram_1867, MEM_stage_inst_dmem_ram_1868, MEM_stage_inst_dmem_ram_1869, MEM_stage_inst_dmem_ram_1870, MEM_stage_inst_dmem_ram_1871, MEM_stage_inst_dmem_ram_1872, MEM_stage_inst_dmem_ram_1873, MEM_stage_inst_dmem_ram_1874, MEM_stage_inst_dmem_ram_1875, MEM_stage_inst_dmem_ram_1876, MEM_stage_inst_dmem_ram_1877, MEM_stage_inst_dmem_ram_1878, MEM_stage_inst_dmem_ram_1879, MEM_stage_inst_dmem_ram_1880, MEM_stage_inst_dmem_ram_1881, MEM_stage_inst_dmem_ram_1882, MEM_stage_inst_dmem_ram_1883, MEM_stage_inst_dmem_ram_1884, MEM_stage_inst_dmem_ram_1885, MEM_stage_inst_dmem_ram_1886, MEM_stage_inst_dmem_ram_1887, MEM_stage_inst_dmem_ram_1888, MEM_stage_inst_dmem_ram_1889, MEM_stage_inst_dmem_ram_1890, MEM_stage_inst_dmem_ram_1891, MEM_stage_inst_dmem_ram_1892, MEM_stage_inst_dmem_ram_1893, MEM_stage_inst_dmem_ram_1894, MEM_stage_inst_dmem_ram_1895, MEM_stage_inst_dmem_ram_1896, MEM_stage_inst_dmem_ram_1897, MEM_stage_inst_dmem_ram_1898, MEM_stage_inst_dmem_ram_1899, MEM_stage_inst_dmem_ram_1900, MEM_stage_inst_dmem_ram_1901, MEM_stage_inst_dmem_ram_1902, MEM_stage_inst_dmem_ram_1903, MEM_stage_inst_dmem_ram_1904, MEM_stage_inst_dmem_ram_1905, MEM_stage_inst_dmem_ram_1906, MEM_stage_inst_dmem_ram_1907, MEM_stage_inst_dmem_ram_1908, MEM_stage_inst_dmem_ram_1909, MEM_stage_inst_dmem_ram_1910, MEM_stage_inst_dmem_ram_1911, MEM_stage_inst_dmem_ram_1912, MEM_stage_inst_dmem_ram_1913, MEM_stage_inst_dmem_ram_1914, MEM_stage_inst_dmem_ram_1915, MEM_stage_inst_dmem_ram_1916, MEM_stage_inst_dmem_ram_1917, MEM_stage_inst_dmem_ram_1918, MEM_stage_inst_dmem_ram_1919, MEM_stage_inst_dmem_ram_1920, MEM_stage_inst_dmem_ram_1921, MEM_stage_inst_dmem_ram_1922, MEM_stage_inst_dmem_ram_1923, MEM_stage_inst_dmem_ram_1924, MEM_stage_inst_dmem_ram_1925, MEM_stage_inst_dmem_ram_1926, MEM_stage_inst_dmem_ram_1927, MEM_stage_inst_dmem_ram_1928, MEM_stage_inst_dmem_ram_1929, MEM_stage_inst_dmem_ram_1930, MEM_stage_inst_dmem_ram_1931, MEM_stage_inst_dmem_ram_1932, MEM_stage_inst_dmem_ram_1933, MEM_stage_inst_dmem_ram_1934, MEM_stage_inst_dmem_ram_1935, MEM_stage_inst_dmem_ram_1936, MEM_stage_inst_dmem_ram_1937, MEM_stage_inst_dmem_ram_1938, MEM_stage_inst_dmem_ram_1939, MEM_stage_inst_dmem_ram_1940, MEM_stage_inst_dmem_ram_1941, MEM_stage_inst_dmem_ram_1942, MEM_stage_inst_dmem_ram_1943, MEM_stage_inst_dmem_ram_1944, MEM_stage_inst_dmem_ram_1945, MEM_stage_inst_dmem_ram_1946, MEM_stage_inst_dmem_ram_1947, MEM_stage_inst_dmem_ram_1948, MEM_stage_inst_dmem_ram_1949, MEM_stage_inst_dmem_ram_1950, MEM_stage_inst_dmem_ram_1951, MEM_stage_inst_dmem_ram_1952, MEM_stage_inst_dmem_ram_1953, MEM_stage_inst_dmem_ram_1954, MEM_stage_inst_dmem_ram_1955, MEM_stage_inst_dmem_ram_1956, MEM_stage_inst_dmem_ram_1957, MEM_stage_inst_dmem_ram_1958, MEM_stage_inst_dmem_ram_1959, MEM_stage_inst_dmem_ram_1960, MEM_stage_inst_dmem_ram_1961, MEM_stage_inst_dmem_ram_1962, MEM_stage_inst_dmem_ram_1963, MEM_stage_inst_dmem_ram_1964, MEM_stage_inst_dmem_ram_1965, MEM_stage_inst_dmem_ram_1966, MEM_stage_inst_dmem_ram_1967, MEM_stage_inst_dmem_ram_1968, MEM_stage_inst_dmem_ram_1969, MEM_stage_inst_dmem_ram_1970, MEM_stage_inst_dmem_ram_1971, MEM_stage_inst_dmem_ram_1972, MEM_stage_inst_dmem_ram_1973, MEM_stage_inst_dmem_ram_1974, MEM_stage_inst_dmem_ram_1975, MEM_stage_inst_dmem_ram_1976, MEM_stage_inst_dmem_ram_1977, MEM_stage_inst_dmem_ram_1978, MEM_stage_inst_dmem_ram_1979, MEM_stage_inst_dmem_ram_1980, MEM_stage_inst_dmem_ram_1981, MEM_stage_inst_dmem_ram_1982, MEM_stage_inst_dmem_ram_1983, MEM_stage_inst_dmem_ram_1984, MEM_stage_inst_dmem_ram_1985, MEM_stage_inst_dmem_ram_1986, MEM_stage_inst_dmem_ram_1987, MEM_stage_inst_dmem_ram_1988, MEM_stage_inst_dmem_ram_1989, MEM_stage_inst_dmem_ram_1990, MEM_stage_inst_dmem_ram_1991, MEM_stage_inst_dmem_ram_1992, MEM_stage_inst_dmem_ram_1993, MEM_stage_inst_dmem_ram_1994, MEM_stage_inst_dmem_ram_1995, MEM_stage_inst_dmem_ram_1996, MEM_stage_inst_dmem_ram_1997, MEM_stage_inst_dmem_ram_1998, MEM_stage_inst_dmem_ram_1999, MEM_stage_inst_dmem_ram_2000, MEM_stage_inst_dmem_ram_2001, MEM_stage_inst_dmem_ram_2002, MEM_stage_inst_dmem_ram_2003, MEM_stage_inst_dmem_ram_2004, MEM_stage_inst_dmem_ram_2005, MEM_stage_inst_dmem_ram_2006, MEM_stage_inst_dmem_ram_2007, MEM_stage_inst_dmem_ram_2008, MEM_stage_inst_dmem_ram_2009, MEM_stage_inst_dmem_ram_2010, MEM_stage_inst_dmem_ram_2011, MEM_stage_inst_dmem_ram_2012, MEM_stage_inst_dmem_ram_2013, MEM_stage_inst_dmem_ram_2014, MEM_stage_inst_dmem_ram_2015, MEM_stage_inst_dmem_ram_2016, MEM_stage_inst_dmem_ram_2017, MEM_stage_inst_dmem_ram_2018, MEM_stage_inst_dmem_ram_2019, MEM_stage_inst_dmem_ram_2020, MEM_stage_inst_dmem_ram_2021, MEM_stage_inst_dmem_ram_2022, MEM_stage_inst_dmem_ram_2023, MEM_stage_inst_dmem_ram_2024, MEM_stage_inst_dmem_ram_2025, MEM_stage_inst_dmem_ram_2026, MEM_stage_inst_dmem_ram_2027, MEM_stage_inst_dmem_ram_2028, MEM_stage_inst_dmem_ram_2029, MEM_stage_inst_dmem_ram_2030, MEM_stage_inst_dmem_ram_2031, MEM_stage_inst_dmem_ram_2032, MEM_stage_inst_dmem_ram_2033, MEM_stage_inst_dmem_ram_2034, MEM_stage_inst_dmem_ram_2035, MEM_stage_inst_dmem_ram_2036, MEM_stage_inst_dmem_ram_2037, MEM_stage_inst_dmem_ram_2038, MEM_stage_inst_dmem_ram_2039, MEM_stage_inst_dmem_ram_2040, MEM_stage_inst_dmem_ram_2041, MEM_stage_inst_dmem_ram_2042, MEM_stage_inst_dmem_ram_2043, MEM_stage_inst_dmem_ram_2044, MEM_stage_inst_dmem_ram_2045, MEM_stage_inst_dmem_ram_2046, MEM_stage_inst_dmem_ram_2047, MEM_stage_inst_dmem_ram_1024, MEM_stage_inst_dmem_ram_1025, MEM_stage_inst_dmem_ram_1026, MEM_stage_inst_dmem_ram_1027, MEM_stage_inst_dmem_ram_1028, MEM_stage_inst_dmem_ram_1029, MEM_stage_inst_dmem_ram_1030, MEM_stage_inst_dmem_ram_1031, MEM_stage_inst_dmem_ram_1032, MEM_stage_inst_dmem_ram_1033, MEM_stage_inst_dmem_ram_1034, MEM_stage_inst_dmem_ram_1035, MEM_stage_inst_dmem_ram_1036, MEM_stage_inst_dmem_ram_1037, MEM_stage_inst_dmem_ram_1038, MEM_stage_inst_dmem_ram_1039, MEM_stage_inst_dmem_ram_1040, MEM_stage_inst_dmem_ram_1041, MEM_stage_inst_dmem_ram_1042, MEM_stage_inst_dmem_ram_1043, MEM_stage_inst_dmem_ram_1044, MEM_stage_inst_dmem_ram_1045, MEM_stage_inst_dmem_ram_1046, MEM_stage_inst_dmem_ram_1047, MEM_stage_inst_dmem_ram_1048, MEM_stage_inst_dmem_ram_1049, MEM_stage_inst_dmem_ram_1050, MEM_stage_inst_dmem_ram_1051, MEM_stage_inst_dmem_ram_1052, MEM_stage_inst_dmem_ram_1053, MEM_stage_inst_dmem_ram_1054, MEM_stage_inst_dmem_ram_1055, MEM_stage_inst_dmem_ram_1056, MEM_stage_inst_dmem_ram_1057, MEM_stage_inst_dmem_ram_1058, MEM_stage_inst_dmem_ram_1059, MEM_stage_inst_dmem_ram_1060, MEM_stage_inst_dmem_ram_1061, MEM_stage_inst_dmem_ram_1062, MEM_stage_inst_dmem_ram_1063, MEM_stage_inst_dmem_ram_1064, MEM_stage_inst_dmem_ram_1065, MEM_stage_inst_dmem_ram_1066, MEM_stage_inst_dmem_ram_1067, MEM_stage_inst_dmem_ram_1068, MEM_stage_inst_dmem_ram_1069, MEM_stage_inst_dmem_ram_1070, MEM_stage_inst_dmem_ram_1071, MEM_stage_inst_dmem_ram_1072, MEM_stage_inst_dmem_ram_1073, MEM_stage_inst_dmem_ram_1074, MEM_stage_inst_dmem_ram_1075, MEM_stage_inst_dmem_ram_1076, MEM_stage_inst_dmem_ram_1077, MEM_stage_inst_dmem_ram_1078, MEM_stage_inst_dmem_ram_1079, MEM_stage_inst_dmem_ram_1080, MEM_stage_inst_dmem_ram_1081, MEM_stage_inst_dmem_ram_1082, MEM_stage_inst_dmem_ram_1083, MEM_stage_inst_dmem_ram_1084, MEM_stage_inst_dmem_ram_1085, MEM_stage_inst_dmem_ram_1086, MEM_stage_inst_dmem_ram_1087, MEM_stage_inst_dmem_ram_1088, MEM_stage_inst_dmem_ram_1089, MEM_stage_inst_dmem_ram_1090, MEM_stage_inst_dmem_ram_1091, MEM_stage_inst_dmem_ram_1092, MEM_stage_inst_dmem_ram_1093, MEM_stage_inst_dmem_ram_1094, MEM_stage_inst_dmem_ram_1095, MEM_stage_inst_dmem_ram_1096, MEM_stage_inst_dmem_ram_1097, MEM_stage_inst_dmem_ram_1098, MEM_stage_inst_dmem_ram_1099, MEM_stage_inst_dmem_ram_1100, MEM_stage_inst_dmem_ram_1101, MEM_stage_inst_dmem_ram_1102, MEM_stage_inst_dmem_ram_1103, MEM_stage_inst_dmem_ram_1104, MEM_stage_inst_dmem_ram_1105, MEM_stage_inst_dmem_ram_1106, MEM_stage_inst_dmem_ram_1107, MEM_stage_inst_dmem_ram_1108, MEM_stage_inst_dmem_ram_1109, MEM_stage_inst_dmem_ram_1110, MEM_stage_inst_dmem_ram_1111, MEM_stage_inst_dmem_ram_1112, MEM_stage_inst_dmem_ram_1113, MEM_stage_inst_dmem_ram_1114, MEM_stage_inst_dmem_ram_1115, MEM_stage_inst_dmem_ram_1116, MEM_stage_inst_dmem_ram_1117, MEM_stage_inst_dmem_ram_1118, MEM_stage_inst_dmem_ram_1119, MEM_stage_inst_dmem_ram_1120, MEM_stage_inst_dmem_ram_1121, MEM_stage_inst_dmem_ram_1122, MEM_stage_inst_dmem_ram_1123, MEM_stage_inst_dmem_ram_1124, MEM_stage_inst_dmem_ram_1125, MEM_stage_inst_dmem_ram_1126, MEM_stage_inst_dmem_ram_1127, MEM_stage_inst_dmem_ram_1128, MEM_stage_inst_dmem_ram_1129, MEM_stage_inst_dmem_ram_1130, MEM_stage_inst_dmem_ram_1131, MEM_stage_inst_dmem_ram_1132, MEM_stage_inst_dmem_ram_1133, MEM_stage_inst_dmem_ram_1134, MEM_stage_inst_dmem_ram_1135, MEM_stage_inst_dmem_ram_1136, MEM_stage_inst_dmem_ram_1137, MEM_stage_inst_dmem_ram_1138, MEM_stage_inst_dmem_ram_1139, MEM_stage_inst_dmem_ram_1140, MEM_stage_inst_dmem_ram_1141, MEM_stage_inst_dmem_ram_1142, MEM_stage_inst_dmem_ram_1143, MEM_stage_inst_dmem_ram_1144, MEM_stage_inst_dmem_ram_1145, MEM_stage_inst_dmem_ram_1146, MEM_stage_inst_dmem_ram_1147, MEM_stage_inst_dmem_ram_1148, MEM_stage_inst_dmem_ram_1149, MEM_stage_inst_dmem_ram_1150, MEM_stage_inst_dmem_ram_1151, MEM_stage_inst_dmem_ram_1152, MEM_stage_inst_dmem_ram_1153, MEM_stage_inst_dmem_ram_1154, MEM_stage_inst_dmem_ram_1155, MEM_stage_inst_dmem_ram_1156, MEM_stage_inst_dmem_ram_1157, MEM_stage_inst_dmem_ram_1158, MEM_stage_inst_dmem_ram_1159, MEM_stage_inst_dmem_ram_1160, MEM_stage_inst_dmem_ram_1161, MEM_stage_inst_dmem_ram_1162, MEM_stage_inst_dmem_ram_1163, MEM_stage_inst_dmem_ram_1164, MEM_stage_inst_dmem_ram_1165, MEM_stage_inst_dmem_ram_1166, MEM_stage_inst_dmem_ram_1167, MEM_stage_inst_dmem_ram_1168, MEM_stage_inst_dmem_ram_1169, MEM_stage_inst_dmem_ram_1170, MEM_stage_inst_dmem_ram_1171, MEM_stage_inst_dmem_ram_1172, MEM_stage_inst_dmem_ram_1173, MEM_stage_inst_dmem_ram_1174, MEM_stage_inst_dmem_ram_1175, MEM_stage_inst_dmem_ram_1176, MEM_stage_inst_dmem_ram_1177, MEM_stage_inst_dmem_ram_1178, MEM_stage_inst_dmem_ram_1179, MEM_stage_inst_dmem_ram_1180, MEM_stage_inst_dmem_ram_1181, MEM_stage_inst_dmem_ram_1182, MEM_stage_inst_dmem_ram_1183, MEM_stage_inst_dmem_ram_1184, MEM_stage_inst_dmem_ram_1185, MEM_stage_inst_dmem_ram_1186, MEM_stage_inst_dmem_ram_1187, MEM_stage_inst_dmem_ram_1188, MEM_stage_inst_dmem_ram_1189, MEM_stage_inst_dmem_ram_1190, MEM_stage_inst_dmem_ram_1191, MEM_stage_inst_dmem_ram_1192, MEM_stage_inst_dmem_ram_1193, MEM_stage_inst_dmem_ram_1194, MEM_stage_inst_dmem_ram_1195, MEM_stage_inst_dmem_ram_1196, MEM_stage_inst_dmem_ram_1197, MEM_stage_inst_dmem_ram_1198, MEM_stage_inst_dmem_ram_1199, MEM_stage_inst_dmem_ram_1200, MEM_stage_inst_dmem_ram_1201, MEM_stage_inst_dmem_ram_1202, MEM_stage_inst_dmem_ram_1203, MEM_stage_inst_dmem_ram_1204, MEM_stage_inst_dmem_ram_1205, MEM_stage_inst_dmem_ram_1206, MEM_stage_inst_dmem_ram_1207, MEM_stage_inst_dmem_ram_1208, MEM_stage_inst_dmem_ram_1209, MEM_stage_inst_dmem_ram_1210, MEM_stage_inst_dmem_ram_1211, MEM_stage_inst_dmem_ram_1212, MEM_stage_inst_dmem_ram_1213, MEM_stage_inst_dmem_ram_1214, MEM_stage_inst_dmem_ram_1215, MEM_stage_inst_dmem_ram_1216, MEM_stage_inst_dmem_ram_1217, MEM_stage_inst_dmem_ram_1218, MEM_stage_inst_dmem_ram_1219, MEM_stage_inst_dmem_ram_1220, MEM_stage_inst_dmem_ram_1221, MEM_stage_inst_dmem_ram_1222, MEM_stage_inst_dmem_ram_1223, MEM_stage_inst_dmem_ram_1224, MEM_stage_inst_dmem_ram_1225, MEM_stage_inst_dmem_ram_1226, MEM_stage_inst_dmem_ram_1227, MEM_stage_inst_dmem_ram_1228, MEM_stage_inst_dmem_ram_1229, MEM_stage_inst_dmem_ram_1230, MEM_stage_inst_dmem_ram_1231, MEM_stage_inst_dmem_ram_1232, MEM_stage_inst_dmem_ram_1233, MEM_stage_inst_dmem_ram_1234, MEM_stage_inst_dmem_ram_1235, MEM_stage_inst_dmem_ram_1236, MEM_stage_inst_dmem_ram_1237, MEM_stage_inst_dmem_ram_1238, MEM_stage_inst_dmem_ram_1239, MEM_stage_inst_dmem_ram_1240, MEM_stage_inst_dmem_ram_1241, MEM_stage_inst_dmem_ram_1242, MEM_stage_inst_dmem_ram_1243, MEM_stage_inst_dmem_ram_1244, MEM_stage_inst_dmem_ram_1245, MEM_stage_inst_dmem_ram_1246, MEM_stage_inst_dmem_ram_1247, MEM_stage_inst_dmem_ram_1248, MEM_stage_inst_dmem_ram_1249, MEM_stage_inst_dmem_ram_1250, MEM_stage_inst_dmem_ram_1251, MEM_stage_inst_dmem_ram_1252, MEM_stage_inst_dmem_ram_1253, MEM_stage_inst_dmem_ram_1254, MEM_stage_inst_dmem_ram_1255, MEM_stage_inst_dmem_ram_1256, MEM_stage_inst_dmem_ram_1257, MEM_stage_inst_dmem_ram_1258, MEM_stage_inst_dmem_ram_1259, MEM_stage_inst_dmem_ram_1260, MEM_stage_inst_dmem_ram_1261, MEM_stage_inst_dmem_ram_1262, MEM_stage_inst_dmem_ram_1263, MEM_stage_inst_dmem_ram_1264, MEM_stage_inst_dmem_ram_1265, MEM_stage_inst_dmem_ram_1266, MEM_stage_inst_dmem_ram_1267, MEM_stage_inst_dmem_ram_1268, MEM_stage_inst_dmem_ram_1269, MEM_stage_inst_dmem_ram_1270, MEM_stage_inst_dmem_ram_1271, MEM_stage_inst_dmem_ram_1272, MEM_stage_inst_dmem_ram_1273, MEM_stage_inst_dmem_ram_1274, MEM_stage_inst_dmem_ram_1275, MEM_stage_inst_dmem_ram_1276, MEM_stage_inst_dmem_ram_1277, MEM_stage_inst_dmem_ram_1278, MEM_stage_inst_dmem_ram_1279, MEM_stage_inst_dmem_ram_1280, MEM_stage_inst_dmem_ram_1281, MEM_stage_inst_dmem_ram_1282, MEM_stage_inst_dmem_ram_1283, MEM_stage_inst_dmem_ram_1284, MEM_stage_inst_dmem_ram_1285, MEM_stage_inst_dmem_ram_1286, MEM_stage_inst_dmem_ram_1287, MEM_stage_inst_dmem_ram_1288, MEM_stage_inst_dmem_ram_1289, MEM_stage_inst_dmem_ram_1290, MEM_stage_inst_dmem_ram_1291, MEM_stage_inst_dmem_ram_1292, MEM_stage_inst_dmem_ram_1293, MEM_stage_inst_dmem_ram_1294, MEM_stage_inst_dmem_ram_1295, MEM_stage_inst_dmem_ram_1296, MEM_stage_inst_dmem_ram_1297, MEM_stage_inst_dmem_ram_1298, MEM_stage_inst_dmem_ram_1299, MEM_stage_inst_dmem_ram_1300, MEM_stage_inst_dmem_ram_1301, MEM_stage_inst_dmem_ram_1302, MEM_stage_inst_dmem_ram_1303, MEM_stage_inst_dmem_ram_1304, MEM_stage_inst_dmem_ram_1305, MEM_stage_inst_dmem_ram_1306, MEM_stage_inst_dmem_ram_1307, MEM_stage_inst_dmem_ram_1308, MEM_stage_inst_dmem_ram_1309, MEM_stage_inst_dmem_ram_1310, MEM_stage_inst_dmem_ram_1311, MEM_stage_inst_dmem_ram_1312, MEM_stage_inst_dmem_ram_1313, MEM_stage_inst_dmem_ram_1314, MEM_stage_inst_dmem_ram_1315, MEM_stage_inst_dmem_ram_1316, MEM_stage_inst_dmem_ram_1317, MEM_stage_inst_dmem_ram_1318, MEM_stage_inst_dmem_ram_1319, MEM_stage_inst_dmem_ram_1320, MEM_stage_inst_dmem_ram_1321, MEM_stage_inst_dmem_ram_1322, MEM_stage_inst_dmem_ram_1323, MEM_stage_inst_dmem_ram_1324, MEM_stage_inst_dmem_ram_1325, MEM_stage_inst_dmem_ram_1326, MEM_stage_inst_dmem_ram_1327, MEM_stage_inst_dmem_ram_1328, MEM_stage_inst_dmem_ram_1329, MEM_stage_inst_dmem_ram_1330, MEM_stage_inst_dmem_ram_1331, MEM_stage_inst_dmem_ram_1332, MEM_stage_inst_dmem_ram_1333, MEM_stage_inst_dmem_ram_1334, MEM_stage_inst_dmem_ram_1335, MEM_stage_inst_dmem_ram_1336, MEM_stage_inst_dmem_ram_1337, MEM_stage_inst_dmem_ram_1338, MEM_stage_inst_dmem_ram_1339, MEM_stage_inst_dmem_ram_1340, MEM_stage_inst_dmem_ram_1341, MEM_stage_inst_dmem_ram_1342, MEM_stage_inst_dmem_ram_1343, MEM_stage_inst_dmem_ram_1344, MEM_stage_inst_dmem_ram_1345, MEM_stage_inst_dmem_ram_1346, MEM_stage_inst_dmem_ram_1347, MEM_stage_inst_dmem_ram_1348, MEM_stage_inst_dmem_ram_1349, MEM_stage_inst_dmem_ram_1350, MEM_stage_inst_dmem_ram_1351, MEM_stage_inst_dmem_ram_1352, MEM_stage_inst_dmem_ram_1353, MEM_stage_inst_dmem_ram_1354, MEM_stage_inst_dmem_ram_1355, MEM_stage_inst_dmem_ram_1356, MEM_stage_inst_dmem_ram_1357, MEM_stage_inst_dmem_ram_1358, MEM_stage_inst_dmem_ram_1359, MEM_stage_inst_dmem_ram_1360, MEM_stage_inst_dmem_ram_1361, MEM_stage_inst_dmem_ram_1362, MEM_stage_inst_dmem_ram_1363, MEM_stage_inst_dmem_ram_1364, MEM_stage_inst_dmem_ram_1365, MEM_stage_inst_dmem_ram_1366, MEM_stage_inst_dmem_ram_1367, MEM_stage_inst_dmem_ram_1368, MEM_stage_inst_dmem_ram_1369, MEM_stage_inst_dmem_ram_1370, MEM_stage_inst_dmem_ram_1371, MEM_stage_inst_dmem_ram_1372, MEM_stage_inst_dmem_ram_1373, MEM_stage_inst_dmem_ram_1374, MEM_stage_inst_dmem_ram_1375, MEM_stage_inst_dmem_ram_1376, MEM_stage_inst_dmem_ram_1377, MEM_stage_inst_dmem_ram_1378, MEM_stage_inst_dmem_ram_1379, MEM_stage_inst_dmem_ram_1380, MEM_stage_inst_dmem_ram_1381, MEM_stage_inst_dmem_ram_1382, MEM_stage_inst_dmem_ram_1383, MEM_stage_inst_dmem_ram_1384, MEM_stage_inst_dmem_ram_1385, MEM_stage_inst_dmem_ram_1386, MEM_stage_inst_dmem_ram_1387, MEM_stage_inst_dmem_ram_1388, MEM_stage_inst_dmem_ram_1389, MEM_stage_inst_dmem_ram_1390, MEM_stage_inst_dmem_ram_1391, MEM_stage_inst_dmem_ram_1392, MEM_stage_inst_dmem_ram_1393, MEM_stage_inst_dmem_ram_1394, MEM_stage_inst_dmem_ram_1395, MEM_stage_inst_dmem_ram_1396, MEM_stage_inst_dmem_ram_1397, MEM_stage_inst_dmem_ram_1398, MEM_stage_inst_dmem_ram_1399, MEM_stage_inst_dmem_ram_1400, MEM_stage_inst_dmem_ram_1401, MEM_stage_inst_dmem_ram_1402, MEM_stage_inst_dmem_ram_1403, MEM_stage_inst_dmem_ram_1404, MEM_stage_inst_dmem_ram_1405, MEM_stage_inst_dmem_ram_1406, MEM_stage_inst_dmem_ram_1407, MEM_stage_inst_dmem_ram_1408, MEM_stage_inst_dmem_ram_1409, MEM_stage_inst_dmem_ram_1410, MEM_stage_inst_dmem_ram_1411, MEM_stage_inst_dmem_ram_1412, MEM_stage_inst_dmem_ram_1413, MEM_stage_inst_dmem_ram_1414, MEM_stage_inst_dmem_ram_1415, MEM_stage_inst_dmem_ram_1416, MEM_stage_inst_dmem_ram_1417, MEM_stage_inst_dmem_ram_1418, MEM_stage_inst_dmem_ram_1419, MEM_stage_inst_dmem_ram_1420, MEM_stage_inst_dmem_ram_1421, MEM_stage_inst_dmem_ram_1422, MEM_stage_inst_dmem_ram_1423, MEM_stage_inst_dmem_ram_1424, MEM_stage_inst_dmem_ram_1425, MEM_stage_inst_dmem_ram_1426, MEM_stage_inst_dmem_ram_1427, MEM_stage_inst_dmem_ram_1428, MEM_stage_inst_dmem_ram_1429, MEM_stage_inst_dmem_ram_1430, MEM_stage_inst_dmem_ram_1431, MEM_stage_inst_dmem_ram_1432, MEM_stage_inst_dmem_ram_1433, MEM_stage_inst_dmem_ram_1434, MEM_stage_inst_dmem_ram_1435, MEM_stage_inst_dmem_ram_1436, MEM_stage_inst_dmem_ram_1437, MEM_stage_inst_dmem_ram_1438, MEM_stage_inst_dmem_ram_1439, MEM_stage_inst_dmem_ram_1440, MEM_stage_inst_dmem_ram_1441, MEM_stage_inst_dmem_ram_1442, MEM_stage_inst_dmem_ram_1443, MEM_stage_inst_dmem_ram_1444, MEM_stage_inst_dmem_ram_1445, MEM_stage_inst_dmem_ram_1446, MEM_stage_inst_dmem_ram_1447, MEM_stage_inst_dmem_ram_1448, MEM_stage_inst_dmem_ram_1449, MEM_stage_inst_dmem_ram_1450, MEM_stage_inst_dmem_ram_1451, MEM_stage_inst_dmem_ram_1452, MEM_stage_inst_dmem_ram_1453, MEM_stage_inst_dmem_ram_1454, MEM_stage_inst_dmem_ram_1455, MEM_stage_inst_dmem_ram_1456, MEM_stage_inst_dmem_ram_1457, MEM_stage_inst_dmem_ram_1458, MEM_stage_inst_dmem_ram_1459, MEM_stage_inst_dmem_ram_1460, MEM_stage_inst_dmem_ram_1461, MEM_stage_inst_dmem_ram_1462, MEM_stage_inst_dmem_ram_1463, MEM_stage_inst_dmem_ram_1464, MEM_stage_inst_dmem_ram_1465, MEM_stage_inst_dmem_ram_1466, MEM_stage_inst_dmem_ram_1467, MEM_stage_inst_dmem_ram_1468, MEM_stage_inst_dmem_ram_1469, MEM_stage_inst_dmem_ram_1470, MEM_stage_inst_dmem_ram_1471, MEM_stage_inst_dmem_ram_1472, MEM_stage_inst_dmem_ram_1473, MEM_stage_inst_dmem_ram_1474, MEM_stage_inst_dmem_ram_1475, MEM_stage_inst_dmem_ram_1476, MEM_stage_inst_dmem_ram_1477, MEM_stage_inst_dmem_ram_1478, MEM_stage_inst_dmem_ram_1479, MEM_stage_inst_dmem_ram_1480, MEM_stage_inst_dmem_ram_1481, MEM_stage_inst_dmem_ram_1482, MEM_stage_inst_dmem_ram_1483, MEM_stage_inst_dmem_ram_1484, MEM_stage_inst_dmem_ram_1485, MEM_stage_inst_dmem_ram_1486, MEM_stage_inst_dmem_ram_1487, MEM_stage_inst_dmem_ram_1488, MEM_stage_inst_dmem_ram_1489, MEM_stage_inst_dmem_ram_1490, MEM_stage_inst_dmem_ram_1491, MEM_stage_inst_dmem_ram_1492, MEM_stage_inst_dmem_ram_1493, MEM_stage_inst_dmem_ram_1494, MEM_stage_inst_dmem_ram_1495, MEM_stage_inst_dmem_ram_1496, MEM_stage_inst_dmem_ram_1497, MEM_stage_inst_dmem_ram_1498, MEM_stage_inst_dmem_ram_1499, MEM_stage_inst_dmem_ram_1500, MEM_stage_inst_dmem_ram_1501, MEM_stage_inst_dmem_ram_1502, MEM_stage_inst_dmem_ram_1503, MEM_stage_inst_dmem_ram_1504, MEM_stage_inst_dmem_ram_1505, MEM_stage_inst_dmem_ram_1506, MEM_stage_inst_dmem_ram_1507, MEM_stage_inst_dmem_ram_1508, MEM_stage_inst_dmem_ram_1509, MEM_stage_inst_dmem_ram_1510, MEM_stage_inst_dmem_ram_1511, MEM_stage_inst_dmem_ram_1512, MEM_stage_inst_dmem_ram_1513, MEM_stage_inst_dmem_ram_1514, MEM_stage_inst_dmem_ram_1515, MEM_stage_inst_dmem_ram_1516, MEM_stage_inst_dmem_ram_1517, MEM_stage_inst_dmem_ram_1518, MEM_stage_inst_dmem_ram_1519, MEM_stage_inst_dmem_ram_1520, MEM_stage_inst_dmem_ram_1521, MEM_stage_inst_dmem_ram_1522, MEM_stage_inst_dmem_ram_1523, MEM_stage_inst_dmem_ram_1524, MEM_stage_inst_dmem_ram_1525, MEM_stage_inst_dmem_ram_1526, MEM_stage_inst_dmem_ram_1527, MEM_stage_inst_dmem_ram_1528, MEM_stage_inst_dmem_ram_1529, MEM_stage_inst_dmem_ram_1530, MEM_stage_inst_dmem_ram_1531, MEM_stage_inst_dmem_ram_1532, MEM_stage_inst_dmem_ram_1533, MEM_stage_inst_dmem_ram_1534, MEM_stage_inst_dmem_ram_1535, MEM_stage_inst_dmem_ram_512, MEM_stage_inst_dmem_ram_513, MEM_stage_inst_dmem_ram_514, MEM_stage_inst_dmem_ram_515, MEM_stage_inst_dmem_ram_516, MEM_stage_inst_dmem_ram_517, MEM_stage_inst_dmem_ram_518, MEM_stage_inst_dmem_ram_519, MEM_stage_inst_dmem_ram_520, MEM_stage_inst_dmem_ram_521, MEM_stage_inst_dmem_ram_522, MEM_stage_inst_dmem_ram_523, MEM_stage_inst_dmem_ram_524, MEM_stage_inst_dmem_ram_525, MEM_stage_inst_dmem_ram_526, MEM_stage_inst_dmem_ram_527, MEM_stage_inst_dmem_ram_528, MEM_stage_inst_dmem_ram_529, MEM_stage_inst_dmem_ram_530, MEM_stage_inst_dmem_ram_531, MEM_stage_inst_dmem_ram_532, MEM_stage_inst_dmem_ram_533, MEM_stage_inst_dmem_ram_534, MEM_stage_inst_dmem_ram_535, MEM_stage_inst_dmem_ram_536, MEM_stage_inst_dmem_ram_537, MEM_stage_inst_dmem_ram_538, MEM_stage_inst_dmem_ram_539, MEM_stage_inst_dmem_ram_540, MEM_stage_inst_dmem_ram_541, MEM_stage_inst_dmem_ram_542, MEM_stage_inst_dmem_ram_543, MEM_stage_inst_dmem_ram_544, MEM_stage_inst_dmem_ram_545, MEM_stage_inst_dmem_ram_546, MEM_stage_inst_dmem_ram_547, MEM_stage_inst_dmem_ram_548, MEM_stage_inst_dmem_ram_549, MEM_stage_inst_dmem_ram_550, MEM_stage_inst_dmem_ram_551, MEM_stage_inst_dmem_ram_552, MEM_stage_inst_dmem_ram_553, MEM_stage_inst_dmem_ram_554, MEM_stage_inst_dmem_ram_555, MEM_stage_inst_dmem_ram_556, MEM_stage_inst_dmem_ram_557, MEM_stage_inst_dmem_ram_558, MEM_stage_inst_dmem_ram_559, MEM_stage_inst_dmem_ram_560, MEM_stage_inst_dmem_ram_561, MEM_stage_inst_dmem_ram_562, MEM_stage_inst_dmem_ram_563, MEM_stage_inst_dmem_ram_564, MEM_stage_inst_dmem_ram_565, MEM_stage_inst_dmem_ram_566, MEM_stage_inst_dmem_ram_567, MEM_stage_inst_dmem_ram_568, MEM_stage_inst_dmem_ram_569, MEM_stage_inst_dmem_ram_570, MEM_stage_inst_dmem_ram_571, MEM_stage_inst_dmem_ram_572, MEM_stage_inst_dmem_ram_573, MEM_stage_inst_dmem_ram_574, MEM_stage_inst_dmem_ram_575, MEM_stage_inst_dmem_ram_576, MEM_stage_inst_dmem_ram_577, MEM_stage_inst_dmem_ram_578, MEM_stage_inst_dmem_ram_579, MEM_stage_inst_dmem_ram_580, MEM_stage_inst_dmem_ram_581, MEM_stage_inst_dmem_ram_582, MEM_stage_inst_dmem_ram_583, MEM_stage_inst_dmem_ram_584, MEM_stage_inst_dmem_ram_585, MEM_stage_inst_dmem_ram_586, MEM_stage_inst_dmem_ram_587, MEM_stage_inst_dmem_ram_588, MEM_stage_inst_dmem_ram_589, MEM_stage_inst_dmem_ram_590, MEM_stage_inst_dmem_ram_591, MEM_stage_inst_dmem_ram_592, MEM_stage_inst_dmem_ram_593, MEM_stage_inst_dmem_ram_594, MEM_stage_inst_dmem_ram_595, MEM_stage_inst_dmem_ram_596, MEM_stage_inst_dmem_ram_597, MEM_stage_inst_dmem_ram_598, MEM_stage_inst_dmem_ram_599, MEM_stage_inst_dmem_ram_600, MEM_stage_inst_dmem_ram_601, MEM_stage_inst_dmem_ram_602, MEM_stage_inst_dmem_ram_603, MEM_stage_inst_dmem_ram_604, MEM_stage_inst_dmem_ram_605, MEM_stage_inst_dmem_ram_606, MEM_stage_inst_dmem_ram_607, MEM_stage_inst_dmem_ram_608, MEM_stage_inst_dmem_ram_609, MEM_stage_inst_dmem_ram_610, MEM_stage_inst_dmem_ram_611, MEM_stage_inst_dmem_ram_612, MEM_stage_inst_dmem_ram_613, MEM_stage_inst_dmem_ram_614, MEM_stage_inst_dmem_ram_615, MEM_stage_inst_dmem_ram_616, MEM_stage_inst_dmem_ram_617, MEM_stage_inst_dmem_ram_618, MEM_stage_inst_dmem_ram_619, MEM_stage_inst_dmem_ram_620, MEM_stage_inst_dmem_ram_621, MEM_stage_inst_dmem_ram_622, MEM_stage_inst_dmem_ram_623, MEM_stage_inst_dmem_ram_624, MEM_stage_inst_dmem_ram_625, MEM_stage_inst_dmem_ram_626, MEM_stage_inst_dmem_ram_627, MEM_stage_inst_dmem_ram_628, MEM_stage_inst_dmem_ram_629, MEM_stage_inst_dmem_ram_630, MEM_stage_inst_dmem_ram_631, MEM_stage_inst_dmem_ram_632, MEM_stage_inst_dmem_ram_633, MEM_stage_inst_dmem_ram_634, MEM_stage_inst_dmem_ram_635, MEM_stage_inst_dmem_ram_636, MEM_stage_inst_dmem_ram_637, MEM_stage_inst_dmem_ram_638, MEM_stage_inst_dmem_ram_639, MEM_stage_inst_dmem_ram_640, MEM_stage_inst_dmem_ram_641, MEM_stage_inst_dmem_ram_642, MEM_stage_inst_dmem_ram_643, MEM_stage_inst_dmem_ram_644, MEM_stage_inst_dmem_ram_645, MEM_stage_inst_dmem_ram_646, MEM_stage_inst_dmem_ram_647, MEM_stage_inst_dmem_ram_648, MEM_stage_inst_dmem_ram_649, MEM_stage_inst_dmem_ram_650, MEM_stage_inst_dmem_ram_651, MEM_stage_inst_dmem_ram_652, MEM_stage_inst_dmem_ram_653, MEM_stage_inst_dmem_ram_654, MEM_stage_inst_dmem_ram_655, MEM_stage_inst_dmem_ram_656, MEM_stage_inst_dmem_ram_657, MEM_stage_inst_dmem_ram_658, MEM_stage_inst_dmem_ram_659, MEM_stage_inst_dmem_ram_660, MEM_stage_inst_dmem_ram_661, MEM_stage_inst_dmem_ram_662, MEM_stage_inst_dmem_ram_663, MEM_stage_inst_dmem_ram_664, MEM_stage_inst_dmem_ram_665, MEM_stage_inst_dmem_ram_666, MEM_stage_inst_dmem_ram_667, MEM_stage_inst_dmem_ram_668, MEM_stage_inst_dmem_ram_669, MEM_stage_inst_dmem_ram_670, MEM_stage_inst_dmem_ram_671, MEM_stage_inst_dmem_ram_672, MEM_stage_inst_dmem_ram_673, MEM_stage_inst_dmem_ram_674, MEM_stage_inst_dmem_ram_675, MEM_stage_inst_dmem_ram_676, MEM_stage_inst_dmem_ram_677, MEM_stage_inst_dmem_ram_678, MEM_stage_inst_dmem_ram_679, MEM_stage_inst_dmem_ram_680, MEM_stage_inst_dmem_ram_681, MEM_stage_inst_dmem_ram_682, MEM_stage_inst_dmem_ram_683, MEM_stage_inst_dmem_ram_684, MEM_stage_inst_dmem_ram_685, MEM_stage_inst_dmem_ram_686, MEM_stage_inst_dmem_ram_687, MEM_stage_inst_dmem_ram_688, MEM_stage_inst_dmem_ram_689, MEM_stage_inst_dmem_ram_690, MEM_stage_inst_dmem_ram_691, MEM_stage_inst_dmem_ram_692, MEM_stage_inst_dmem_ram_693, MEM_stage_inst_dmem_ram_694, MEM_stage_inst_dmem_ram_695, MEM_stage_inst_dmem_ram_696, MEM_stage_inst_dmem_ram_697, MEM_stage_inst_dmem_ram_698, MEM_stage_inst_dmem_ram_699, MEM_stage_inst_dmem_ram_700, MEM_stage_inst_dmem_ram_701, MEM_stage_inst_dmem_ram_702, MEM_stage_inst_dmem_ram_703, MEM_stage_inst_dmem_ram_704, MEM_stage_inst_dmem_ram_705, MEM_stage_inst_dmem_ram_706, MEM_stage_inst_dmem_ram_707, MEM_stage_inst_dmem_ram_708, MEM_stage_inst_dmem_ram_709, MEM_stage_inst_dmem_ram_710, MEM_stage_inst_dmem_ram_711, MEM_stage_inst_dmem_ram_712, MEM_stage_inst_dmem_ram_713, MEM_stage_inst_dmem_ram_714, MEM_stage_inst_dmem_ram_715, MEM_stage_inst_dmem_ram_716, MEM_stage_inst_dmem_ram_717, MEM_stage_inst_dmem_ram_718, MEM_stage_inst_dmem_ram_719, MEM_stage_inst_dmem_ram_720, MEM_stage_inst_dmem_ram_721, MEM_stage_inst_dmem_ram_722, MEM_stage_inst_dmem_ram_723, MEM_stage_inst_dmem_ram_724, MEM_stage_inst_dmem_ram_725, MEM_stage_inst_dmem_ram_726, MEM_stage_inst_dmem_ram_727, MEM_stage_inst_dmem_ram_728, MEM_stage_inst_dmem_ram_729, MEM_stage_inst_dmem_ram_730, MEM_stage_inst_dmem_ram_731, MEM_stage_inst_dmem_ram_732, MEM_stage_inst_dmem_ram_733, MEM_stage_inst_dmem_ram_734, MEM_stage_inst_dmem_ram_735, MEM_stage_inst_dmem_ram_736, MEM_stage_inst_dmem_ram_737, MEM_stage_inst_dmem_ram_738, MEM_stage_inst_dmem_ram_739, MEM_stage_inst_dmem_ram_740, MEM_stage_inst_dmem_ram_741, MEM_stage_inst_dmem_ram_742, MEM_stage_inst_dmem_ram_743, MEM_stage_inst_dmem_ram_744, MEM_stage_inst_dmem_ram_745, MEM_stage_inst_dmem_ram_746, MEM_stage_inst_dmem_ram_747, MEM_stage_inst_dmem_ram_748, MEM_stage_inst_dmem_ram_749, MEM_stage_inst_dmem_ram_750, MEM_stage_inst_dmem_ram_751, MEM_stage_inst_dmem_ram_752, MEM_stage_inst_dmem_ram_753, MEM_stage_inst_dmem_ram_754, MEM_stage_inst_dmem_ram_755, MEM_stage_inst_dmem_ram_756, MEM_stage_inst_dmem_ram_757, MEM_stage_inst_dmem_ram_758, MEM_stage_inst_dmem_ram_759, MEM_stage_inst_dmem_ram_760, MEM_stage_inst_dmem_ram_761, MEM_stage_inst_dmem_ram_762, MEM_stage_inst_dmem_ram_763, MEM_stage_inst_dmem_ram_764, MEM_stage_inst_dmem_ram_765, MEM_stage_inst_dmem_ram_766, MEM_stage_inst_dmem_ram_767, MEM_stage_inst_dmem_ram_768, MEM_stage_inst_dmem_ram_769, MEM_stage_inst_dmem_ram_770, MEM_stage_inst_dmem_ram_771, MEM_stage_inst_dmem_ram_772, MEM_stage_inst_dmem_ram_773, MEM_stage_inst_dmem_ram_774, MEM_stage_inst_dmem_ram_775, MEM_stage_inst_dmem_ram_776, MEM_stage_inst_dmem_ram_777, MEM_stage_inst_dmem_ram_778, MEM_stage_inst_dmem_ram_779, MEM_stage_inst_dmem_ram_780, MEM_stage_inst_dmem_ram_781, MEM_stage_inst_dmem_ram_782, MEM_stage_inst_dmem_ram_783, MEM_stage_inst_dmem_ram_784, MEM_stage_inst_dmem_ram_785, MEM_stage_inst_dmem_ram_786, MEM_stage_inst_dmem_ram_787, MEM_stage_inst_dmem_ram_788, MEM_stage_inst_dmem_ram_789, MEM_stage_inst_dmem_ram_790, MEM_stage_inst_dmem_ram_791, MEM_stage_inst_dmem_ram_792, MEM_stage_inst_dmem_ram_793, MEM_stage_inst_dmem_ram_794, MEM_stage_inst_dmem_ram_795, MEM_stage_inst_dmem_ram_796, MEM_stage_inst_dmem_ram_797, MEM_stage_inst_dmem_ram_798, MEM_stage_inst_dmem_ram_799, MEM_stage_inst_dmem_ram_800, MEM_stage_inst_dmem_ram_801, MEM_stage_inst_dmem_ram_802, MEM_stage_inst_dmem_ram_803, MEM_stage_inst_dmem_ram_804, MEM_stage_inst_dmem_ram_805, MEM_stage_inst_dmem_ram_806, MEM_stage_inst_dmem_ram_807, MEM_stage_inst_dmem_ram_808, MEM_stage_inst_dmem_ram_809, MEM_stage_inst_dmem_ram_810, MEM_stage_inst_dmem_ram_811, MEM_stage_inst_dmem_ram_812, MEM_stage_inst_dmem_ram_813, MEM_stage_inst_dmem_ram_814, MEM_stage_inst_dmem_ram_815, MEM_stage_inst_dmem_ram_816, MEM_stage_inst_dmem_ram_817, MEM_stage_inst_dmem_ram_818, MEM_stage_inst_dmem_ram_819, MEM_stage_inst_dmem_ram_820, MEM_stage_inst_dmem_ram_821, MEM_stage_inst_dmem_ram_822, MEM_stage_inst_dmem_ram_823, MEM_stage_inst_dmem_ram_824, MEM_stage_inst_dmem_ram_825, MEM_stage_inst_dmem_ram_826, MEM_stage_inst_dmem_ram_827, MEM_stage_inst_dmem_ram_828, MEM_stage_inst_dmem_ram_829, MEM_stage_inst_dmem_ram_830, MEM_stage_inst_dmem_ram_831, MEM_stage_inst_dmem_ram_832, MEM_stage_inst_dmem_ram_833, MEM_stage_inst_dmem_ram_834, MEM_stage_inst_dmem_ram_835, MEM_stage_inst_dmem_ram_836, MEM_stage_inst_dmem_ram_837, MEM_stage_inst_dmem_ram_838, MEM_stage_inst_dmem_ram_839, MEM_stage_inst_dmem_ram_840, MEM_stage_inst_dmem_ram_841, MEM_stage_inst_dmem_ram_842, MEM_stage_inst_dmem_ram_843, MEM_stage_inst_dmem_ram_844, MEM_stage_inst_dmem_ram_845, MEM_stage_inst_dmem_ram_846, MEM_stage_inst_dmem_ram_847, MEM_stage_inst_dmem_ram_848, MEM_stage_inst_dmem_ram_849, MEM_stage_inst_dmem_ram_850, MEM_stage_inst_dmem_ram_851, MEM_stage_inst_dmem_ram_852, MEM_stage_inst_dmem_ram_853, MEM_stage_inst_dmem_ram_854, MEM_stage_inst_dmem_ram_855, MEM_stage_inst_dmem_ram_856, MEM_stage_inst_dmem_ram_857, MEM_stage_inst_dmem_ram_858, MEM_stage_inst_dmem_ram_859, MEM_stage_inst_dmem_ram_860, MEM_stage_inst_dmem_ram_861, MEM_stage_inst_dmem_ram_862, MEM_stage_inst_dmem_ram_863, MEM_stage_inst_dmem_ram_864, MEM_stage_inst_dmem_ram_865, MEM_stage_inst_dmem_ram_866, MEM_stage_inst_dmem_ram_867, MEM_stage_inst_dmem_ram_868, MEM_stage_inst_dmem_ram_869, MEM_stage_inst_dmem_ram_870, MEM_stage_inst_dmem_ram_871, MEM_stage_inst_dmem_ram_872, MEM_stage_inst_dmem_ram_873, MEM_stage_inst_dmem_ram_874, MEM_stage_inst_dmem_ram_875, MEM_stage_inst_dmem_ram_876, MEM_stage_inst_dmem_ram_877, MEM_stage_inst_dmem_ram_878, MEM_stage_inst_dmem_ram_879, MEM_stage_inst_dmem_ram_880, MEM_stage_inst_dmem_ram_881, MEM_stage_inst_dmem_ram_882, MEM_stage_inst_dmem_ram_883, MEM_stage_inst_dmem_ram_884, MEM_stage_inst_dmem_ram_885, MEM_stage_inst_dmem_ram_886, MEM_stage_inst_dmem_ram_887, MEM_stage_inst_dmem_ram_888, MEM_stage_inst_dmem_ram_889, MEM_stage_inst_dmem_ram_890, MEM_stage_inst_dmem_ram_891, MEM_stage_inst_dmem_ram_892, MEM_stage_inst_dmem_ram_893, MEM_stage_inst_dmem_ram_894, MEM_stage_inst_dmem_ram_895, MEM_stage_inst_dmem_ram_896, MEM_stage_inst_dmem_ram_897, MEM_stage_inst_dmem_ram_898, MEM_stage_inst_dmem_ram_899, MEM_stage_inst_dmem_ram_900, MEM_stage_inst_dmem_ram_901, MEM_stage_inst_dmem_ram_902, MEM_stage_inst_dmem_ram_903, MEM_stage_inst_dmem_ram_904, MEM_stage_inst_dmem_ram_905, MEM_stage_inst_dmem_ram_906, MEM_stage_inst_dmem_ram_907, MEM_stage_inst_dmem_ram_908, MEM_stage_inst_dmem_ram_909, MEM_stage_inst_dmem_ram_910, MEM_stage_inst_dmem_ram_911, MEM_stage_inst_dmem_ram_912, MEM_stage_inst_dmem_ram_913, MEM_stage_inst_dmem_ram_914, MEM_stage_inst_dmem_ram_915, MEM_stage_inst_dmem_ram_916, MEM_stage_inst_dmem_ram_917, MEM_stage_inst_dmem_ram_918, MEM_stage_inst_dmem_ram_919, MEM_stage_inst_dmem_ram_920, MEM_stage_inst_dmem_ram_921, MEM_stage_inst_dmem_ram_922, MEM_stage_inst_dmem_ram_923, MEM_stage_inst_dmem_ram_924, MEM_stage_inst_dmem_ram_925, MEM_stage_inst_dmem_ram_926, MEM_stage_inst_dmem_ram_927, MEM_stage_inst_dmem_ram_928, MEM_stage_inst_dmem_ram_929, MEM_stage_inst_dmem_ram_930, MEM_stage_inst_dmem_ram_931, MEM_stage_inst_dmem_ram_932, MEM_stage_inst_dmem_ram_933, MEM_stage_inst_dmem_ram_934, MEM_stage_inst_dmem_ram_935, MEM_stage_inst_dmem_ram_936, MEM_stage_inst_dmem_ram_937, MEM_stage_inst_dmem_ram_938, MEM_stage_inst_dmem_ram_939, MEM_stage_inst_dmem_ram_940, MEM_stage_inst_dmem_ram_941, MEM_stage_inst_dmem_ram_942, MEM_stage_inst_dmem_ram_943, MEM_stage_inst_dmem_ram_944, MEM_stage_inst_dmem_ram_945, MEM_stage_inst_dmem_ram_946, MEM_stage_inst_dmem_ram_947, MEM_stage_inst_dmem_ram_948, MEM_stage_inst_dmem_ram_949, MEM_stage_inst_dmem_ram_950, MEM_stage_inst_dmem_ram_951, MEM_stage_inst_dmem_ram_952, MEM_stage_inst_dmem_ram_953, MEM_stage_inst_dmem_ram_954, MEM_stage_inst_dmem_ram_955, MEM_stage_inst_dmem_ram_956, MEM_stage_inst_dmem_ram_957, MEM_stage_inst_dmem_ram_958, MEM_stage_inst_dmem_ram_959, MEM_stage_inst_dmem_ram_960, MEM_stage_inst_dmem_ram_961, MEM_stage_inst_dmem_ram_962, MEM_stage_inst_dmem_ram_963, MEM_stage_inst_dmem_ram_964, MEM_stage_inst_dmem_ram_965, MEM_stage_inst_dmem_ram_966, MEM_stage_inst_dmem_ram_967, MEM_stage_inst_dmem_ram_968, MEM_stage_inst_dmem_ram_969, MEM_stage_inst_dmem_ram_970, MEM_stage_inst_dmem_ram_971, MEM_stage_inst_dmem_ram_972, MEM_stage_inst_dmem_ram_973, MEM_stage_inst_dmem_ram_974, MEM_stage_inst_dmem_ram_975, MEM_stage_inst_dmem_ram_976, MEM_stage_inst_dmem_ram_977, MEM_stage_inst_dmem_ram_978, MEM_stage_inst_dmem_ram_979, MEM_stage_inst_dmem_ram_980, MEM_stage_inst_dmem_ram_981, MEM_stage_inst_dmem_ram_982, MEM_stage_inst_dmem_ram_983, MEM_stage_inst_dmem_ram_984, MEM_stage_inst_dmem_ram_985, MEM_stage_inst_dmem_ram_986, MEM_stage_inst_dmem_ram_987, MEM_stage_inst_dmem_ram_988, MEM_stage_inst_dmem_ram_989, MEM_stage_inst_dmem_ram_990, MEM_stage_inst_dmem_ram_991, MEM_stage_inst_dmem_ram_992, MEM_stage_inst_dmem_ram_993, MEM_stage_inst_dmem_ram_994, MEM_stage_inst_dmem_ram_995, MEM_stage_inst_dmem_ram_996, MEM_stage_inst_dmem_ram_997, MEM_stage_inst_dmem_ram_998, MEM_stage_inst_dmem_ram_999, MEM_stage_inst_dmem_ram_1000, MEM_stage_inst_dmem_ram_1001, MEM_stage_inst_dmem_ram_1002, MEM_stage_inst_dmem_ram_1003, MEM_stage_inst_dmem_ram_1004, MEM_stage_inst_dmem_ram_1005, MEM_stage_inst_dmem_ram_1006, MEM_stage_inst_dmem_ram_1007, MEM_stage_inst_dmem_ram_1008, MEM_stage_inst_dmem_ram_1009, MEM_stage_inst_dmem_ram_1010, MEM_stage_inst_dmem_ram_1011, MEM_stage_inst_dmem_ram_1012, MEM_stage_inst_dmem_ram_1013, MEM_stage_inst_dmem_ram_1014, MEM_stage_inst_dmem_ram_1015, MEM_stage_inst_dmem_ram_1016, MEM_stage_inst_dmem_ram_1017, MEM_stage_inst_dmem_ram_1018, MEM_stage_inst_dmem_ram_1019, MEM_stage_inst_dmem_ram_1020, MEM_stage_inst_dmem_ram_1021, MEM_stage_inst_dmem_ram_1022, MEM_stage_inst_dmem_ram_1023, MEM_stage_inst_dmem_ram_1, MEM_stage_inst_dmem_ram_2, MEM_stage_inst_dmem_ram_3, MEM_stage_inst_dmem_ram_4, MEM_stage_inst_dmem_ram_5, MEM_stage_inst_dmem_ram_6, MEM_stage_inst_dmem_ram_7, MEM_stage_inst_dmem_ram_8, MEM_stage_inst_dmem_ram_9, MEM_stage_inst_dmem_ram_10, MEM_stage_inst_dmem_ram_11, MEM_stage_inst_dmem_ram_12, MEM_stage_inst_dmem_ram_13, MEM_stage_inst_dmem_ram_14, MEM_stage_inst_dmem_ram_15, MEM_stage_inst_dmem_ram_16, MEM_stage_inst_dmem_ram_17, MEM_stage_inst_dmem_ram_18, MEM_stage_inst_dmem_ram_19, MEM_stage_inst_dmem_ram_20, MEM_stage_inst_dmem_ram_21, MEM_stage_inst_dmem_ram_22, MEM_stage_inst_dmem_ram_23, MEM_stage_inst_dmem_ram_24, MEM_stage_inst_dmem_ram_25, MEM_stage_inst_dmem_ram_26, MEM_stage_inst_dmem_ram_27, MEM_stage_inst_dmem_ram_28, MEM_stage_inst_dmem_ram_29, MEM_stage_inst_dmem_ram_30, MEM_stage_inst_dmem_ram_31, MEM_stage_inst_dmem_ram_32, MEM_stage_inst_dmem_ram_33, MEM_stage_inst_dmem_ram_34, MEM_stage_inst_dmem_ram_35, MEM_stage_inst_dmem_ram_36, MEM_stage_inst_dmem_ram_37, MEM_stage_inst_dmem_ram_38, MEM_stage_inst_dmem_ram_39, MEM_stage_inst_dmem_ram_40, MEM_stage_inst_dmem_ram_41, MEM_stage_inst_dmem_ram_42, MEM_stage_inst_dmem_ram_43, MEM_stage_inst_dmem_ram_44, MEM_stage_inst_dmem_ram_45, MEM_stage_inst_dmem_ram_46, MEM_stage_inst_dmem_ram_47, MEM_stage_inst_dmem_ram_48, MEM_stage_inst_dmem_ram_49, MEM_stage_inst_dmem_ram_50, MEM_stage_inst_dmem_ram_51, MEM_stage_inst_dmem_ram_52, MEM_stage_inst_dmem_ram_53, MEM_stage_inst_dmem_ram_54, MEM_stage_inst_dmem_ram_55, MEM_stage_inst_dmem_ram_56, MEM_stage_inst_dmem_ram_57, MEM_stage_inst_dmem_ram_58, MEM_stage_inst_dmem_ram_59, MEM_stage_inst_dmem_ram_60, MEM_stage_inst_dmem_ram_61, MEM_stage_inst_dmem_ram_62, MEM_stage_inst_dmem_ram_63, MEM_stage_inst_dmem_ram_64, MEM_stage_inst_dmem_ram_65, MEM_stage_inst_dmem_ram_66, MEM_stage_inst_dmem_ram_67, MEM_stage_inst_dmem_ram_68, MEM_stage_inst_dmem_ram_69, MEM_stage_inst_dmem_ram_70, MEM_stage_inst_dmem_ram_71, MEM_stage_inst_dmem_ram_72, MEM_stage_inst_dmem_ram_73, MEM_stage_inst_dmem_ram_74, MEM_stage_inst_dmem_ram_75, MEM_stage_inst_dmem_ram_76, MEM_stage_inst_dmem_ram_77, MEM_stage_inst_dmem_ram_78, MEM_stage_inst_dmem_ram_79, MEM_stage_inst_dmem_ram_80, MEM_stage_inst_dmem_ram_81, MEM_stage_inst_dmem_ram_82, MEM_stage_inst_dmem_ram_83, MEM_stage_inst_dmem_ram_84, MEM_stage_inst_dmem_ram_85, MEM_stage_inst_dmem_ram_86, MEM_stage_inst_dmem_ram_87, MEM_stage_inst_dmem_ram_88, MEM_stage_inst_dmem_ram_89, MEM_stage_inst_dmem_ram_90, MEM_stage_inst_dmem_ram_91, MEM_stage_inst_dmem_ram_92, MEM_stage_inst_dmem_ram_93, MEM_stage_inst_dmem_ram_94, MEM_stage_inst_dmem_ram_95, MEM_stage_inst_dmem_ram_96, MEM_stage_inst_dmem_ram_97, MEM_stage_inst_dmem_ram_98, MEM_stage_inst_dmem_ram_99, MEM_stage_inst_dmem_ram_100, MEM_stage_inst_dmem_ram_101, MEM_stage_inst_dmem_ram_102, MEM_stage_inst_dmem_ram_103, MEM_stage_inst_dmem_ram_104, MEM_stage_inst_dmem_ram_105, MEM_stage_inst_dmem_ram_106, MEM_stage_inst_dmem_ram_107, MEM_stage_inst_dmem_ram_108, MEM_stage_inst_dmem_ram_109, MEM_stage_inst_dmem_ram_110, MEM_stage_inst_dmem_ram_111, MEM_stage_inst_dmem_ram_112, MEM_stage_inst_dmem_ram_113, MEM_stage_inst_dmem_ram_114, MEM_stage_inst_dmem_ram_115, MEM_stage_inst_dmem_ram_116, MEM_stage_inst_dmem_ram_117, MEM_stage_inst_dmem_ram_118, MEM_stage_inst_dmem_ram_119, MEM_stage_inst_dmem_ram_120, MEM_stage_inst_dmem_ram_121, MEM_stage_inst_dmem_ram_122, MEM_stage_inst_dmem_ram_123, MEM_stage_inst_dmem_ram_124, MEM_stage_inst_dmem_ram_125, MEM_stage_inst_dmem_ram_126, MEM_stage_inst_dmem_ram_127, MEM_stage_inst_dmem_ram_128, MEM_stage_inst_dmem_ram_129, MEM_stage_inst_dmem_ram_130, MEM_stage_inst_dmem_ram_131, MEM_stage_inst_dmem_ram_132, MEM_stage_inst_dmem_ram_133, MEM_stage_inst_dmem_ram_134, MEM_stage_inst_dmem_ram_135, MEM_stage_inst_dmem_ram_136, MEM_stage_inst_dmem_ram_137, MEM_stage_inst_dmem_ram_138, MEM_stage_inst_dmem_ram_139, MEM_stage_inst_dmem_ram_140, MEM_stage_inst_dmem_ram_141, MEM_stage_inst_dmem_ram_142, MEM_stage_inst_dmem_ram_143, MEM_stage_inst_dmem_ram_144, MEM_stage_inst_dmem_ram_145, MEM_stage_inst_dmem_ram_146, MEM_stage_inst_dmem_ram_147, MEM_stage_inst_dmem_ram_148, MEM_stage_inst_dmem_ram_149, MEM_stage_inst_dmem_ram_150, MEM_stage_inst_dmem_ram_151, MEM_stage_inst_dmem_ram_152, MEM_stage_inst_dmem_ram_153, MEM_stage_inst_dmem_ram_154, MEM_stage_inst_dmem_ram_155, MEM_stage_inst_dmem_ram_156, MEM_stage_inst_dmem_ram_157, MEM_stage_inst_dmem_ram_158, MEM_stage_inst_dmem_ram_159, MEM_stage_inst_dmem_ram_160, MEM_stage_inst_dmem_ram_161, MEM_stage_inst_dmem_ram_162, MEM_stage_inst_dmem_ram_163, MEM_stage_inst_dmem_ram_164, MEM_stage_inst_dmem_ram_165, MEM_stage_inst_dmem_ram_166, MEM_stage_inst_dmem_ram_167, MEM_stage_inst_dmem_ram_168, MEM_stage_inst_dmem_ram_169, MEM_stage_inst_dmem_ram_170, MEM_stage_inst_dmem_ram_171, MEM_stage_inst_dmem_ram_172, MEM_stage_inst_dmem_ram_173, MEM_stage_inst_dmem_ram_174, MEM_stage_inst_dmem_ram_175, MEM_stage_inst_dmem_ram_176, MEM_stage_inst_dmem_ram_177, MEM_stage_inst_dmem_ram_178, MEM_stage_inst_dmem_ram_179, MEM_stage_inst_dmem_ram_180, MEM_stage_inst_dmem_ram_181, MEM_stage_inst_dmem_ram_182, MEM_stage_inst_dmem_ram_183, MEM_stage_inst_dmem_ram_184, MEM_stage_inst_dmem_ram_185, MEM_stage_inst_dmem_ram_186, MEM_stage_inst_dmem_ram_187, MEM_stage_inst_dmem_ram_188, MEM_stage_inst_dmem_ram_189, MEM_stage_inst_dmem_ram_190, MEM_stage_inst_dmem_ram_191, MEM_stage_inst_dmem_ram_192, MEM_stage_inst_dmem_ram_193, MEM_stage_inst_dmem_ram_194, MEM_stage_inst_dmem_ram_195, MEM_stage_inst_dmem_ram_196, MEM_stage_inst_dmem_ram_197, MEM_stage_inst_dmem_ram_198, MEM_stage_inst_dmem_ram_199, MEM_stage_inst_dmem_ram_200, MEM_stage_inst_dmem_ram_201, MEM_stage_inst_dmem_ram_202, MEM_stage_inst_dmem_ram_203, MEM_stage_inst_dmem_ram_204, MEM_stage_inst_dmem_ram_205, MEM_stage_inst_dmem_ram_206, MEM_stage_inst_dmem_ram_207, MEM_stage_inst_dmem_ram_208, MEM_stage_inst_dmem_ram_209, MEM_stage_inst_dmem_ram_210, MEM_stage_inst_dmem_ram_211, MEM_stage_inst_dmem_ram_212, MEM_stage_inst_dmem_ram_213, MEM_stage_inst_dmem_ram_214, MEM_stage_inst_dmem_ram_215, MEM_stage_inst_dmem_ram_216, MEM_stage_inst_dmem_ram_217, MEM_stage_inst_dmem_ram_218, MEM_stage_inst_dmem_ram_219, MEM_stage_inst_dmem_ram_220, MEM_stage_inst_dmem_ram_221, MEM_stage_inst_dmem_ram_222, MEM_stage_inst_dmem_ram_223, MEM_stage_inst_dmem_ram_224, MEM_stage_inst_dmem_ram_225, MEM_stage_inst_dmem_ram_226, MEM_stage_inst_dmem_ram_227, MEM_stage_inst_dmem_ram_228, MEM_stage_inst_dmem_ram_229, MEM_stage_inst_dmem_ram_230, MEM_stage_inst_dmem_ram_231, MEM_stage_inst_dmem_ram_232, MEM_stage_inst_dmem_ram_233, MEM_stage_inst_dmem_ram_234, MEM_stage_inst_dmem_ram_235, MEM_stage_inst_dmem_ram_236, MEM_stage_inst_dmem_ram_237, MEM_stage_inst_dmem_ram_238, MEM_stage_inst_dmem_ram_239, MEM_stage_inst_dmem_ram_240, MEM_stage_inst_dmem_ram_241, MEM_stage_inst_dmem_ram_242, MEM_stage_inst_dmem_ram_243, MEM_stage_inst_dmem_ram_244, MEM_stage_inst_dmem_ram_245, MEM_stage_inst_dmem_ram_246, MEM_stage_inst_dmem_ram_247, MEM_stage_inst_dmem_ram_248, MEM_stage_inst_dmem_ram_249, MEM_stage_inst_dmem_ram_250, MEM_stage_inst_dmem_ram_251, MEM_stage_inst_dmem_ram_252, MEM_stage_inst_dmem_ram_253, MEM_stage_inst_dmem_ram_254, MEM_stage_inst_dmem_ram_255, MEM_stage_inst_dmem_ram_256, MEM_stage_inst_dmem_ram_257, MEM_stage_inst_dmem_ram_258, MEM_stage_inst_dmem_ram_259, MEM_stage_inst_dmem_ram_260, MEM_stage_inst_dmem_ram_261, MEM_stage_inst_dmem_ram_262, MEM_stage_inst_dmem_ram_263, MEM_stage_inst_dmem_ram_264, MEM_stage_inst_dmem_ram_265, MEM_stage_inst_dmem_ram_266, MEM_stage_inst_dmem_ram_267, MEM_stage_inst_dmem_ram_268, MEM_stage_inst_dmem_ram_269, MEM_stage_inst_dmem_ram_270, MEM_stage_inst_dmem_ram_271, MEM_stage_inst_dmem_ram_272, MEM_stage_inst_dmem_ram_273, MEM_stage_inst_dmem_ram_274, MEM_stage_inst_dmem_ram_275, MEM_stage_inst_dmem_ram_276, MEM_stage_inst_dmem_ram_277, MEM_stage_inst_dmem_ram_278, MEM_stage_inst_dmem_ram_279, MEM_stage_inst_dmem_ram_280, MEM_stage_inst_dmem_ram_281, MEM_stage_inst_dmem_ram_282, MEM_stage_inst_dmem_ram_283, MEM_stage_inst_dmem_ram_284, MEM_stage_inst_dmem_ram_285, MEM_stage_inst_dmem_ram_286, MEM_stage_inst_dmem_ram_287, MEM_stage_inst_dmem_ram_288, MEM_stage_inst_dmem_ram_289, MEM_stage_inst_dmem_ram_290, MEM_stage_inst_dmem_ram_291, MEM_stage_inst_dmem_ram_292, MEM_stage_inst_dmem_ram_293, MEM_stage_inst_dmem_ram_294, MEM_stage_inst_dmem_ram_295, MEM_stage_inst_dmem_ram_296, MEM_stage_inst_dmem_ram_297, MEM_stage_inst_dmem_ram_298, MEM_stage_inst_dmem_ram_299, MEM_stage_inst_dmem_ram_300, MEM_stage_inst_dmem_ram_301, MEM_stage_inst_dmem_ram_302, MEM_stage_inst_dmem_ram_303, MEM_stage_inst_dmem_ram_304, MEM_stage_inst_dmem_ram_305, MEM_stage_inst_dmem_ram_306, MEM_stage_inst_dmem_ram_307, MEM_stage_inst_dmem_ram_308, MEM_stage_inst_dmem_ram_309, MEM_stage_inst_dmem_ram_310, MEM_stage_inst_dmem_ram_311, MEM_stage_inst_dmem_ram_312, MEM_stage_inst_dmem_ram_313, MEM_stage_inst_dmem_ram_314, MEM_stage_inst_dmem_ram_315, MEM_stage_inst_dmem_ram_316, MEM_stage_inst_dmem_ram_317, MEM_stage_inst_dmem_ram_318, MEM_stage_inst_dmem_ram_319, MEM_stage_inst_dmem_ram_320, MEM_stage_inst_dmem_ram_321, MEM_stage_inst_dmem_ram_322, MEM_stage_inst_dmem_ram_323, MEM_stage_inst_dmem_ram_324, MEM_stage_inst_dmem_ram_325, MEM_stage_inst_dmem_ram_326, MEM_stage_inst_dmem_ram_327, MEM_stage_inst_dmem_ram_328, MEM_stage_inst_dmem_ram_329, MEM_stage_inst_dmem_ram_330, MEM_stage_inst_dmem_ram_331, MEM_stage_inst_dmem_ram_332, MEM_stage_inst_dmem_ram_333, MEM_stage_inst_dmem_ram_334, MEM_stage_inst_dmem_ram_335, MEM_stage_inst_dmem_ram_336, MEM_stage_inst_dmem_ram_337, MEM_stage_inst_dmem_ram_338, MEM_stage_inst_dmem_ram_339, MEM_stage_inst_dmem_ram_340, MEM_stage_inst_dmem_ram_341, MEM_stage_inst_dmem_ram_342, MEM_stage_inst_dmem_ram_343, MEM_stage_inst_dmem_ram_344, MEM_stage_inst_dmem_ram_345, MEM_stage_inst_dmem_ram_346, MEM_stage_inst_dmem_ram_347, MEM_stage_inst_dmem_ram_348, MEM_stage_inst_dmem_ram_349, MEM_stage_inst_dmem_ram_350, MEM_stage_inst_dmem_ram_351, MEM_stage_inst_dmem_ram_352, MEM_stage_inst_dmem_ram_353, MEM_stage_inst_dmem_ram_354, MEM_stage_inst_dmem_ram_355, MEM_stage_inst_dmem_ram_356, MEM_stage_inst_dmem_ram_357, MEM_stage_inst_dmem_ram_358, MEM_stage_inst_dmem_ram_359, MEM_stage_inst_dmem_ram_360, MEM_stage_inst_dmem_ram_361, MEM_stage_inst_dmem_ram_362, MEM_stage_inst_dmem_ram_363, MEM_stage_inst_dmem_ram_364, MEM_stage_inst_dmem_ram_365, MEM_stage_inst_dmem_ram_366, MEM_stage_inst_dmem_ram_367, MEM_stage_inst_dmem_ram_368, MEM_stage_inst_dmem_ram_369, MEM_stage_inst_dmem_ram_370, MEM_stage_inst_dmem_ram_371, MEM_stage_inst_dmem_ram_372, MEM_stage_inst_dmem_ram_373, MEM_stage_inst_dmem_ram_374, MEM_stage_inst_dmem_ram_375, MEM_stage_inst_dmem_ram_376, MEM_stage_inst_dmem_ram_377, MEM_stage_inst_dmem_ram_378, MEM_stage_inst_dmem_ram_379, MEM_stage_inst_dmem_ram_380, MEM_stage_inst_dmem_ram_381, MEM_stage_inst_dmem_ram_382, MEM_stage_inst_dmem_ram_383, MEM_stage_inst_dmem_ram_384, MEM_stage_inst_dmem_ram_385, MEM_stage_inst_dmem_ram_386, MEM_stage_inst_dmem_ram_387, MEM_stage_inst_dmem_ram_388, MEM_stage_inst_dmem_ram_389, MEM_stage_inst_dmem_ram_390, MEM_stage_inst_dmem_ram_391, MEM_stage_inst_dmem_ram_392, MEM_stage_inst_dmem_ram_393, MEM_stage_inst_dmem_ram_394, MEM_stage_inst_dmem_ram_395, MEM_stage_inst_dmem_ram_396, MEM_stage_inst_dmem_ram_397, MEM_stage_inst_dmem_ram_398, MEM_stage_inst_dmem_ram_399, MEM_stage_inst_dmem_ram_400, MEM_stage_inst_dmem_ram_401, MEM_stage_inst_dmem_ram_402, MEM_stage_inst_dmem_ram_403, MEM_stage_inst_dmem_ram_404, MEM_stage_inst_dmem_ram_405, MEM_stage_inst_dmem_ram_406, MEM_stage_inst_dmem_ram_407, MEM_stage_inst_dmem_ram_408, MEM_stage_inst_dmem_ram_409, MEM_stage_inst_dmem_ram_410, MEM_stage_inst_dmem_ram_411, MEM_stage_inst_dmem_ram_412, MEM_stage_inst_dmem_ram_413, MEM_stage_inst_dmem_ram_414, MEM_stage_inst_dmem_ram_415, MEM_stage_inst_dmem_ram_416, MEM_stage_inst_dmem_ram_417, MEM_stage_inst_dmem_ram_418, MEM_stage_inst_dmem_ram_419, MEM_stage_inst_dmem_ram_420, MEM_stage_inst_dmem_ram_421, MEM_stage_inst_dmem_ram_422, MEM_stage_inst_dmem_ram_423, MEM_stage_inst_dmem_ram_424, MEM_stage_inst_dmem_ram_425, MEM_stage_inst_dmem_ram_426, MEM_stage_inst_dmem_ram_427, MEM_stage_inst_dmem_ram_428, MEM_stage_inst_dmem_ram_429, MEM_stage_inst_dmem_ram_430, MEM_stage_inst_dmem_ram_431, MEM_stage_inst_dmem_ram_432, MEM_stage_inst_dmem_ram_433, MEM_stage_inst_dmem_ram_434, MEM_stage_inst_dmem_ram_435, MEM_stage_inst_dmem_ram_436, MEM_stage_inst_dmem_ram_437, MEM_stage_inst_dmem_ram_438, MEM_stage_inst_dmem_ram_439, MEM_stage_inst_dmem_ram_440, MEM_stage_inst_dmem_ram_441, MEM_stage_inst_dmem_ram_442, MEM_stage_inst_dmem_ram_443, MEM_stage_inst_dmem_ram_444, MEM_stage_inst_dmem_ram_445, MEM_stage_inst_dmem_ram_446, MEM_stage_inst_dmem_ram_447, MEM_stage_inst_dmem_ram_448, MEM_stage_inst_dmem_ram_449, MEM_stage_inst_dmem_ram_450, MEM_stage_inst_dmem_ram_451, MEM_stage_inst_dmem_ram_452, MEM_stage_inst_dmem_ram_453, MEM_stage_inst_dmem_ram_454, MEM_stage_inst_dmem_ram_455, MEM_stage_inst_dmem_ram_456, MEM_stage_inst_dmem_ram_457, MEM_stage_inst_dmem_ram_458, MEM_stage_inst_dmem_ram_459, MEM_stage_inst_dmem_ram_460, MEM_stage_inst_dmem_ram_461, MEM_stage_inst_dmem_ram_462, MEM_stage_inst_dmem_ram_463, MEM_stage_inst_dmem_ram_464, MEM_stage_inst_dmem_ram_465, MEM_stage_inst_dmem_ram_466, MEM_stage_inst_dmem_ram_467, MEM_stage_inst_dmem_ram_468, MEM_stage_inst_dmem_ram_469, MEM_stage_inst_dmem_ram_470, MEM_stage_inst_dmem_ram_471, MEM_stage_inst_dmem_ram_472, MEM_stage_inst_dmem_ram_473, MEM_stage_inst_dmem_ram_474, MEM_stage_inst_dmem_ram_475, MEM_stage_inst_dmem_ram_476, MEM_stage_inst_dmem_ram_477, MEM_stage_inst_dmem_ram_478, MEM_stage_inst_dmem_ram_479, MEM_stage_inst_dmem_ram_480, MEM_stage_inst_dmem_ram_481, MEM_stage_inst_dmem_ram_482, MEM_stage_inst_dmem_ram_483, MEM_stage_inst_dmem_ram_484, MEM_stage_inst_dmem_ram_485, MEM_stage_inst_dmem_ram_486, MEM_stage_inst_dmem_ram_487, MEM_stage_inst_dmem_ram_488, MEM_stage_inst_dmem_ram_489, MEM_stage_inst_dmem_ram_490, MEM_stage_inst_dmem_ram_491, MEM_stage_inst_dmem_ram_492, MEM_stage_inst_dmem_ram_493, MEM_stage_inst_dmem_ram_494, MEM_stage_inst_dmem_ram_495, MEM_stage_inst_dmem_ram_496, MEM_stage_inst_dmem_ram_497, MEM_stage_inst_dmem_ram_498, MEM_stage_inst_dmem_ram_499, MEM_stage_inst_dmem_ram_500, MEM_stage_inst_dmem_ram_501, MEM_stage_inst_dmem_ram_502, MEM_stage_inst_dmem_ram_503, MEM_stage_inst_dmem_ram_504, MEM_stage_inst_dmem_ram_505, MEM_stage_inst_dmem_ram_506, MEM_stage_inst_dmem_ram_507, MEM_stage_inst_dmem_ram_508, MEM_stage_inst_dmem_ram_509, MEM_stage_inst_dmem_ram_510, MEM_stage_inst_dmem_ram_511, MEM_stage_inst_dmem_ram_0, pc_7_, pc_6_, pc_5_, pc_4_, pc_3_, pc_2_, pc_1_, pc_0_ ;
output MEM_stage_inst_N6, EX_stage_inst_N4, MEM_stage_inst_N4, EX_stage_inst_N5, MEM_stage_inst_N5, EX_stage_inst_N6, EX_stage_inst_N3, EX_stage_inst_N7, EX_stage_inst_N24, MEM_stage_inst_N7, EX_stage_inst_N40, MEM_stage_inst_N39, EX_stage_inst_N23, EX_stage_inst_N25, MEM_stage_inst_N24, EX_stage_inst_N8, EX_stage_inst_N33, MEM_stage_inst_N32, EX_stage_inst_N16, EX_stage_inst_N35, MEM_stage_inst_N34, EX_stage_inst_N18, EX_stage_inst_N37, MEM_stage_inst_N36, EX_stage_inst_N20, EX_stage_inst_N39, MEM_stage_inst_N38, EX_stage_inst_N22, EX_stage_inst_N29, MEM_stage_inst_N28, EX_stage_inst_N12, EX_stage_inst_N31, MEM_stage_inst_N30, EX_stage_inst_N14, EX_stage_inst_N36, MEM_stage_inst_N35, EX_stage_inst_N19, EX_stage_inst_N38, MEM_stage_inst_N37, EX_stage_inst_N21, EX_stage_inst_N27, MEM_stage_inst_N26, EX_stage_inst_N10, EX_stage_inst_N28, MEM_stage_inst_N27, EX_stage_inst_N11, EX_stage_inst_N26, MEM_stage_inst_N25, EX_stage_inst_N9, EX_stage_inst_N30, MEM_stage_inst_N29, EX_stage_inst_N13, EX_stage_inst_N34, MEM_stage_inst_N33, EX_stage_inst_N17, EX_stage_inst_N32, MEM_stage_inst_N31, EX_stage_inst_N15, MEM_stage_inst_N8, MEM_stage_inst_N9, MEM_stage_inst_N10, MEM_stage_inst_N11, MEM_stage_inst_N12, MEM_stage_inst_N13, MEM_stage_inst_N14, MEM_stage_inst_N15, MEM_stage_inst_N16, MEM_stage_inst_N17, MEM_stage_inst_N18, MEM_stage_inst_N19, MEM_stage_inst_N20, MEM_stage_inst_N21, MEM_stage_inst_N22, MEM_stage_inst_N23, n1734, n3520, n1731, n3517, n1730, n1741, n1729, n1739, n1728, n1727, n1724, n3521, n1722, n3518, n1725, n1723, n1713, n1714, n1726, n1721, n1720, n1719, n1718, ID_stage_inst_ir_dest_with_bubble_0, n1717, ID_stage_inst_ir_dest_with_bubble_1, n1716, ID_stage_inst_ir_dest_with_bubble_2, n1715, n1712, ID_stage_inst_ex_alu_cmd_1, ID_stage_inst_ex_alu_cmd_0, ID_stage_inst_ex_alu_cmd_2, ID_stage_inst_write_back_result_mux, ID_stage_inst_write_back_en, n1738, n1735, reg_read_data_1_15, n1606, n1605, n3519, n1604, n1603, n1602, n1601, reg_read_data_2_15, ID_stage_inst_ex_alu_src2_15, n1711, n1710, n1709, n1708, n1707, n1706, n1705, reg_read_data_2_0, reg_read_data_1_0, n1655, n1654, n1653, n1652, n1651, n1650, n1649, reg_read_data_2_8, ID_stage_inst_ex_alu_src2_8, reg_read_data_1_8, n1641, n1640, n1639, n1638, n1637, n1636, n1635, reg_read_data_2_10, ID_stage_inst_ex_alu_src2_10, reg_read_data_1_10, n1627, n1626, n1625, n1624, n1623, n1622, n1621, reg_read_data_2_12, ID_stage_inst_ex_alu_src2_12, reg_read_data_1_12, n1613, n1612, n1611, n1610, n1609, n1608, n1607, reg_read_data_2_14, ID_stage_inst_ex_alu_src2_14, reg_read_data_1_14, n1683, n1682, n1681, n1680, n1679, n1678, n1677, reg_read_data_2_4, ID_stage_inst_ex_alu_src2_4, reg_read_data_1_4, n1669, n1668, n1667, n1666, n1665, n1664, n1663, reg_read_data_2_6, ID_stage_inst_ex_alu_src2_6, reg_read_data_1_6, n1634, n1633, n1632, n1631, n1630, n1629, n1628, reg_read_data_2_11, ID_stage_inst_ex_alu_src2_11, reg_read_data_1_11, n1620, n1619, n1618, n1617, n1616, n1615, n1614, reg_read_data_2_13, ID_stage_inst_ex_alu_src2_13, reg_read_data_1_13, n1697, n1696, n1695, n1694, n1693, n1692, n1691, reg_read_data_2_2, reg_read_data_1_2, n1690, n1689, n1688, n1687, n1686, n1685, n1684, reg_read_data_2_3, reg_read_data_1_3, n1704, n1703, n1702, n1701, n1700, n1699, n1698, reg_read_data_2_1, reg_read_data_1_1, n1676, n1675, n1674, n1673, n1672, n1671, n1670, reg_read_data_2_5, ID_stage_inst_ex_alu_src2_5, reg_read_data_1_5, n1648, n1647, n1646, n1645, n1644, n1643, n1642, reg_read_data_2_9, ID_stage_inst_ex_alu_src2_9, reg_read_data_1_9, n1662, n1661, n1660, n1659, n1658, n1657, n1656, reg_read_data_2_7, ID_stage_inst_ex_alu_src2_7, reg_read_data_1_7, n1732, ID_stage_inst_ex_alu_src2_1, MEM_stage_inst_N3, ID_stage_inst_ex_alu_src2_2, ID_stage_inst_ex_alu_src2_0, ID_stage_inst_ex_alu_src2_3, n1733, MEM_stage_inst_dmem_n8763, MEM_stage_inst_dmem_n21529, MEM_stage_inst_dmem_n8764, MEM_stage_inst_dmem_n21573, MEM_stage_inst_dmem_n8765, MEM_stage_inst_dmem_n21564, MEM_stage_inst_dmem_n8766, MEM_stage_inst_dmem_n21580, MEM_stage_inst_dmem_n8767, MEM_stage_inst_dmem_n21538, MEM_stage_inst_dmem_n8768, MEM_stage_inst_dmem_n21540, MEM_stage_inst_dmem_n8769, MEM_stage_inst_dmem_n21605, MEM_stage_inst_dmem_n8770, MEM_stage_inst_dmem_n21579, MEM_stage_inst_dmem_n8771, MEM_stage_inst_dmem_n21575, MEM_stage_inst_dmem_n8772, MEM_stage_inst_dmem_n21584, MEM_stage_inst_dmem_n8773, MEM_stage_inst_dmem_n21597, MEM_stage_inst_dmem_n8774, MEM_stage_inst_dmem_n21542, MEM_stage_inst_dmem_n8775, MEM_stage_inst_dmem_n21586, MEM_stage_inst_dmem_n8776, MEM_stage_inst_dmem_n21570, MEM_stage_inst_dmem_n8777, MEM_stage_inst_dmem_n21546, MEM_stage_inst_dmem_n8778, MEM_stage_inst_dmem_n21532, MEM_stage_inst_dmem_n8779, MEM_stage_inst_dmem_n21549, MEM_stage_inst_dmem_n8780, MEM_stage_inst_dmem_n21553, MEM_stage_inst_dmem_n8781, MEM_stage_inst_dmem_n21629, MEM_stage_inst_dmem_n8782, MEM_stage_inst_dmem_n21547, MEM_stage_inst_dmem_n8783, MEM_stage_inst_dmem_n21572, MEM_stage_inst_dmem_n8784, MEM_stage_inst_dmem_n21559, MEM_stage_inst_dmem_n8785, MEM_stage_inst_dmem_n21600, MEM_stage_inst_dmem_n8786, MEM_stage_inst_dmem_n21554, MEM_stage_inst_dmem_n8787, MEM_stage_inst_dmem_n8788, MEM_stage_inst_dmem_n8789, MEM_stage_inst_dmem_n8790, MEM_stage_inst_dmem_n21591, MEM_stage_inst_dmem_n8791, MEM_stage_inst_dmem_n21527, MEM_stage_inst_dmem_n8792, MEM_stage_inst_dmem_n21622, MEM_stage_inst_dmem_n8793, MEM_stage_inst_dmem_n8794, MEM_stage_inst_dmem_n21590, MEM_stage_inst_dmem_n8795, MEM_stage_inst_dmem_n21610, MEM_stage_inst_dmem_n8796, MEM_stage_inst_dmem_n21612, MEM_stage_inst_dmem_n8797, MEM_stage_inst_dmem_n21616, MEM_stage_inst_dmem_n8798, MEM_stage_inst_dmem_n21582, MEM_stage_inst_dmem_n8799, MEM_stage_inst_dmem_n21537, MEM_stage_inst_dmem_n8800, MEM_stage_inst_dmem_n21602, MEM_stage_inst_dmem_n8801, MEM_stage_inst_dmem_n21574, MEM_stage_inst_dmem_n8802, MEM_stage_inst_dmem_n21566, MEM_stage_inst_dmem_n8803, MEM_stage_inst_dmem_n8804, MEM_stage_inst_dmem_n21543, MEM_stage_inst_dmem_n8805, MEM_stage_inst_dmem_n8806, MEM_stage_inst_dmem_n8807, MEM_stage_inst_dmem_n8808, MEM_stage_inst_dmem_n8809, MEM_stage_inst_dmem_n8810, MEM_stage_inst_dmem_n8811, MEM_stage_inst_dmem_n21619, MEM_stage_inst_dmem_n8812, MEM_stage_inst_dmem_n21525, MEM_stage_inst_dmem_n8813, MEM_stage_inst_dmem_n21593, MEM_stage_inst_dmem_n8814, MEM_stage_inst_dmem_n8815, MEM_stage_inst_dmem_n21524, MEM_stage_inst_dmem_n8816, MEM_stage_inst_dmem_n21511, MEM_stage_inst_dmem_n8817, MEM_stage_inst_dmem_n21556, MEM_stage_inst_dmem_n8818, MEM_stage_inst_dmem_n8819, MEM_stage_inst_dmem_n21576, MEM_stage_inst_dmem_n8820, MEM_stage_inst_dmem_n8821, MEM_stage_inst_dmem_n8822, MEM_stage_inst_dmem_n21544, MEM_stage_inst_dmem_n8823, MEM_stage_inst_dmem_n8824, MEM_stage_inst_dmem_n21519, MEM_stage_inst_dmem_n8825, MEM_stage_inst_dmem_n21510, MEM_stage_inst_dmem_n8826, MEM_stage_inst_dmem_n8827, MEM_stage_inst_dmem_n21569, MEM_stage_inst_dmem_n8828, MEM_stage_inst_dmem_n21625, MEM_stage_inst_dmem_n8829, MEM_stage_inst_dmem_n21608, MEM_stage_inst_dmem_n8830, MEM_stage_inst_dmem_n21563, MEM_stage_inst_dmem_n8831, MEM_stage_inst_dmem_n21526, MEM_stage_inst_dmem_n8832, MEM_stage_inst_dmem_n21588, MEM_stage_inst_dmem_n8833, MEM_stage_inst_dmem_n21618, MEM_stage_inst_dmem_n8834, MEM_stage_inst_dmem_n21624, MEM_stage_inst_dmem_n8835, MEM_stage_inst_dmem_n21522, MEM_stage_inst_dmem_n8836, MEM_stage_inst_dmem_n21615, MEM_stage_inst_dmem_n8837, MEM_stage_inst_dmem_n21617, MEM_stage_inst_dmem_n8838, MEM_stage_inst_dmem_n8839, MEM_stage_inst_dmem_n21555, MEM_stage_inst_dmem_n8840, MEM_stage_inst_dmem_n21606, MEM_stage_inst_dmem_n8841, MEM_stage_inst_dmem_n21539, MEM_stage_inst_dmem_n8842, MEM_stage_inst_dmem_n21568, MEM_stage_inst_dmem_n8843, MEM_stage_inst_dmem_n8844, MEM_stage_inst_dmem_n8845, MEM_stage_inst_dmem_n8846, MEM_stage_inst_dmem_n21594, MEM_stage_inst_dmem_n8847, MEM_stage_inst_dmem_n21548, MEM_stage_inst_dmem_n8848, MEM_stage_inst_dmem_n21565, MEM_stage_inst_dmem_n8849, MEM_stage_inst_dmem_n8850, MEM_stage_inst_dmem_n8851, MEM_stage_inst_dmem_n21534, MEM_stage_inst_dmem_n8852, MEM_stage_inst_dmem_n8853, MEM_stage_inst_dmem_n21609, MEM_stage_inst_dmem_n8854, MEM_stage_inst_dmem_n8855, MEM_stage_inst_dmem_n21621, MEM_stage_inst_dmem_n8856, MEM_stage_inst_dmem_n8857, MEM_stage_inst_dmem_n21633, MEM_stage_inst_dmem_n8858, MEM_stage_inst_dmem_n21604, MEM_stage_inst_dmem_n8859, MEM_stage_inst_dmem_n21518, MEM_stage_inst_dmem_n8860, MEM_stage_inst_dmem_n8861, MEM_stage_inst_dmem_n8862, MEM_stage_inst_dmem_n8863, MEM_stage_inst_dmem_n21636, MEM_stage_inst_dmem_n8864, MEM_stage_inst_dmem_n8865, MEM_stage_inst_dmem_n8866, MEM_stage_inst_dmem_n8867, MEM_stage_inst_dmem_n21589, MEM_stage_inst_dmem_n8868, MEM_stage_inst_dmem_n8869, MEM_stage_inst_dmem_n8870, MEM_stage_inst_dmem_n8871, MEM_stage_inst_dmem_n8872, MEM_stage_inst_dmem_n8873, MEM_stage_inst_dmem_n8874, MEM_stage_inst_dmem_n21514, MEM_stage_inst_dmem_n8875, MEM_stage_inst_dmem_n21592, MEM_stage_inst_dmem_n8876, MEM_stage_inst_dmem_n21628, MEM_stage_inst_dmem_n8877, MEM_stage_inst_dmem_n21513, MEM_stage_inst_dmem_n8878, MEM_stage_inst_dmem_n8879, MEM_stage_inst_dmem_n21623, MEM_stage_inst_dmem_n8880, MEM_stage_inst_dmem_n21583, MEM_stage_inst_dmem_n8881, MEM_stage_inst_dmem_n21613, MEM_stage_inst_dmem_n8882, MEM_stage_inst_dmem_n8883, MEM_stage_inst_dmem_n21516, MEM_stage_inst_dmem_n8884, MEM_stage_inst_dmem_n8885, MEM_stage_inst_dmem_n21509, MEM_stage_inst_dmem_n8886, MEM_stage_inst_dmem_n8887, MEM_stage_inst_dmem_n21558, MEM_stage_inst_dmem_n8888, MEM_stage_inst_dmem_n8889, MEM_stage_inst_dmem_n8890, MEM_stage_inst_dmem_n8891, MEM_stage_inst_dmem_n8892, MEM_stage_inst_dmem_n8893, MEM_stage_inst_dmem_n8894, MEM_stage_inst_dmem_n8895, MEM_stage_inst_dmem_n8896, MEM_stage_inst_dmem_n21587, MEM_stage_inst_dmem_n8897, MEM_stage_inst_dmem_n8898, MEM_stage_inst_dmem_n21626, MEM_stage_inst_dmem_n8899, MEM_stage_inst_dmem_n21599, MEM_stage_inst_dmem_n8900, MEM_stage_inst_dmem_n8901, MEM_stage_inst_dmem_n21598, MEM_stage_inst_dmem_n8902, MEM_stage_inst_dmem_n21552, MEM_stage_inst_dmem_n8903, MEM_stage_inst_dmem_n8904, MEM_stage_inst_dmem_n8905, MEM_stage_inst_dmem_n21523, MEM_stage_inst_dmem_n8906, MEM_stage_inst_dmem_n21517, MEM_stage_inst_dmem_n8907, MEM_stage_inst_dmem_n21601, MEM_stage_inst_dmem_n8908, MEM_stage_inst_dmem_n21603, MEM_stage_inst_dmem_n8909, MEM_stage_inst_dmem_n8910, MEM_stage_inst_dmem_n8911, MEM_stage_inst_dmem_n8912, MEM_stage_inst_dmem_n21515, MEM_stage_inst_dmem_n8913, MEM_stage_inst_dmem_n8914, MEM_stage_inst_dmem_n21578, MEM_stage_inst_dmem_n8915, MEM_stage_inst_dmem_n8916, MEM_stage_inst_dmem_n8917, MEM_stage_inst_dmem_n8918, MEM_stage_inst_dmem_n8919, MEM_stage_inst_dmem_n8920, MEM_stage_inst_dmem_n8921, MEM_stage_inst_dmem_n8922, MEM_stage_inst_dmem_n21551, MEM_stage_inst_dmem_n8923, MEM_stage_inst_dmem_n8924, MEM_stage_inst_dmem_n21620, MEM_stage_inst_dmem_n8925, MEM_stage_inst_dmem_n8926, MEM_stage_inst_dmem_n8927, MEM_stage_inst_dmem_n8928, MEM_stage_inst_dmem_n8929, MEM_stage_inst_dmem_n8930, MEM_stage_inst_dmem_n8931, MEM_stage_inst_dmem_n8932, MEM_stage_inst_dmem_n21596, MEM_stage_inst_dmem_n8933, MEM_stage_inst_dmem_n8934, MEM_stage_inst_dmem_n8935, MEM_stage_inst_dmem_n8936, MEM_stage_inst_dmem_n8937, MEM_stage_inst_dmem_n21550, MEM_stage_inst_dmem_n8938, MEM_stage_inst_dmem_n8939, MEM_stage_inst_dmem_n8940, MEM_stage_inst_dmem_n21632, MEM_stage_inst_dmem_n8941, MEM_stage_inst_dmem_n21635, MEM_stage_inst_dmem_n8942, MEM_stage_inst_dmem_n8943, MEM_stage_inst_dmem_n8944, MEM_stage_inst_dmem_n8945, MEM_stage_inst_dmem_n8946, MEM_stage_inst_dmem_n8947, MEM_stage_inst_dmem_n8948, MEM_stage_inst_dmem_n8949, MEM_stage_inst_dmem_n8950, MEM_stage_inst_dmem_n8951, MEM_stage_inst_dmem_n21611, MEM_stage_inst_dmem_n8952, MEM_stage_inst_dmem_n8953, MEM_stage_inst_dmem_n8954, MEM_stage_inst_dmem_n21512, MEM_stage_inst_dmem_n8955, MEM_stage_inst_dmem_n8956, MEM_stage_inst_dmem_n21607, MEM_stage_inst_dmem_n8957, MEM_stage_inst_dmem_n21545, MEM_stage_inst_dmem_n8958, MEM_stage_inst_dmem_n8959, MEM_stage_inst_dmem_n8960, MEM_stage_inst_dmem_n8961, MEM_stage_inst_dmem_n8962, MEM_stage_inst_dmem_n8963, MEM_stage_inst_dmem_n8964, MEM_stage_inst_dmem_n8965, MEM_stage_inst_dmem_n21581, MEM_stage_inst_dmem_n8966, MEM_stage_inst_dmem_n8967, MEM_stage_inst_dmem_n8968, MEM_stage_inst_dmem_n8969, MEM_stage_inst_dmem_n8970, MEM_stage_inst_dmem_n8971, MEM_stage_inst_dmem_n8972, MEM_stage_inst_dmem_n8973, MEM_stage_inst_dmem_n21520, MEM_stage_inst_dmem_n8974, MEM_stage_inst_dmem_n8975, MEM_stage_inst_dmem_n21560, MEM_stage_inst_dmem_n8976, MEM_stage_inst_dmem_n8977, MEM_stage_inst_dmem_n8978, MEM_stage_inst_dmem_n8979, MEM_stage_inst_dmem_n8980, MEM_stage_inst_dmem_n8981, MEM_stage_inst_dmem_n8982, MEM_stage_inst_dmem_n8983, MEM_stage_inst_dmem_n8984, MEM_stage_inst_dmem_n8985, MEM_stage_inst_dmem_n8986, MEM_stage_inst_dmem_n8987, MEM_stage_inst_dmem_n8988, MEM_stage_inst_dmem_n21585, MEM_stage_inst_dmem_n8989, MEM_stage_inst_dmem_n8990, MEM_stage_inst_dmem_n8991, MEM_stage_inst_dmem_n8992, MEM_stage_inst_dmem_n8993, MEM_stage_inst_dmem_n8994, MEM_stage_inst_dmem_n8995, MEM_stage_inst_dmem_n8996, MEM_stage_inst_dmem_n8997, MEM_stage_inst_dmem_n21530, MEM_stage_inst_dmem_n8998, MEM_stage_inst_dmem_n8999, MEM_stage_inst_dmem_n21535, MEM_stage_inst_dmem_n9000, MEM_stage_inst_dmem_n9001, MEM_stage_inst_dmem_n9002, MEM_stage_inst_dmem_n9003, MEM_stage_inst_dmem_n9004, MEM_stage_inst_dmem_n9005, MEM_stage_inst_dmem_n9006, MEM_stage_inst_dmem_n9007, MEM_stage_inst_dmem_n9008, MEM_stage_inst_dmem_n9009, MEM_stage_inst_dmem_n9010, MEM_stage_inst_dmem_n9011, MEM_stage_inst_dmem_n21614, MEM_stage_inst_dmem_n9012, MEM_stage_inst_dmem_n9013, MEM_stage_inst_dmem_n9014, MEM_stage_inst_dmem_n9015, MEM_stage_inst_dmem_n9016, MEM_stage_inst_dmem_n9017, MEM_stage_inst_dmem_n21577, MEM_stage_inst_dmem_n9018, MEM_stage_inst_dmem_n9019, MEM_stage_inst_dmem_n9020, MEM_stage_inst_dmem_n9021, MEM_stage_inst_dmem_n9022, MEM_stage_inst_dmem_n9023, MEM_stage_inst_dmem_n9024, MEM_stage_inst_dmem_n9025, MEM_stage_inst_dmem_n9026, MEM_stage_inst_dmem_n9027, MEM_stage_inst_dmem_n9028, MEM_stage_inst_dmem_n9029, MEM_stage_inst_dmem_n9030, MEM_stage_inst_dmem_n9031, MEM_stage_inst_dmem_n21595, MEM_stage_inst_dmem_n9032, MEM_stage_inst_dmem_n9033, MEM_stage_inst_dmem_n9034, MEM_stage_inst_dmem_n9035, MEM_stage_inst_dmem_n21531, MEM_stage_inst_dmem_n9036, MEM_stage_inst_dmem_n9037, MEM_stage_inst_dmem_n9038, MEM_stage_inst_dmem_n9039, MEM_stage_inst_dmem_n9040, MEM_stage_inst_dmem_n9041, MEM_stage_inst_dmem_n9042, MEM_stage_inst_dmem_n9043, MEM_stage_inst_dmem_n9044, MEM_stage_inst_dmem_n9045, MEM_stage_inst_dmem_n9046, MEM_stage_inst_dmem_n9047, MEM_stage_inst_dmem_n9048, MEM_stage_inst_dmem_n9049, MEM_stage_inst_dmem_n9050, MEM_stage_inst_dmem_n9051, MEM_stage_inst_dmem_n21528, MEM_stage_inst_dmem_n9052, MEM_stage_inst_dmem_n9053, MEM_stage_inst_dmem_n9054, MEM_stage_inst_dmem_n9055, MEM_stage_inst_dmem_n9056, MEM_stage_inst_dmem_n9057, MEM_stage_inst_dmem_n9058, MEM_stage_inst_dmem_n9059, MEM_stage_inst_dmem_n9060, MEM_stage_inst_dmem_n9061, MEM_stage_inst_dmem_n9062, MEM_stage_inst_dmem_n9063, MEM_stage_inst_dmem_n9064, MEM_stage_inst_dmem_n21631, MEM_stage_inst_dmem_n9065, MEM_stage_inst_dmem_n9066, MEM_stage_inst_dmem_n21634, MEM_stage_inst_dmem_n9067, MEM_stage_inst_dmem_n9068, MEM_stage_inst_dmem_n9069, MEM_stage_inst_dmem_n9070, MEM_stage_inst_dmem_n21627, MEM_stage_inst_dmem_n9071, MEM_stage_inst_dmem_n9072, MEM_stage_inst_dmem_n9073, MEM_stage_inst_dmem_n9074, MEM_stage_inst_dmem_n9075, MEM_stage_inst_dmem_n9076, MEM_stage_inst_dmem_n9077, MEM_stage_inst_dmem_n9078, MEM_stage_inst_dmem_n9079, MEM_stage_inst_dmem_n21562, MEM_stage_inst_dmem_n9080, MEM_stage_inst_dmem_n9081, MEM_stage_inst_dmem_n21557, MEM_stage_inst_dmem_n9082, MEM_stage_inst_dmem_n9083, MEM_stage_inst_dmem_n9084, MEM_stage_inst_dmem_n9085, MEM_stage_inst_dmem_n9086, MEM_stage_inst_dmem_n9087, MEM_stage_inst_dmem_n9088, MEM_stage_inst_dmem_n9089, MEM_stage_inst_dmem_n9090, MEM_stage_inst_dmem_n9091, MEM_stage_inst_dmem_n9092, MEM_stage_inst_dmem_n9093, MEM_stage_inst_dmem_n9094, MEM_stage_inst_dmem_n9095, MEM_stage_inst_dmem_n21571, MEM_stage_inst_dmem_n9096, MEM_stage_inst_dmem_n9097, MEM_stage_inst_dmem_n9098, MEM_stage_inst_dmem_n9099, MEM_stage_inst_dmem_n9100, MEM_stage_inst_dmem_n9101, MEM_stage_inst_dmem_n9102, MEM_stage_inst_dmem_n9103, MEM_stage_inst_dmem_n9104, MEM_stage_inst_dmem_n9105, MEM_stage_inst_dmem_n9106, MEM_stage_inst_dmem_n9107, MEM_stage_inst_dmem_n9108, MEM_stage_inst_dmem_n9109, MEM_stage_inst_dmem_n9110, MEM_stage_inst_dmem_n9111, MEM_stage_inst_dmem_n9112, MEM_stage_inst_dmem_n9113, MEM_stage_inst_dmem_n21561, MEM_stage_inst_dmem_n9114, MEM_stage_inst_dmem_n9115, MEM_stage_inst_dmem_n9116, MEM_stage_inst_dmem_n9117, MEM_stage_inst_dmem_n9118, MEM_stage_inst_dmem_n9119, MEM_stage_inst_dmem_n9120, MEM_stage_inst_dmem_n9121, MEM_stage_inst_dmem_n9122, MEM_stage_inst_dmem_n9123, MEM_stage_inst_dmem_n9124, MEM_stage_inst_dmem_n9125, MEM_stage_inst_dmem_n9126, MEM_stage_inst_dmem_n9127, MEM_stage_inst_dmem_n9128, MEM_stage_inst_dmem_n9129, MEM_stage_inst_dmem_n9130, MEM_stage_inst_dmem_n9131, MEM_stage_inst_dmem_n21541, MEM_stage_inst_dmem_n9132, MEM_stage_inst_dmem_n9133, MEM_stage_inst_dmem_n9134, MEM_stage_inst_dmem_n9135, MEM_stage_inst_dmem_n21567, MEM_stage_inst_dmem_n9136, MEM_stage_inst_dmem_n9137, MEM_stage_inst_dmem_n9138, MEM_stage_inst_dmem_n9139, MEM_stage_inst_dmem_n9140, MEM_stage_inst_dmem_n9141, MEM_stage_inst_dmem_n9142, MEM_stage_inst_dmem_n9143, MEM_stage_inst_dmem_n9144, MEM_stage_inst_dmem_n9145, MEM_stage_inst_dmem_n9146, MEM_stage_inst_dmem_n9147, MEM_stage_inst_dmem_n9148, MEM_stage_inst_dmem_n9149, MEM_stage_inst_dmem_n9150, MEM_stage_inst_dmem_n9151, MEM_stage_inst_dmem_n9152, MEM_stage_inst_dmem_n9153, MEM_stage_inst_dmem_n9154, MEM_stage_inst_dmem_n9155, MEM_stage_inst_dmem_n9156, MEM_stage_inst_dmem_n9157, MEM_stage_inst_dmem_n9158, MEM_stage_inst_dmem_n9159, MEM_stage_inst_dmem_n9160, MEM_stage_inst_dmem_n9161, MEM_stage_inst_dmem_n9162, MEM_stage_inst_dmem_n9163, MEM_stage_inst_dmem_n9164, MEM_stage_inst_dmem_n9165, MEM_stage_inst_dmem_n9166, MEM_stage_inst_dmem_n9167, MEM_stage_inst_dmem_n9168, MEM_stage_inst_dmem_n9169, MEM_stage_inst_dmem_n9170, MEM_stage_inst_dmem_n9171, MEM_stage_inst_dmem_n9172, MEM_stage_inst_dmem_n9173, MEM_stage_inst_dmem_n9174, MEM_stage_inst_dmem_n9175, MEM_stage_inst_dmem_n9176, MEM_stage_inst_dmem_n9177, MEM_stage_inst_dmem_n9178, MEM_stage_inst_dmem_n9179, MEM_stage_inst_dmem_n9180, MEM_stage_inst_dmem_n9181, MEM_stage_inst_dmem_n9182, MEM_stage_inst_dmem_n9183, MEM_stage_inst_dmem_n9184, MEM_stage_inst_dmem_n9185, MEM_stage_inst_dmem_n9186, MEM_stage_inst_dmem_n9187, MEM_stage_inst_dmem_n9188, MEM_stage_inst_dmem_n9189, MEM_stage_inst_dmem_n9190, MEM_stage_inst_dmem_n9191, MEM_stage_inst_dmem_n9192, MEM_stage_inst_dmem_n9193, MEM_stage_inst_dmem_n9194, MEM_stage_inst_dmem_n9195, MEM_stage_inst_dmem_n21630, MEM_stage_inst_dmem_n9196, MEM_stage_inst_dmem_n9197, MEM_stage_inst_dmem_n9198, MEM_stage_inst_dmem_n9199, MEM_stage_inst_dmem_n9200, MEM_stage_inst_dmem_n9201, MEM_stage_inst_dmem_n9202, MEM_stage_inst_dmem_n9203, MEM_stage_inst_dmem_n9204, MEM_stage_inst_dmem_n9205, MEM_stage_inst_dmem_n9206, MEM_stage_inst_dmem_n9207, MEM_stage_inst_dmem_n9208, MEM_stage_inst_dmem_n9209, MEM_stage_inst_dmem_n9210, MEM_stage_inst_dmem_n9211, MEM_stage_inst_dmem_n9212, MEM_stage_inst_dmem_n9213, MEM_stage_inst_dmem_n9214, MEM_stage_inst_dmem_n9215, MEM_stage_inst_dmem_n9216, MEM_stage_inst_dmem_n9217, MEM_stage_inst_dmem_n9218, MEM_stage_inst_dmem_n9219, MEM_stage_inst_dmem_n9220, MEM_stage_inst_dmem_n9221, MEM_stage_inst_dmem_n9222, MEM_stage_inst_dmem_n9223, MEM_stage_inst_dmem_n9224, MEM_stage_inst_dmem_n9225, MEM_stage_inst_dmem_n9226, MEM_stage_inst_dmem_n9227, MEM_stage_inst_dmem_n9228, MEM_stage_inst_dmem_n9229, MEM_stage_inst_dmem_n9230, MEM_stage_inst_dmem_n9231, MEM_stage_inst_dmem_n9232, MEM_stage_inst_dmem_n9233, MEM_stage_inst_dmem_n9234, MEM_stage_inst_dmem_n9235, MEM_stage_inst_dmem_n9236, MEM_stage_inst_dmem_n9237, MEM_stage_inst_dmem_n9238, MEM_stage_inst_dmem_n9239, MEM_stage_inst_dmem_n9240, MEM_stage_inst_dmem_n9241, MEM_stage_inst_dmem_n21521, MEM_stage_inst_dmem_n9242, MEM_stage_inst_dmem_n9243, MEM_stage_inst_dmem_n9244, MEM_stage_inst_dmem_n9245, MEM_stage_inst_dmem_n9246, MEM_stage_inst_dmem_n9247, MEM_stage_inst_dmem_n9248, MEM_stage_inst_dmem_n9249, MEM_stage_inst_dmem_n9250, MEM_stage_inst_dmem_n9251, MEM_stage_inst_dmem_n9252, MEM_stage_inst_dmem_n9253, MEM_stage_inst_dmem_n9254, MEM_stage_inst_dmem_n9255, MEM_stage_inst_dmem_n9256, MEM_stage_inst_dmem_n9257, MEM_stage_inst_dmem_n9258, MEM_stage_inst_dmem_n9259, MEM_stage_inst_dmem_n9260, MEM_stage_inst_dmem_n9261, MEM_stage_inst_dmem_n9262, MEM_stage_inst_dmem_n9263, MEM_stage_inst_dmem_n9264, MEM_stage_inst_dmem_n9265, MEM_stage_inst_dmem_n9266, MEM_stage_inst_dmem_n9267, MEM_stage_inst_dmem_n9268, MEM_stage_inst_dmem_n9269, MEM_stage_inst_dmem_n9270, MEM_stage_inst_dmem_n9271, MEM_stage_inst_dmem_n9272, MEM_stage_inst_dmem_n9273, MEM_stage_inst_dmem_n9274, MEM_stage_inst_dmem_n9275, MEM_stage_inst_dmem_n9276, MEM_stage_inst_dmem_n9277, MEM_stage_inst_dmem_n9278, MEM_stage_inst_dmem_n9279, MEM_stage_inst_dmem_n9280, MEM_stage_inst_dmem_n9281, MEM_stage_inst_dmem_n9282, MEM_stage_inst_dmem_n9283, MEM_stage_inst_dmem_n9284, MEM_stage_inst_dmem_n9285, MEM_stage_inst_dmem_n9286, MEM_stage_inst_dmem_n9287, MEM_stage_inst_dmem_n9288, MEM_stage_inst_dmem_n9289, MEM_stage_inst_dmem_n9290, MEM_stage_inst_dmem_n9291, MEM_stage_inst_dmem_n9292, MEM_stage_inst_dmem_n9293, MEM_stage_inst_dmem_n9294, MEM_stage_inst_dmem_n9295, MEM_stage_inst_dmem_n9296, MEM_stage_inst_dmem_n9297, MEM_stage_inst_dmem_n9298, MEM_stage_inst_dmem_n9299, MEM_stage_inst_dmem_n9300, MEM_stage_inst_dmem_n9301, MEM_stage_inst_dmem_n9302, MEM_stage_inst_dmem_n9303, MEM_stage_inst_dmem_n9304, MEM_stage_inst_dmem_n9305, MEM_stage_inst_dmem_n9306, MEM_stage_inst_dmem_n9307, MEM_stage_inst_dmem_n9308, MEM_stage_inst_dmem_n9309, MEM_stage_inst_dmem_n9310, MEM_stage_inst_dmem_n9311, MEM_stage_inst_dmem_n9312, MEM_stage_inst_dmem_n9313, MEM_stage_inst_dmem_n9314, MEM_stage_inst_dmem_n9315, MEM_stage_inst_dmem_n9316, MEM_stage_inst_dmem_n9317, MEM_stage_inst_dmem_n9318, MEM_stage_inst_dmem_n9319, MEM_stage_inst_dmem_n9320, MEM_stage_inst_dmem_n9321, MEM_stage_inst_dmem_n9322, MEM_stage_inst_dmem_n9323, MEM_stage_inst_dmem_n9324, MEM_stage_inst_dmem_n9325, MEM_stage_inst_dmem_n9326, MEM_stage_inst_dmem_n9327, MEM_stage_inst_dmem_n9328, MEM_stage_inst_dmem_n9329, MEM_stage_inst_dmem_n9330, MEM_stage_inst_dmem_n9331, MEM_stage_inst_dmem_n9332, MEM_stage_inst_dmem_n9333, MEM_stage_inst_dmem_n9334, MEM_stage_inst_dmem_n9335, MEM_stage_inst_dmem_n9336, MEM_stage_inst_dmem_n9337, MEM_stage_inst_dmem_n9338, MEM_stage_inst_dmem_n9339, MEM_stage_inst_dmem_n9340, MEM_stage_inst_dmem_n9341, MEM_stage_inst_dmem_n9342, MEM_stage_inst_dmem_n9343, MEM_stage_inst_dmem_n9344, MEM_stage_inst_dmem_n9345, MEM_stage_inst_dmem_n9346, MEM_stage_inst_dmem_n9347, MEM_stage_inst_dmem_n9348, MEM_stage_inst_dmem_n9349, MEM_stage_inst_dmem_n9350, MEM_stage_inst_dmem_n9351, MEM_stage_inst_dmem_n9352, MEM_stage_inst_dmem_n9353, MEM_stage_inst_dmem_n9354, MEM_stage_inst_dmem_n9355, MEM_stage_inst_dmem_n9356, MEM_stage_inst_dmem_n9357, MEM_stage_inst_dmem_n9358, MEM_stage_inst_dmem_n9359, MEM_stage_inst_dmem_n9360, MEM_stage_inst_dmem_n9361, MEM_stage_inst_dmem_n9362, MEM_stage_inst_dmem_n9363, MEM_stage_inst_dmem_n9364, MEM_stage_inst_dmem_n9365, MEM_stage_inst_dmem_n9366, MEM_stage_inst_dmem_n9367, MEM_stage_inst_dmem_n9368, MEM_stage_inst_dmem_n9369, MEM_stage_inst_dmem_n9370, MEM_stage_inst_dmem_n9371, MEM_stage_inst_dmem_n9372, MEM_stage_inst_dmem_n9373, MEM_stage_inst_dmem_n9374, MEM_stage_inst_dmem_n9375, MEM_stage_inst_dmem_n9376, MEM_stage_inst_dmem_n9377, MEM_stage_inst_dmem_n9378, MEM_stage_inst_dmem_n9379, MEM_stage_inst_dmem_n9380, MEM_stage_inst_dmem_n9381, MEM_stage_inst_dmem_n9382, MEM_stage_inst_dmem_n9383, MEM_stage_inst_dmem_n9384, MEM_stage_inst_dmem_n9385, MEM_stage_inst_dmem_n9386, MEM_stage_inst_dmem_n9387, MEM_stage_inst_dmem_n9388, MEM_stage_inst_dmem_n9389, MEM_stage_inst_dmem_n9390, MEM_stage_inst_dmem_n9391, MEM_stage_inst_dmem_n9392, MEM_stage_inst_dmem_n9393, MEM_stage_inst_dmem_n9394, MEM_stage_inst_dmem_n9395, MEM_stage_inst_dmem_n9396, MEM_stage_inst_dmem_n21533, MEM_stage_inst_dmem_n9397, MEM_stage_inst_dmem_n9398, MEM_stage_inst_dmem_n9399, MEM_stage_inst_dmem_n9400, MEM_stage_inst_dmem_n9401, MEM_stage_inst_dmem_n9402, MEM_stage_inst_dmem_n21637, MEM_stage_inst_dmem_n9403, MEM_stage_inst_dmem_n9404, MEM_stage_inst_dmem_n9405, MEM_stage_inst_dmem_n9406, MEM_stage_inst_dmem_n9407, MEM_stage_inst_dmem_n9408, MEM_stage_inst_dmem_n9409, MEM_stage_inst_dmem_n9410, MEM_stage_inst_dmem_n9411, MEM_stage_inst_dmem_n9412, MEM_stage_inst_dmem_n9413, MEM_stage_inst_dmem_n9414, MEM_stage_inst_dmem_n9415, MEM_stage_inst_dmem_n9416, MEM_stage_inst_dmem_n9417, MEM_stage_inst_dmem_n9418, MEM_stage_inst_dmem_n9419, MEM_stage_inst_dmem_n9420, MEM_stage_inst_dmem_n9421, MEM_stage_inst_dmem_n9422, MEM_stage_inst_dmem_n9423, MEM_stage_inst_dmem_n9424, MEM_stage_inst_dmem_n9425, MEM_stage_inst_dmem_n9426, MEM_stage_inst_dmem_n9427, MEM_stage_inst_dmem_n9428, MEM_stage_inst_dmem_n9429, MEM_stage_inst_dmem_n9430, MEM_stage_inst_dmem_n9431, MEM_stage_inst_dmem_n9432, MEM_stage_inst_dmem_n9433, MEM_stage_inst_dmem_n9434, MEM_stage_inst_dmem_n9435, MEM_stage_inst_dmem_n9436, MEM_stage_inst_dmem_n9437, MEM_stage_inst_dmem_n9438, MEM_stage_inst_dmem_n9439, MEM_stage_inst_dmem_n9440, MEM_stage_inst_dmem_n9441, MEM_stage_inst_dmem_n9442, MEM_stage_inst_dmem_n9443, MEM_stage_inst_dmem_n9444, MEM_stage_inst_dmem_n9445, MEM_stage_inst_dmem_n9446, MEM_stage_inst_dmem_n9447, MEM_stage_inst_dmem_n9448, MEM_stage_inst_dmem_n9449, MEM_stage_inst_dmem_n9450, MEM_stage_inst_dmem_n9451, MEM_stage_inst_dmem_n9452, MEM_stage_inst_dmem_n9453, MEM_stage_inst_dmem_n9454, MEM_stage_inst_dmem_n9455, MEM_stage_inst_dmem_n9456, MEM_stage_inst_dmem_n9457, MEM_stage_inst_dmem_n9458, MEM_stage_inst_dmem_n9459, MEM_stage_inst_dmem_n9460, MEM_stage_inst_dmem_n9461, MEM_stage_inst_dmem_n9462, MEM_stage_inst_dmem_n9463, MEM_stage_inst_dmem_n9464, MEM_stage_inst_dmem_n9465, MEM_stage_inst_dmem_n9466, MEM_stage_inst_dmem_n9467, MEM_stage_inst_dmem_n9468, MEM_stage_inst_dmem_n9469, MEM_stage_inst_dmem_n9470, MEM_stage_inst_dmem_n9471, MEM_stage_inst_dmem_n9472, MEM_stage_inst_dmem_n9473, MEM_stage_inst_dmem_n9474, MEM_stage_inst_dmem_n9475, MEM_stage_inst_dmem_n9476, MEM_stage_inst_dmem_n9477, MEM_stage_inst_dmem_n9478, MEM_stage_inst_dmem_n9479, MEM_stage_inst_dmem_n9480, MEM_stage_inst_dmem_n9481, MEM_stage_inst_dmem_n9482, MEM_stage_inst_dmem_n9483, MEM_stage_inst_dmem_n9484, MEM_stage_inst_dmem_n9485, MEM_stage_inst_dmem_n9486, MEM_stage_inst_dmem_n9487, MEM_stage_inst_dmem_n9488, MEM_stage_inst_dmem_n9489, MEM_stage_inst_dmem_n9490, MEM_stage_inst_dmem_n9491, MEM_stage_inst_dmem_n9492, MEM_stage_inst_dmem_n9493, MEM_stage_inst_dmem_n9494, MEM_stage_inst_dmem_n9495, MEM_stage_inst_dmem_n9496, MEM_stage_inst_dmem_n9497, MEM_stage_inst_dmem_n21536, MEM_stage_inst_dmem_n9498, MEM_stage_inst_dmem_n9499, MEM_stage_inst_dmem_n9500, MEM_stage_inst_dmem_n9501, MEM_stage_inst_dmem_n9502, MEM_stage_inst_dmem_n9503, MEM_stage_inst_dmem_n9504, MEM_stage_inst_dmem_n9505, MEM_stage_inst_dmem_n9506, MEM_stage_inst_dmem_n9507, MEM_stage_inst_dmem_n9508, MEM_stage_inst_dmem_n9509, MEM_stage_inst_dmem_n9510, MEM_stage_inst_dmem_n9511, MEM_stage_inst_dmem_n9512, MEM_stage_inst_dmem_n9513, MEM_stage_inst_dmem_n9514, MEM_stage_inst_dmem_n9515, MEM_stage_inst_dmem_n9516, MEM_stage_inst_dmem_n9517, MEM_stage_inst_dmem_n9518, MEM_stage_inst_dmem_n9519, MEM_stage_inst_dmem_n9520, MEM_stage_inst_dmem_n9521, MEM_stage_inst_dmem_n9522, MEM_stage_inst_dmem_n9523, MEM_stage_inst_dmem_n9524, MEM_stage_inst_dmem_n9525, MEM_stage_inst_dmem_n9526, MEM_stage_inst_dmem_n9527, MEM_stage_inst_dmem_n9528, MEM_stage_inst_dmem_n9529, MEM_stage_inst_dmem_n9530, MEM_stage_inst_dmem_n9531, MEM_stage_inst_dmem_n9532, MEM_stage_inst_dmem_n9533, MEM_stage_inst_dmem_n9534, MEM_stage_inst_dmem_n9535, MEM_stage_inst_dmem_n9536, MEM_stage_inst_dmem_n9537, MEM_stage_inst_dmem_n9538, MEM_stage_inst_dmem_n9539, MEM_stage_inst_dmem_n9540, MEM_stage_inst_dmem_n9541, MEM_stage_inst_dmem_n9542, MEM_stage_inst_dmem_n9543, MEM_stage_inst_dmem_n9544, MEM_stage_inst_dmem_n9545, MEM_stage_inst_dmem_n9546, MEM_stage_inst_dmem_n9547, MEM_stage_inst_dmem_n9548, MEM_stage_inst_dmem_n9549, MEM_stage_inst_dmem_n9550, MEM_stage_inst_dmem_n9551, MEM_stage_inst_dmem_n9552, MEM_stage_inst_dmem_n9553, MEM_stage_inst_dmem_n9554, MEM_stage_inst_dmem_n9555, MEM_stage_inst_dmem_n9556, MEM_stage_inst_dmem_n9557, MEM_stage_inst_dmem_n9558, MEM_stage_inst_dmem_n9559, MEM_stage_inst_dmem_n9560, MEM_stage_inst_dmem_n9561, MEM_stage_inst_dmem_n9562, MEM_stage_inst_dmem_n9563, MEM_stage_inst_dmem_n9564, MEM_stage_inst_dmem_n9565, MEM_stage_inst_dmem_n9566, MEM_stage_inst_dmem_n9567, MEM_stage_inst_dmem_n9568, MEM_stage_inst_dmem_n9569, MEM_stage_inst_dmem_n9570, MEM_stage_inst_dmem_n9571, MEM_stage_inst_dmem_n9572, MEM_stage_inst_dmem_n9573, MEM_stage_inst_dmem_n9574, MEM_stage_inst_dmem_n9575, MEM_stage_inst_dmem_n9576, MEM_stage_inst_dmem_n9577, MEM_stage_inst_dmem_n9578, MEM_stage_inst_dmem_n9579, MEM_stage_inst_dmem_n9580, MEM_stage_inst_dmem_n9581, MEM_stage_inst_dmem_n9582, MEM_stage_inst_dmem_n9583, MEM_stage_inst_dmem_n9584, MEM_stage_inst_dmem_n9585, MEM_stage_inst_dmem_n9586, MEM_stage_inst_dmem_n9587, MEM_stage_inst_dmem_n9588, MEM_stage_inst_dmem_n9589, MEM_stage_inst_dmem_n9590, MEM_stage_inst_dmem_n9591, MEM_stage_inst_dmem_n9592, MEM_stage_inst_dmem_n9593, MEM_stage_inst_dmem_n9594, MEM_stage_inst_dmem_n9595, MEM_stage_inst_dmem_n9596, MEM_stage_inst_dmem_n9597, MEM_stage_inst_dmem_n9598, MEM_stage_inst_dmem_n9599, MEM_stage_inst_dmem_n9600, MEM_stage_inst_dmem_n9601, MEM_stage_inst_dmem_n9602, MEM_stage_inst_dmem_n9603, MEM_stage_inst_dmem_n9604, MEM_stage_inst_dmem_n9605, MEM_stage_inst_dmem_n9606, MEM_stage_inst_dmem_n9607, MEM_stage_inst_dmem_n9608, MEM_stage_inst_dmem_n9609, MEM_stage_inst_dmem_n9610, MEM_stage_inst_dmem_n9611, MEM_stage_inst_dmem_n9612, MEM_stage_inst_dmem_n9613, MEM_stage_inst_dmem_n9614, MEM_stage_inst_dmem_n9615, MEM_stage_inst_dmem_n9616, MEM_stage_inst_dmem_n9617, MEM_stage_inst_dmem_n9618, MEM_stage_inst_dmem_n9619, MEM_stage_inst_dmem_n9620, MEM_stage_inst_dmem_n9621, MEM_stage_inst_dmem_n9622, MEM_stage_inst_dmem_n9623, MEM_stage_inst_dmem_n9624, MEM_stage_inst_dmem_n9625, MEM_stage_inst_dmem_n9626, MEM_stage_inst_dmem_n9627, MEM_stage_inst_dmem_n9628, MEM_stage_inst_dmem_n9629, MEM_stage_inst_dmem_n9630, MEM_stage_inst_dmem_n9631, MEM_stage_inst_dmem_n9632, MEM_stage_inst_dmem_n9633, MEM_stage_inst_dmem_n9634, MEM_stage_inst_dmem_n9635, MEM_stage_inst_dmem_n9636, MEM_stage_inst_dmem_n9637, MEM_stage_inst_dmem_n9638, MEM_stage_inst_dmem_n9639, MEM_stage_inst_dmem_n9640, MEM_stage_inst_dmem_n9641, MEM_stage_inst_dmem_n9642, MEM_stage_inst_dmem_n9643, MEM_stage_inst_dmem_n9644, MEM_stage_inst_dmem_n9645, MEM_stage_inst_dmem_n9646, MEM_stage_inst_dmem_n9647, MEM_stage_inst_dmem_n9648, MEM_stage_inst_dmem_n9649, MEM_stage_inst_dmem_n9650, MEM_stage_inst_dmem_n9651, MEM_stage_inst_dmem_n9652, MEM_stage_inst_dmem_n9653, MEM_stage_inst_dmem_n9654, MEM_stage_inst_dmem_n9655, MEM_stage_inst_dmem_n9656, MEM_stage_inst_dmem_n9657, MEM_stage_inst_dmem_n9658, MEM_stage_inst_dmem_n9659, MEM_stage_inst_dmem_n9660, MEM_stage_inst_dmem_n9661, MEM_stage_inst_dmem_n9662, MEM_stage_inst_dmem_n9663, MEM_stage_inst_dmem_n9664, MEM_stage_inst_dmem_n9665, MEM_stage_inst_dmem_n9666, MEM_stage_inst_dmem_n9667, MEM_stage_inst_dmem_n9668, MEM_stage_inst_dmem_n9669, MEM_stage_inst_dmem_n9670, MEM_stage_inst_dmem_n9671, MEM_stage_inst_dmem_n9672, MEM_stage_inst_dmem_n9673, MEM_stage_inst_dmem_n9674, MEM_stage_inst_dmem_n9675, MEM_stage_inst_dmem_n9676, MEM_stage_inst_dmem_n9677, MEM_stage_inst_dmem_n9678, MEM_stage_inst_dmem_n9679, MEM_stage_inst_dmem_n9680, MEM_stage_inst_dmem_n9681, MEM_stage_inst_dmem_n9682, MEM_stage_inst_dmem_n9683, MEM_stage_inst_dmem_n9684, MEM_stage_inst_dmem_n9685, MEM_stage_inst_dmem_n9686, MEM_stage_inst_dmem_n9687, MEM_stage_inst_dmem_n9688, MEM_stage_inst_dmem_n9689, MEM_stage_inst_dmem_n9690, MEM_stage_inst_dmem_n9691, MEM_stage_inst_dmem_n9692, MEM_stage_inst_dmem_n9693, MEM_stage_inst_dmem_n9694, MEM_stage_inst_dmem_n9695, MEM_stage_inst_dmem_n9696, MEM_stage_inst_dmem_n9697, MEM_stage_inst_dmem_n9698, MEM_stage_inst_dmem_n9699, MEM_stage_inst_dmem_n9700, MEM_stage_inst_dmem_n9701, MEM_stage_inst_dmem_n9702, MEM_stage_inst_dmem_n9703, MEM_stage_inst_dmem_n9704, MEM_stage_inst_dmem_n9705, MEM_stage_inst_dmem_n9706, MEM_stage_inst_dmem_n9707, MEM_stage_inst_dmem_n9708, MEM_stage_inst_dmem_n9709, MEM_stage_inst_dmem_n9710, MEM_stage_inst_dmem_n9711, MEM_stage_inst_dmem_n9712, MEM_stage_inst_dmem_n9713, MEM_stage_inst_dmem_n9714, MEM_stage_inst_dmem_n9715, MEM_stage_inst_dmem_n9716, MEM_stage_inst_dmem_n9717, MEM_stage_inst_dmem_n9718, MEM_stage_inst_dmem_n9719, MEM_stage_inst_dmem_n9720, MEM_stage_inst_dmem_n9721, MEM_stage_inst_dmem_n9722, MEM_stage_inst_dmem_n9723, MEM_stage_inst_dmem_n9724, MEM_stage_inst_dmem_n9725, MEM_stage_inst_dmem_n9726, MEM_stage_inst_dmem_n9727, MEM_stage_inst_dmem_n9728, MEM_stage_inst_dmem_n9729, MEM_stage_inst_dmem_n9730, MEM_stage_inst_dmem_n9731, MEM_stage_inst_dmem_n9732, MEM_stage_inst_dmem_n9733, MEM_stage_inst_dmem_n9734, MEM_stage_inst_dmem_n9735, MEM_stage_inst_dmem_n9736, MEM_stage_inst_dmem_n9737, MEM_stage_inst_dmem_n9738, MEM_stage_inst_dmem_n9739, MEM_stage_inst_dmem_n9740, MEM_stage_inst_dmem_n9741, MEM_stage_inst_dmem_n9742, MEM_stage_inst_dmem_n9743, MEM_stage_inst_dmem_n9744, MEM_stage_inst_dmem_n9745, MEM_stage_inst_dmem_n9746, MEM_stage_inst_dmem_n9747, MEM_stage_inst_dmem_n9748, MEM_stage_inst_dmem_n9749, MEM_stage_inst_dmem_n9750, MEM_stage_inst_dmem_n9751, MEM_stage_inst_dmem_n9752, MEM_stage_inst_dmem_n9753, MEM_stage_inst_dmem_n9754, MEM_stage_inst_dmem_n9755, MEM_stage_inst_dmem_n9756, MEM_stage_inst_dmem_n9757, MEM_stage_inst_dmem_n9758, MEM_stage_inst_dmem_n9759, MEM_stage_inst_dmem_n9760, MEM_stage_inst_dmem_n9761, MEM_stage_inst_dmem_n9762, MEM_stage_inst_dmem_n9763, MEM_stage_inst_dmem_n9764, MEM_stage_inst_dmem_n9765, MEM_stage_inst_dmem_n9766, MEM_stage_inst_dmem_n9767, MEM_stage_inst_dmem_n9768, MEM_stage_inst_dmem_n9769, MEM_stage_inst_dmem_n9770, MEM_stage_inst_dmem_n9771, MEM_stage_inst_dmem_n9772, MEM_stage_inst_dmem_n9773, MEM_stage_inst_dmem_n9774, MEM_stage_inst_dmem_n9775, MEM_stage_inst_dmem_n9776, MEM_stage_inst_dmem_n9777, MEM_stage_inst_dmem_n9778, MEM_stage_inst_dmem_n9779, MEM_stage_inst_dmem_n9780, MEM_stage_inst_dmem_n9781, MEM_stage_inst_dmem_n9782, MEM_stage_inst_dmem_n9783, MEM_stage_inst_dmem_n9784, MEM_stage_inst_dmem_n9785, MEM_stage_inst_dmem_n9786, MEM_stage_inst_dmem_n9787, MEM_stage_inst_dmem_n9788, MEM_stage_inst_dmem_n9789, MEM_stage_inst_dmem_n9790, MEM_stage_inst_dmem_n9791, MEM_stage_inst_dmem_n9792, MEM_stage_inst_dmem_n9793, MEM_stage_inst_dmem_n9794, MEM_stage_inst_dmem_n9795, MEM_stage_inst_dmem_n9796, MEM_stage_inst_dmem_n9797, MEM_stage_inst_dmem_n9798, MEM_stage_inst_dmem_n9799, MEM_stage_inst_dmem_n9800, MEM_stage_inst_dmem_n9801, MEM_stage_inst_dmem_n9802, MEM_stage_inst_dmem_n9803, MEM_stage_inst_dmem_n9804, MEM_stage_inst_dmem_n9805, MEM_stage_inst_dmem_n9806, MEM_stage_inst_dmem_n9807, MEM_stage_inst_dmem_n9808, MEM_stage_inst_dmem_n9809, MEM_stage_inst_dmem_n9810, MEM_stage_inst_dmem_n9811, MEM_stage_inst_dmem_n9812, MEM_stage_inst_dmem_n9813, MEM_stage_inst_dmem_n9814, MEM_stage_inst_dmem_n9815, MEM_stage_inst_dmem_n9816, MEM_stage_inst_dmem_n9817, MEM_stage_inst_dmem_n9818, MEM_stage_inst_dmem_n9819, MEM_stage_inst_dmem_n9820, MEM_stage_inst_dmem_n9821, MEM_stage_inst_dmem_n9822, MEM_stage_inst_dmem_n9823, MEM_stage_inst_dmem_n9824, MEM_stage_inst_dmem_n9825, MEM_stage_inst_dmem_n9826, MEM_stage_inst_dmem_n9827, MEM_stage_inst_dmem_n9828, MEM_stage_inst_dmem_n9829, MEM_stage_inst_dmem_n9830, MEM_stage_inst_dmem_n9831, MEM_stage_inst_dmem_n9832, MEM_stage_inst_dmem_n9833, MEM_stage_inst_dmem_n9834, MEM_stage_inst_dmem_n9835, MEM_stage_inst_dmem_n9836, MEM_stage_inst_dmem_n9837, MEM_stage_inst_dmem_n9838, MEM_stage_inst_dmem_n9839, MEM_stage_inst_dmem_n9840, MEM_stage_inst_dmem_n9841, MEM_stage_inst_dmem_n9842, MEM_stage_inst_dmem_n9843, MEM_stage_inst_dmem_n9844, MEM_stage_inst_dmem_n9845, MEM_stage_inst_dmem_n9846, MEM_stage_inst_dmem_n9847, MEM_stage_inst_dmem_n9848, MEM_stage_inst_dmem_n9849, MEM_stage_inst_dmem_n9850, MEM_stage_inst_dmem_n9851, MEM_stage_inst_dmem_n9852, MEM_stage_inst_dmem_n9853, MEM_stage_inst_dmem_n9854, MEM_stage_inst_dmem_n9855, MEM_stage_inst_dmem_n9856, MEM_stage_inst_dmem_n9857, MEM_stage_inst_dmem_n9858, MEM_stage_inst_dmem_n9859, MEM_stage_inst_dmem_n9860, MEM_stage_inst_dmem_n9861, MEM_stage_inst_dmem_n9862, MEM_stage_inst_dmem_n9863, MEM_stage_inst_dmem_n9864, MEM_stage_inst_dmem_n9865, MEM_stage_inst_dmem_n9866, MEM_stage_inst_dmem_n9867, MEM_stage_inst_dmem_n9868, MEM_stage_inst_dmem_n9869, MEM_stage_inst_dmem_n9870, MEM_stage_inst_dmem_n9871, MEM_stage_inst_dmem_n9872, MEM_stage_inst_dmem_n9873, MEM_stage_inst_dmem_n9874, MEM_stage_inst_dmem_n9875, MEM_stage_inst_dmem_n9876, MEM_stage_inst_dmem_n9877, MEM_stage_inst_dmem_n9878, MEM_stage_inst_dmem_n9879, MEM_stage_inst_dmem_n9880, MEM_stage_inst_dmem_n9881, MEM_stage_inst_dmem_n9882, MEM_stage_inst_dmem_n9883, MEM_stage_inst_dmem_n9884, MEM_stage_inst_dmem_n9885, MEM_stage_inst_dmem_n9886, MEM_stage_inst_dmem_n9887, MEM_stage_inst_dmem_n9888, MEM_stage_inst_dmem_n9889, MEM_stage_inst_dmem_n9890, MEM_stage_inst_dmem_n9891, MEM_stage_inst_dmem_n9892, MEM_stage_inst_dmem_n9893, MEM_stage_inst_dmem_n9894, MEM_stage_inst_dmem_n9895, MEM_stage_inst_dmem_n9896, MEM_stage_inst_dmem_n9897, MEM_stage_inst_dmem_n9898, MEM_stage_inst_dmem_n9899, MEM_stage_inst_dmem_n9900, MEM_stage_inst_dmem_n9901, MEM_stage_inst_dmem_n9902, MEM_stage_inst_dmem_n9903, MEM_stage_inst_dmem_n9904, MEM_stage_inst_dmem_n9905, MEM_stage_inst_dmem_n9906, MEM_stage_inst_dmem_n9907, MEM_stage_inst_dmem_n9908, MEM_stage_inst_dmem_n9909, MEM_stage_inst_dmem_n9910, MEM_stage_inst_dmem_n9911, MEM_stage_inst_dmem_n9912, MEM_stage_inst_dmem_n9913, MEM_stage_inst_dmem_n9914, MEM_stage_inst_dmem_n9915, MEM_stage_inst_dmem_n9916, MEM_stage_inst_dmem_n9917, MEM_stage_inst_dmem_n9918, MEM_stage_inst_dmem_n9919, MEM_stage_inst_dmem_n9920, MEM_stage_inst_dmem_n9921, MEM_stage_inst_dmem_n9922, MEM_stage_inst_dmem_n9923, MEM_stage_inst_dmem_n9924, MEM_stage_inst_dmem_n9925, MEM_stage_inst_dmem_n9926, MEM_stage_inst_dmem_n9927, MEM_stage_inst_dmem_n9928, MEM_stage_inst_dmem_n9929, MEM_stage_inst_dmem_n9930, MEM_stage_inst_dmem_n9931, MEM_stage_inst_dmem_n9932, MEM_stage_inst_dmem_n9933, MEM_stage_inst_dmem_n9934, MEM_stage_inst_dmem_n9935, MEM_stage_inst_dmem_n9936, MEM_stage_inst_dmem_n9937, MEM_stage_inst_dmem_n9938, MEM_stage_inst_dmem_n9939, MEM_stage_inst_dmem_n9940, MEM_stage_inst_dmem_n9941, MEM_stage_inst_dmem_n9942, MEM_stage_inst_dmem_n9943, MEM_stage_inst_dmem_n9944, MEM_stage_inst_dmem_n9945, MEM_stage_inst_dmem_n9946, MEM_stage_inst_dmem_n9947, MEM_stage_inst_dmem_n9948, MEM_stage_inst_dmem_n9949, MEM_stage_inst_dmem_n9950, MEM_stage_inst_dmem_n9951, MEM_stage_inst_dmem_n9952, MEM_stage_inst_dmem_n9953, MEM_stage_inst_dmem_n9954, MEM_stage_inst_dmem_n9955, MEM_stage_inst_dmem_n9956, MEM_stage_inst_dmem_n9957, MEM_stage_inst_dmem_n9958, MEM_stage_inst_dmem_n9959, MEM_stage_inst_dmem_n9960, MEM_stage_inst_dmem_n9961, MEM_stage_inst_dmem_n9962, MEM_stage_inst_dmem_n9963, MEM_stage_inst_dmem_n9964, MEM_stage_inst_dmem_n9965, MEM_stage_inst_dmem_n9966, MEM_stage_inst_dmem_n9967, MEM_stage_inst_dmem_n9968, MEM_stage_inst_dmem_n9969, MEM_stage_inst_dmem_n9970, MEM_stage_inst_dmem_n9971, MEM_stage_inst_dmem_n9972, MEM_stage_inst_dmem_n9973, MEM_stage_inst_dmem_n9974, MEM_stage_inst_dmem_n9975, MEM_stage_inst_dmem_n9976, MEM_stage_inst_dmem_n9977, MEM_stage_inst_dmem_n9978, MEM_stage_inst_dmem_n9979, MEM_stage_inst_dmem_n9980, MEM_stage_inst_dmem_n9981, MEM_stage_inst_dmem_n9982, MEM_stage_inst_dmem_n9983, MEM_stage_inst_dmem_n9984, MEM_stage_inst_dmem_n9985, MEM_stage_inst_dmem_n9986, MEM_stage_inst_dmem_n9987, MEM_stage_inst_dmem_n9988, MEM_stage_inst_dmem_n9989, MEM_stage_inst_dmem_n9990, MEM_stage_inst_dmem_n9991, MEM_stage_inst_dmem_n9992, MEM_stage_inst_dmem_n9993, MEM_stage_inst_dmem_n9994, MEM_stage_inst_dmem_n9995, MEM_stage_inst_dmem_n9996, MEM_stage_inst_dmem_n9997, MEM_stage_inst_dmem_n9998, MEM_stage_inst_dmem_n9999, MEM_stage_inst_dmem_n10000, MEM_stage_inst_dmem_n10001, MEM_stage_inst_dmem_n10002, MEM_stage_inst_dmem_n10003, MEM_stage_inst_dmem_n10004, MEM_stage_inst_dmem_n10005, MEM_stage_inst_dmem_n10006, MEM_stage_inst_dmem_n10007, MEM_stage_inst_dmem_n10008, MEM_stage_inst_dmem_n10009, MEM_stage_inst_dmem_n10010, MEM_stage_inst_dmem_n10011, MEM_stage_inst_dmem_n10012, MEM_stage_inst_dmem_n10013, MEM_stage_inst_dmem_n10014, MEM_stage_inst_dmem_n10015, MEM_stage_inst_dmem_n10016, MEM_stage_inst_dmem_n10017, MEM_stage_inst_dmem_n10018, MEM_stage_inst_dmem_n10019, MEM_stage_inst_dmem_n10020, MEM_stage_inst_dmem_n10021, MEM_stage_inst_dmem_n10022, MEM_stage_inst_dmem_n10023, MEM_stage_inst_dmem_n10024, MEM_stage_inst_dmem_n10025, MEM_stage_inst_dmem_n10026, MEM_stage_inst_dmem_n10027, MEM_stage_inst_dmem_n10028, MEM_stage_inst_dmem_n10029, MEM_stage_inst_dmem_n10030, MEM_stage_inst_dmem_n10031, MEM_stage_inst_dmem_n10032, MEM_stage_inst_dmem_n10033, MEM_stage_inst_dmem_n10034, MEM_stage_inst_dmem_n10035, MEM_stage_inst_dmem_n10036, MEM_stage_inst_dmem_n10037, MEM_stage_inst_dmem_n10038, MEM_stage_inst_dmem_n10039, MEM_stage_inst_dmem_n10040, MEM_stage_inst_dmem_n10041, MEM_stage_inst_dmem_n10042, MEM_stage_inst_dmem_n10043, MEM_stage_inst_dmem_n10044, MEM_stage_inst_dmem_n10045, MEM_stage_inst_dmem_n10046, MEM_stage_inst_dmem_n10047, MEM_stage_inst_dmem_n10048, MEM_stage_inst_dmem_n10049, MEM_stage_inst_dmem_n10050, MEM_stage_inst_dmem_n10051, MEM_stage_inst_dmem_n10052, MEM_stage_inst_dmem_n10053, MEM_stage_inst_dmem_n10054, MEM_stage_inst_dmem_n10055, MEM_stage_inst_dmem_n10056, MEM_stage_inst_dmem_n10057, MEM_stage_inst_dmem_n10058, MEM_stage_inst_dmem_n10059, MEM_stage_inst_dmem_n10060, MEM_stage_inst_dmem_n10061, MEM_stage_inst_dmem_n10062, MEM_stage_inst_dmem_n10063, MEM_stage_inst_dmem_n10064, MEM_stage_inst_dmem_n10065, MEM_stage_inst_dmem_n10066, MEM_stage_inst_dmem_n10067, MEM_stage_inst_dmem_n10068, MEM_stage_inst_dmem_n10069, MEM_stage_inst_dmem_n10070, MEM_stage_inst_dmem_n10071, MEM_stage_inst_dmem_n10072, MEM_stage_inst_dmem_n10073, MEM_stage_inst_dmem_n10074, MEM_stage_inst_dmem_n10075, MEM_stage_inst_dmem_n10076, MEM_stage_inst_dmem_n10077, MEM_stage_inst_dmem_n10078, MEM_stage_inst_dmem_n10079, MEM_stage_inst_dmem_n10080, MEM_stage_inst_dmem_n10081, MEM_stage_inst_dmem_n10082, MEM_stage_inst_dmem_n10083, MEM_stage_inst_dmem_n10084, MEM_stage_inst_dmem_n10085, MEM_stage_inst_dmem_n10086, MEM_stage_inst_dmem_n10087, MEM_stage_inst_dmem_n10088, MEM_stage_inst_dmem_n10089, MEM_stage_inst_dmem_n10090, MEM_stage_inst_dmem_n10091, MEM_stage_inst_dmem_n10092, MEM_stage_inst_dmem_n10093, MEM_stage_inst_dmem_n10094, MEM_stage_inst_dmem_n10095, MEM_stage_inst_dmem_n10096, MEM_stage_inst_dmem_n10097, MEM_stage_inst_dmem_n10098, MEM_stage_inst_dmem_n10099, MEM_stage_inst_dmem_n10100, MEM_stage_inst_dmem_n10101, MEM_stage_inst_dmem_n10102, MEM_stage_inst_dmem_n10103, MEM_stage_inst_dmem_n10104, MEM_stage_inst_dmem_n10105, MEM_stage_inst_dmem_n10106, MEM_stage_inst_dmem_n10107, MEM_stage_inst_dmem_n10108, MEM_stage_inst_dmem_n10109, MEM_stage_inst_dmem_n10110, MEM_stage_inst_dmem_n10111, MEM_stage_inst_dmem_n10112, MEM_stage_inst_dmem_n10113, MEM_stage_inst_dmem_n10114, MEM_stage_inst_dmem_n10115, MEM_stage_inst_dmem_n10116, MEM_stage_inst_dmem_n10117, MEM_stage_inst_dmem_n10118, MEM_stage_inst_dmem_n10119, MEM_stage_inst_dmem_n10120, MEM_stage_inst_dmem_n10121, MEM_stage_inst_dmem_n10122, MEM_stage_inst_dmem_n10123, MEM_stage_inst_dmem_n10124, MEM_stage_inst_dmem_n10125, MEM_stage_inst_dmem_n10126, MEM_stage_inst_dmem_n10127, MEM_stage_inst_dmem_n10128, MEM_stage_inst_dmem_n10129, MEM_stage_inst_dmem_n10130, MEM_stage_inst_dmem_n10131, MEM_stage_inst_dmem_n10132, MEM_stage_inst_dmem_n10133, MEM_stage_inst_dmem_n10134, MEM_stage_inst_dmem_n10135, MEM_stage_inst_dmem_n10136, MEM_stage_inst_dmem_n10137, MEM_stage_inst_dmem_n10138, MEM_stage_inst_dmem_n10139, MEM_stage_inst_dmem_n10140, MEM_stage_inst_dmem_n10141, MEM_stage_inst_dmem_n10142, MEM_stage_inst_dmem_n10143, MEM_stage_inst_dmem_n10144, MEM_stage_inst_dmem_n10145, MEM_stage_inst_dmem_n10146, MEM_stage_inst_dmem_n10147, MEM_stage_inst_dmem_n10148, MEM_stage_inst_dmem_n10149, MEM_stage_inst_dmem_n10150, MEM_stage_inst_dmem_n10151, MEM_stage_inst_dmem_n10152, MEM_stage_inst_dmem_n10153, MEM_stage_inst_dmem_n10154, MEM_stage_inst_dmem_n10155, MEM_stage_inst_dmem_n10156, MEM_stage_inst_dmem_n10157, MEM_stage_inst_dmem_n10158, MEM_stage_inst_dmem_n10159, MEM_stage_inst_dmem_n10160, MEM_stage_inst_dmem_n10161, MEM_stage_inst_dmem_n10162, MEM_stage_inst_dmem_n10163, MEM_stage_inst_dmem_n10164, MEM_stage_inst_dmem_n10165, MEM_stage_inst_dmem_n10166, MEM_stage_inst_dmem_n10167, MEM_stage_inst_dmem_n10168, MEM_stage_inst_dmem_n10169, MEM_stage_inst_dmem_n10170, MEM_stage_inst_dmem_n10171, MEM_stage_inst_dmem_n10172, MEM_stage_inst_dmem_n10173, MEM_stage_inst_dmem_n10174, MEM_stage_inst_dmem_n10175, MEM_stage_inst_dmem_n10176, MEM_stage_inst_dmem_n10177, MEM_stage_inst_dmem_n10178, MEM_stage_inst_dmem_n10179, MEM_stage_inst_dmem_n10180, MEM_stage_inst_dmem_n10181, MEM_stage_inst_dmem_n10182, MEM_stage_inst_dmem_n10183, MEM_stage_inst_dmem_n10184, MEM_stage_inst_dmem_n10185, MEM_stage_inst_dmem_n10186, MEM_stage_inst_dmem_n10187, MEM_stage_inst_dmem_n10188, MEM_stage_inst_dmem_n10189, MEM_stage_inst_dmem_n10190, MEM_stage_inst_dmem_n10191, MEM_stage_inst_dmem_n10192, MEM_stage_inst_dmem_n10193, MEM_stage_inst_dmem_n10194, MEM_stage_inst_dmem_n10195, MEM_stage_inst_dmem_n10196, MEM_stage_inst_dmem_n10197, MEM_stage_inst_dmem_n10198, MEM_stage_inst_dmem_n10199, MEM_stage_inst_dmem_n10200, MEM_stage_inst_dmem_n10201, MEM_stage_inst_dmem_n10202, MEM_stage_inst_dmem_n10203, MEM_stage_inst_dmem_n10204, MEM_stage_inst_dmem_n10205, MEM_stage_inst_dmem_n10206, MEM_stage_inst_dmem_n10207, MEM_stage_inst_dmem_n10208, MEM_stage_inst_dmem_n10209, MEM_stage_inst_dmem_n10210, MEM_stage_inst_dmem_n10211, MEM_stage_inst_dmem_n10212, MEM_stage_inst_dmem_n10213, MEM_stage_inst_dmem_n10214, MEM_stage_inst_dmem_n10215, MEM_stage_inst_dmem_n10216, MEM_stage_inst_dmem_n10217, MEM_stage_inst_dmem_n10218, MEM_stage_inst_dmem_n10219, MEM_stage_inst_dmem_n10220, MEM_stage_inst_dmem_n10221, MEM_stage_inst_dmem_n10222, MEM_stage_inst_dmem_n10223, MEM_stage_inst_dmem_n10224, MEM_stage_inst_dmem_n10225, MEM_stage_inst_dmem_n10226, MEM_stage_inst_dmem_n10227, MEM_stage_inst_dmem_n10228, MEM_stage_inst_dmem_n10229, MEM_stage_inst_dmem_n10230, MEM_stage_inst_dmem_n10231, MEM_stage_inst_dmem_n10232, MEM_stage_inst_dmem_n10233, MEM_stage_inst_dmem_n10234, MEM_stage_inst_dmem_n10235, MEM_stage_inst_dmem_n10236, MEM_stage_inst_dmem_n10237, MEM_stage_inst_dmem_n10238, MEM_stage_inst_dmem_n10239, MEM_stage_inst_dmem_n10240, MEM_stage_inst_dmem_n10241, MEM_stage_inst_dmem_n10242, MEM_stage_inst_dmem_n10243, MEM_stage_inst_dmem_n10244, MEM_stage_inst_dmem_n10245, MEM_stage_inst_dmem_n10246, MEM_stage_inst_dmem_n10247, MEM_stage_inst_dmem_n10248, MEM_stage_inst_dmem_n10249, MEM_stage_inst_dmem_n10250, MEM_stage_inst_dmem_n10251, MEM_stage_inst_dmem_n10252, MEM_stage_inst_dmem_n10253, MEM_stage_inst_dmem_n10254, MEM_stage_inst_dmem_n10255, MEM_stage_inst_dmem_n10256, MEM_stage_inst_dmem_n10257, MEM_stage_inst_dmem_n10258, MEM_stage_inst_dmem_n10259, MEM_stage_inst_dmem_n10260, MEM_stage_inst_dmem_n10261, MEM_stage_inst_dmem_n10262, MEM_stage_inst_dmem_n10263, MEM_stage_inst_dmem_n10264, MEM_stage_inst_dmem_n10265, MEM_stage_inst_dmem_n10266, MEM_stage_inst_dmem_n10267, MEM_stage_inst_dmem_n10268, MEM_stage_inst_dmem_n10269, MEM_stage_inst_dmem_n10270, MEM_stage_inst_dmem_n10271, MEM_stage_inst_dmem_n10272, MEM_stage_inst_dmem_n10273, MEM_stage_inst_dmem_n10274, MEM_stage_inst_dmem_n10275, MEM_stage_inst_dmem_n10276, MEM_stage_inst_dmem_n10277, MEM_stage_inst_dmem_n10278, MEM_stage_inst_dmem_n10279, MEM_stage_inst_dmem_n10280, MEM_stage_inst_dmem_n10281, MEM_stage_inst_dmem_n10282, MEM_stage_inst_dmem_n10283, MEM_stage_inst_dmem_n10284, MEM_stage_inst_dmem_n10285, MEM_stage_inst_dmem_n10286, MEM_stage_inst_dmem_n10287, MEM_stage_inst_dmem_n10288, MEM_stage_inst_dmem_n10289, MEM_stage_inst_dmem_n10290, MEM_stage_inst_dmem_n10291, MEM_stage_inst_dmem_n10292, MEM_stage_inst_dmem_n10293, MEM_stage_inst_dmem_n10294, MEM_stage_inst_dmem_n10295, MEM_stage_inst_dmem_n10296, MEM_stage_inst_dmem_n10297, MEM_stage_inst_dmem_n10298, MEM_stage_inst_dmem_n10299, MEM_stage_inst_dmem_n10300, MEM_stage_inst_dmem_n10301, MEM_stage_inst_dmem_n10302, MEM_stage_inst_dmem_n10303, MEM_stage_inst_dmem_n10304, MEM_stage_inst_dmem_n10305, MEM_stage_inst_dmem_n10306, MEM_stage_inst_dmem_n10307, MEM_stage_inst_dmem_n10308, MEM_stage_inst_dmem_n10309, MEM_stage_inst_dmem_n10310, MEM_stage_inst_dmem_n10311, MEM_stage_inst_dmem_n10312, MEM_stage_inst_dmem_n10313, MEM_stage_inst_dmem_n10314, MEM_stage_inst_dmem_n10315, MEM_stage_inst_dmem_n10316, MEM_stage_inst_dmem_n10317, MEM_stage_inst_dmem_n10318, MEM_stage_inst_dmem_n10319, MEM_stage_inst_dmem_n10320, MEM_stage_inst_dmem_n10321, MEM_stage_inst_dmem_n10322, MEM_stage_inst_dmem_n10323, MEM_stage_inst_dmem_n10324, MEM_stage_inst_dmem_n10325, MEM_stage_inst_dmem_n10326, MEM_stage_inst_dmem_n10327, MEM_stage_inst_dmem_n10328, MEM_stage_inst_dmem_n10329, MEM_stage_inst_dmem_n10330, MEM_stage_inst_dmem_n10331, MEM_stage_inst_dmem_n10332, MEM_stage_inst_dmem_n10333, MEM_stage_inst_dmem_n10334, MEM_stage_inst_dmem_n10335, MEM_stage_inst_dmem_n10336, MEM_stage_inst_dmem_n10337, MEM_stage_inst_dmem_n10338, MEM_stage_inst_dmem_n10339, MEM_stage_inst_dmem_n10340, MEM_stage_inst_dmem_n10341, MEM_stage_inst_dmem_n10342, MEM_stage_inst_dmem_n10343, MEM_stage_inst_dmem_n10344, MEM_stage_inst_dmem_n10345, MEM_stage_inst_dmem_n10346, MEM_stage_inst_dmem_n10347, MEM_stage_inst_dmem_n10348, MEM_stage_inst_dmem_n10349, MEM_stage_inst_dmem_n10350, MEM_stage_inst_dmem_n10351, MEM_stage_inst_dmem_n10352, MEM_stage_inst_dmem_n10353, MEM_stage_inst_dmem_n10354, MEM_stage_inst_dmem_n10355, MEM_stage_inst_dmem_n10356, MEM_stage_inst_dmem_n10357, MEM_stage_inst_dmem_n10358, MEM_stage_inst_dmem_n10359, MEM_stage_inst_dmem_n10360, MEM_stage_inst_dmem_n10361, MEM_stage_inst_dmem_n10362, MEM_stage_inst_dmem_n10363, MEM_stage_inst_dmem_n10364, MEM_stage_inst_dmem_n10365, MEM_stage_inst_dmem_n10366, MEM_stage_inst_dmem_n10367, MEM_stage_inst_dmem_n10368, MEM_stage_inst_dmem_n10369, MEM_stage_inst_dmem_n10370, MEM_stage_inst_dmem_n10371, MEM_stage_inst_dmem_n10372, MEM_stage_inst_dmem_n10373, MEM_stage_inst_dmem_n10374, MEM_stage_inst_dmem_n10375, MEM_stage_inst_dmem_n10376, MEM_stage_inst_dmem_n10377, MEM_stage_inst_dmem_n10378, MEM_stage_inst_dmem_n10379, MEM_stage_inst_dmem_n10380, MEM_stage_inst_dmem_n10381, MEM_stage_inst_dmem_n10382, MEM_stage_inst_dmem_n10383, MEM_stage_inst_dmem_n10384, MEM_stage_inst_dmem_n10385, MEM_stage_inst_dmem_n10386, MEM_stage_inst_dmem_n10387, MEM_stage_inst_dmem_n10388, MEM_stage_inst_dmem_n10389, MEM_stage_inst_dmem_n10390, MEM_stage_inst_dmem_n10391, MEM_stage_inst_dmem_n10392, MEM_stage_inst_dmem_n10393, MEM_stage_inst_dmem_n10394, MEM_stage_inst_dmem_n10395, MEM_stage_inst_dmem_n10396, MEM_stage_inst_dmem_n10397, MEM_stage_inst_dmem_n10398, MEM_stage_inst_dmem_n10399, MEM_stage_inst_dmem_n10400, MEM_stage_inst_dmem_n10401, MEM_stage_inst_dmem_n10402, MEM_stage_inst_dmem_n10403, MEM_stage_inst_dmem_n10404, MEM_stage_inst_dmem_n10405, MEM_stage_inst_dmem_n10406, MEM_stage_inst_dmem_n10407, MEM_stage_inst_dmem_n10408, MEM_stage_inst_dmem_n10409, MEM_stage_inst_dmem_n10410, MEM_stage_inst_dmem_n10411, MEM_stage_inst_dmem_n10412, MEM_stage_inst_dmem_n10413, MEM_stage_inst_dmem_n10414, MEM_stage_inst_dmem_n10415, MEM_stage_inst_dmem_n10416, MEM_stage_inst_dmem_n10417, MEM_stage_inst_dmem_n10418, MEM_stage_inst_dmem_n10419, MEM_stage_inst_dmem_n10420, MEM_stage_inst_dmem_n10421, MEM_stage_inst_dmem_n10422, MEM_stage_inst_dmem_n10423, MEM_stage_inst_dmem_n10424, MEM_stage_inst_dmem_n10425, MEM_stage_inst_dmem_n10426, MEM_stage_inst_dmem_n10427, MEM_stage_inst_dmem_n10428, MEM_stage_inst_dmem_n10429, MEM_stage_inst_dmem_n10430, MEM_stage_inst_dmem_n10431, MEM_stage_inst_dmem_n10432, MEM_stage_inst_dmem_n10433, MEM_stage_inst_dmem_n10434, MEM_stage_inst_dmem_n10435, MEM_stage_inst_dmem_n10436, MEM_stage_inst_dmem_n10437, MEM_stage_inst_dmem_n10438, MEM_stage_inst_dmem_n10439, MEM_stage_inst_dmem_n10440, MEM_stage_inst_dmem_n10441, MEM_stage_inst_dmem_n10442, MEM_stage_inst_dmem_n10443, MEM_stage_inst_dmem_n10444, MEM_stage_inst_dmem_n10445, MEM_stage_inst_dmem_n10446, MEM_stage_inst_dmem_n10447, MEM_stage_inst_dmem_n10448, MEM_stage_inst_dmem_n10449, MEM_stage_inst_dmem_n10450, MEM_stage_inst_dmem_n10451, MEM_stage_inst_dmem_n10452, MEM_stage_inst_dmem_n10453, MEM_stage_inst_dmem_n10454, MEM_stage_inst_dmem_n10455, MEM_stage_inst_dmem_n10456, MEM_stage_inst_dmem_n10457, MEM_stage_inst_dmem_n10458, MEM_stage_inst_dmem_n10459, MEM_stage_inst_dmem_n10460, MEM_stage_inst_dmem_n10461, MEM_stage_inst_dmem_n10462, MEM_stage_inst_dmem_n10463, MEM_stage_inst_dmem_n10464, MEM_stage_inst_dmem_n10465, MEM_stage_inst_dmem_n10466, MEM_stage_inst_dmem_n10467, MEM_stage_inst_dmem_n10468, MEM_stage_inst_dmem_n10469, MEM_stage_inst_dmem_n10470, MEM_stage_inst_dmem_n10471, MEM_stage_inst_dmem_n10472, MEM_stage_inst_dmem_n10473, MEM_stage_inst_dmem_n10474, MEM_stage_inst_dmem_n10475, MEM_stage_inst_dmem_n10476, MEM_stage_inst_dmem_n10477, MEM_stage_inst_dmem_n10478, MEM_stage_inst_dmem_n10479, MEM_stage_inst_dmem_n10480, MEM_stage_inst_dmem_n10481, MEM_stage_inst_dmem_n10482, MEM_stage_inst_dmem_n10483, MEM_stage_inst_dmem_n10484, MEM_stage_inst_dmem_n10485, MEM_stage_inst_dmem_n10486, MEM_stage_inst_dmem_n10487, MEM_stage_inst_dmem_n10488, MEM_stage_inst_dmem_n10489, MEM_stage_inst_dmem_n10490, MEM_stage_inst_dmem_n10491, MEM_stage_inst_dmem_n10492, MEM_stage_inst_dmem_n10493, MEM_stage_inst_dmem_n10494, MEM_stage_inst_dmem_n10495, MEM_stage_inst_dmem_n10496, MEM_stage_inst_dmem_n10497, MEM_stage_inst_dmem_n10498, MEM_stage_inst_dmem_n10499, MEM_stage_inst_dmem_n10500, MEM_stage_inst_dmem_n10501, MEM_stage_inst_dmem_n10502, MEM_stage_inst_dmem_n10503, MEM_stage_inst_dmem_n10504, MEM_stage_inst_dmem_n10505, MEM_stage_inst_dmem_n10506, MEM_stage_inst_dmem_n10507, MEM_stage_inst_dmem_n10508, MEM_stage_inst_dmem_n10509, MEM_stage_inst_dmem_n10510, MEM_stage_inst_dmem_n10511, MEM_stage_inst_dmem_n10512, MEM_stage_inst_dmem_n10513, MEM_stage_inst_dmem_n10514, MEM_stage_inst_dmem_n10515, MEM_stage_inst_dmem_n10516, MEM_stage_inst_dmem_n10517, MEM_stage_inst_dmem_n10518, MEM_stage_inst_dmem_n10519, MEM_stage_inst_dmem_n10520, MEM_stage_inst_dmem_n10521, MEM_stage_inst_dmem_n10522, MEM_stage_inst_dmem_n10523, MEM_stage_inst_dmem_n10524, MEM_stage_inst_dmem_n10525, MEM_stage_inst_dmem_n10526, MEM_stage_inst_dmem_n10527, MEM_stage_inst_dmem_n10528, MEM_stage_inst_dmem_n10529, MEM_stage_inst_dmem_n10530, MEM_stage_inst_dmem_n10531, MEM_stage_inst_dmem_n10532, MEM_stage_inst_dmem_n10533, MEM_stage_inst_dmem_n10534, MEM_stage_inst_dmem_n10535, MEM_stage_inst_dmem_n10536, MEM_stage_inst_dmem_n10537, MEM_stage_inst_dmem_n10538, MEM_stage_inst_dmem_n10539, MEM_stage_inst_dmem_n10540, MEM_stage_inst_dmem_n10541, MEM_stage_inst_dmem_n10542, MEM_stage_inst_dmem_n10543, MEM_stage_inst_dmem_n10544, MEM_stage_inst_dmem_n10545, MEM_stage_inst_dmem_n10546, MEM_stage_inst_dmem_n10547, MEM_stage_inst_dmem_n10548, MEM_stage_inst_dmem_n10549, MEM_stage_inst_dmem_n10550, MEM_stage_inst_dmem_n10551, MEM_stage_inst_dmem_n10552, MEM_stage_inst_dmem_n10553, MEM_stage_inst_dmem_n10554, MEM_stage_inst_dmem_n10555, MEM_stage_inst_dmem_n10556, MEM_stage_inst_dmem_n10557, MEM_stage_inst_dmem_n10558, MEM_stage_inst_dmem_n10559, MEM_stage_inst_dmem_n10560, MEM_stage_inst_dmem_n10561, MEM_stage_inst_dmem_n10562, MEM_stage_inst_dmem_n10563, MEM_stage_inst_dmem_n10564, MEM_stage_inst_dmem_n10565, MEM_stage_inst_dmem_n10566, MEM_stage_inst_dmem_n10567, MEM_stage_inst_dmem_n10568, MEM_stage_inst_dmem_n10569, MEM_stage_inst_dmem_n10570, MEM_stage_inst_dmem_n10571, MEM_stage_inst_dmem_n10572, MEM_stage_inst_dmem_n10573, MEM_stage_inst_dmem_n10574, MEM_stage_inst_dmem_n10575, MEM_stage_inst_dmem_n10576, MEM_stage_inst_dmem_n10577, MEM_stage_inst_dmem_n10578, MEM_stage_inst_dmem_n10579, MEM_stage_inst_dmem_n10580, MEM_stage_inst_dmem_n10581, MEM_stage_inst_dmem_n10582, MEM_stage_inst_dmem_n10583, MEM_stage_inst_dmem_n10584, MEM_stage_inst_dmem_n10585, MEM_stage_inst_dmem_n10586, MEM_stage_inst_dmem_n10587, MEM_stage_inst_dmem_n10588, MEM_stage_inst_dmem_n10589, MEM_stage_inst_dmem_n10590, MEM_stage_inst_dmem_n10591, MEM_stage_inst_dmem_n10592, MEM_stage_inst_dmem_n10593, MEM_stage_inst_dmem_n10594, MEM_stage_inst_dmem_n10595, MEM_stage_inst_dmem_n10596, MEM_stage_inst_dmem_n10597, MEM_stage_inst_dmem_n10598, MEM_stage_inst_dmem_n10599, MEM_stage_inst_dmem_n10600, MEM_stage_inst_dmem_n10601, MEM_stage_inst_dmem_n10602, MEM_stage_inst_dmem_n10603, MEM_stage_inst_dmem_n10604, MEM_stage_inst_dmem_n10605, MEM_stage_inst_dmem_n10606, MEM_stage_inst_dmem_n10607, MEM_stage_inst_dmem_n10608, MEM_stage_inst_dmem_n10609, MEM_stage_inst_dmem_n10610, MEM_stage_inst_dmem_n10611, MEM_stage_inst_dmem_n10612, MEM_stage_inst_dmem_n10613, MEM_stage_inst_dmem_n10614, MEM_stage_inst_dmem_n10615, MEM_stage_inst_dmem_n10616, MEM_stage_inst_dmem_n10617, MEM_stage_inst_dmem_n10618, MEM_stage_inst_dmem_n10619, MEM_stage_inst_dmem_n10620, MEM_stage_inst_dmem_n10621, MEM_stage_inst_dmem_n10622, MEM_stage_inst_dmem_n10623, MEM_stage_inst_dmem_n10624, MEM_stage_inst_dmem_n10625, MEM_stage_inst_dmem_n10626, MEM_stage_inst_dmem_n10627, MEM_stage_inst_dmem_n10628, MEM_stage_inst_dmem_n10629, MEM_stage_inst_dmem_n10630, MEM_stage_inst_dmem_n10631, MEM_stage_inst_dmem_n10632, MEM_stage_inst_dmem_n10633, MEM_stage_inst_dmem_n10634, MEM_stage_inst_dmem_n10635, MEM_stage_inst_dmem_n10636, MEM_stage_inst_dmem_n10637, MEM_stage_inst_dmem_n10638, MEM_stage_inst_dmem_n10639, MEM_stage_inst_dmem_n10640, MEM_stage_inst_dmem_n10641, MEM_stage_inst_dmem_n10642, MEM_stage_inst_dmem_n10643, MEM_stage_inst_dmem_n10644, MEM_stage_inst_dmem_n10645, MEM_stage_inst_dmem_n10646, MEM_stage_inst_dmem_n10647, MEM_stage_inst_dmem_n10648, MEM_stage_inst_dmem_n10649, MEM_stage_inst_dmem_n10650, MEM_stage_inst_dmem_n10651, MEM_stage_inst_dmem_n10652, MEM_stage_inst_dmem_n10653, MEM_stage_inst_dmem_n10654, MEM_stage_inst_dmem_n10655, MEM_stage_inst_dmem_n10656, MEM_stage_inst_dmem_n10657, MEM_stage_inst_dmem_n10658, MEM_stage_inst_dmem_n10659, MEM_stage_inst_dmem_n10660, MEM_stage_inst_dmem_n10661, MEM_stage_inst_dmem_n10662, MEM_stage_inst_dmem_n10663, MEM_stage_inst_dmem_n10664, MEM_stage_inst_dmem_n10665, MEM_stage_inst_dmem_n10666, MEM_stage_inst_dmem_n10667, MEM_stage_inst_dmem_n10668, MEM_stage_inst_dmem_n10669, MEM_stage_inst_dmem_n10670, MEM_stage_inst_dmem_n10671, MEM_stage_inst_dmem_n10672, MEM_stage_inst_dmem_n10673, MEM_stage_inst_dmem_n10674, MEM_stage_inst_dmem_n10675, MEM_stage_inst_dmem_n10676, MEM_stage_inst_dmem_n10677, MEM_stage_inst_dmem_n10678, MEM_stage_inst_dmem_n10679, MEM_stage_inst_dmem_n10680, MEM_stage_inst_dmem_n10681, MEM_stage_inst_dmem_n10682, MEM_stage_inst_dmem_n10683, MEM_stage_inst_dmem_n10684, MEM_stage_inst_dmem_n10685, MEM_stage_inst_dmem_n10686, MEM_stage_inst_dmem_n10687, MEM_stage_inst_dmem_n10688, MEM_stage_inst_dmem_n10689, MEM_stage_inst_dmem_n10690, MEM_stage_inst_dmem_n10691, MEM_stage_inst_dmem_n10692, MEM_stage_inst_dmem_n10693, MEM_stage_inst_dmem_n10694, MEM_stage_inst_dmem_n10695, MEM_stage_inst_dmem_n10696, MEM_stage_inst_dmem_n10697, MEM_stage_inst_dmem_n10698, MEM_stage_inst_dmem_n10699, MEM_stage_inst_dmem_n10700, MEM_stage_inst_dmem_n10701, MEM_stage_inst_dmem_n10702, MEM_stage_inst_dmem_n10703, MEM_stage_inst_dmem_n10704, MEM_stage_inst_dmem_n10705, MEM_stage_inst_dmem_n10706, MEM_stage_inst_dmem_n10707, MEM_stage_inst_dmem_n10708, MEM_stage_inst_dmem_n10709, MEM_stage_inst_dmem_n10710, MEM_stage_inst_dmem_n10711, MEM_stage_inst_dmem_n10712, MEM_stage_inst_dmem_n10713, MEM_stage_inst_dmem_n10714, MEM_stage_inst_dmem_n10715, MEM_stage_inst_dmem_n10716, MEM_stage_inst_dmem_n10717, MEM_stage_inst_dmem_n10718, MEM_stage_inst_dmem_n10719, MEM_stage_inst_dmem_n10720, MEM_stage_inst_dmem_n10721, MEM_stage_inst_dmem_n10722, MEM_stage_inst_dmem_n10723, MEM_stage_inst_dmem_n10724, MEM_stage_inst_dmem_n10725, MEM_stage_inst_dmem_n10726, MEM_stage_inst_dmem_n10727, MEM_stage_inst_dmem_n10728, MEM_stage_inst_dmem_n10729, MEM_stage_inst_dmem_n10730, MEM_stage_inst_dmem_n10731, MEM_stage_inst_dmem_n10732, MEM_stage_inst_dmem_n10733, MEM_stage_inst_dmem_n10734, MEM_stage_inst_dmem_n10735, MEM_stage_inst_dmem_n10736, MEM_stage_inst_dmem_n10737, MEM_stage_inst_dmem_n10738, MEM_stage_inst_dmem_n10739, MEM_stage_inst_dmem_n10740, MEM_stage_inst_dmem_n10741, MEM_stage_inst_dmem_n10742, MEM_stage_inst_dmem_n10743, MEM_stage_inst_dmem_n10744, MEM_stage_inst_dmem_n10745, MEM_stage_inst_dmem_n10746, MEM_stage_inst_dmem_n10747, MEM_stage_inst_dmem_n10748, MEM_stage_inst_dmem_n10749, MEM_stage_inst_dmem_n10750, MEM_stage_inst_dmem_n10751, MEM_stage_inst_dmem_n10752, MEM_stage_inst_dmem_n10753, MEM_stage_inst_dmem_n10754, MEM_stage_inst_dmem_n10755, MEM_stage_inst_dmem_n10756, MEM_stage_inst_dmem_n10757, MEM_stage_inst_dmem_n10758, MEM_stage_inst_dmem_n10759, MEM_stage_inst_dmem_n10760, MEM_stage_inst_dmem_n10761, MEM_stage_inst_dmem_n10762, MEM_stage_inst_dmem_n10763, MEM_stage_inst_dmem_n10764, MEM_stage_inst_dmem_n10765, MEM_stage_inst_dmem_n10766, MEM_stage_inst_dmem_n10767, MEM_stage_inst_dmem_n10768, MEM_stage_inst_dmem_n10769, MEM_stage_inst_dmem_n10770, MEM_stage_inst_dmem_n10771, MEM_stage_inst_dmem_n10772, MEM_stage_inst_dmem_n10773, MEM_stage_inst_dmem_n10774, MEM_stage_inst_dmem_n10775, MEM_stage_inst_dmem_n10776, MEM_stage_inst_dmem_n10777, MEM_stage_inst_dmem_n10778, MEM_stage_inst_dmem_n10779, MEM_stage_inst_dmem_n10780, MEM_stage_inst_dmem_n10781, MEM_stage_inst_dmem_n10782, MEM_stage_inst_dmem_n10783, MEM_stage_inst_dmem_n10784, MEM_stage_inst_dmem_n10785, MEM_stage_inst_dmem_n10786, MEM_stage_inst_dmem_n10787, MEM_stage_inst_dmem_n10788, MEM_stage_inst_dmem_n10789, MEM_stage_inst_dmem_n10790, MEM_stage_inst_dmem_n10791, MEM_stage_inst_dmem_n10792, MEM_stage_inst_dmem_n10793, MEM_stage_inst_dmem_n10794, MEM_stage_inst_dmem_n10795, MEM_stage_inst_dmem_n10796, MEM_stage_inst_dmem_n10797, MEM_stage_inst_dmem_n10798, MEM_stage_inst_dmem_n10799, MEM_stage_inst_dmem_n10800, MEM_stage_inst_dmem_n10801, MEM_stage_inst_dmem_n10802, MEM_stage_inst_dmem_n10803, MEM_stage_inst_dmem_n10804, MEM_stage_inst_dmem_n10805, MEM_stage_inst_dmem_n10806, MEM_stage_inst_dmem_n10807, MEM_stage_inst_dmem_n10808, MEM_stage_inst_dmem_n10809, MEM_stage_inst_dmem_n10810, MEM_stage_inst_dmem_n10811, MEM_stage_inst_dmem_n10812, MEM_stage_inst_dmem_n10813, MEM_stage_inst_dmem_n10814, MEM_stage_inst_dmem_n10815, MEM_stage_inst_dmem_n10816, MEM_stage_inst_dmem_n10817, MEM_stage_inst_dmem_n10818, MEM_stage_inst_dmem_n10819, MEM_stage_inst_dmem_n10820, MEM_stage_inst_dmem_n10821, MEM_stage_inst_dmem_n10822, MEM_stage_inst_dmem_n10823, MEM_stage_inst_dmem_n10824, MEM_stage_inst_dmem_n10825, MEM_stage_inst_dmem_n10826, MEM_stage_inst_dmem_n10827, MEM_stage_inst_dmem_n10828, MEM_stage_inst_dmem_n10829, MEM_stage_inst_dmem_n10830, MEM_stage_inst_dmem_n10831, MEM_stage_inst_dmem_n10832, MEM_stage_inst_dmem_n10833, MEM_stage_inst_dmem_n10834, MEM_stage_inst_dmem_n10835, MEM_stage_inst_dmem_n10836, MEM_stage_inst_dmem_n10837, MEM_stage_inst_dmem_n10838, MEM_stage_inst_dmem_n10839, MEM_stage_inst_dmem_n10840, MEM_stage_inst_dmem_n10841, MEM_stage_inst_dmem_n10842, MEM_stage_inst_dmem_n10843, MEM_stage_inst_dmem_n10844, MEM_stage_inst_dmem_n10845, MEM_stage_inst_dmem_n10846, MEM_stage_inst_dmem_n10847, MEM_stage_inst_dmem_n10848, MEM_stage_inst_dmem_n10849, MEM_stage_inst_dmem_n10850, MEM_stage_inst_dmem_n10851, MEM_stage_inst_dmem_n10852, MEM_stage_inst_dmem_n10853, MEM_stage_inst_dmem_n10854, MEM_stage_inst_dmem_n10855, MEM_stage_inst_dmem_n10856, MEM_stage_inst_dmem_n10857, MEM_stage_inst_dmem_n10858, MEM_stage_inst_dmem_n10859, MEM_stage_inst_dmem_n10860, MEM_stage_inst_dmem_n10861, MEM_stage_inst_dmem_n10862, MEM_stage_inst_dmem_n10863, MEM_stage_inst_dmem_n10864, MEM_stage_inst_dmem_n10865, MEM_stage_inst_dmem_n10866, MEM_stage_inst_dmem_n10867, MEM_stage_inst_dmem_n10868, MEM_stage_inst_dmem_n10869, MEM_stage_inst_dmem_n10870, MEM_stage_inst_dmem_n10871, MEM_stage_inst_dmem_n10872, MEM_stage_inst_dmem_n10873, MEM_stage_inst_dmem_n10874, MEM_stage_inst_dmem_n10875, MEM_stage_inst_dmem_n10876, MEM_stage_inst_dmem_n10877, MEM_stage_inst_dmem_n10878, MEM_stage_inst_dmem_n10879, MEM_stage_inst_dmem_n10880, MEM_stage_inst_dmem_n10881, MEM_stage_inst_dmem_n10882, MEM_stage_inst_dmem_n10883, MEM_stage_inst_dmem_n10884, MEM_stage_inst_dmem_n10885, MEM_stage_inst_dmem_n10886, MEM_stage_inst_dmem_n10887, MEM_stage_inst_dmem_n10888, MEM_stage_inst_dmem_n10889, MEM_stage_inst_dmem_n10890, MEM_stage_inst_dmem_n10891, MEM_stage_inst_dmem_n10892, MEM_stage_inst_dmem_n10893, MEM_stage_inst_dmem_n10894, MEM_stage_inst_dmem_n10895, MEM_stage_inst_dmem_n10896, MEM_stage_inst_dmem_n10897, MEM_stage_inst_dmem_n10898, MEM_stage_inst_dmem_n10899, MEM_stage_inst_dmem_n10900, MEM_stage_inst_dmem_n10901, MEM_stage_inst_dmem_n10902, MEM_stage_inst_dmem_n10903, MEM_stage_inst_dmem_n10904, MEM_stage_inst_dmem_n10905, MEM_stage_inst_dmem_n10906, MEM_stage_inst_dmem_n10907, MEM_stage_inst_dmem_n10908, MEM_stage_inst_dmem_n10909, MEM_stage_inst_dmem_n10910, MEM_stage_inst_dmem_n10911, MEM_stage_inst_dmem_n10912, MEM_stage_inst_dmem_n10913, MEM_stage_inst_dmem_n10914, MEM_stage_inst_dmem_n10915, MEM_stage_inst_dmem_n10916, MEM_stage_inst_dmem_n10917, MEM_stage_inst_dmem_n10918, MEM_stage_inst_dmem_n10919, MEM_stage_inst_dmem_n10920, MEM_stage_inst_dmem_n10921, MEM_stage_inst_dmem_n10922, MEM_stage_inst_dmem_n10923, MEM_stage_inst_dmem_n10924, MEM_stage_inst_dmem_n10925, MEM_stage_inst_dmem_n10926, MEM_stage_inst_dmem_n10927, MEM_stage_inst_dmem_n10928, MEM_stage_inst_dmem_n10929, MEM_stage_inst_dmem_n10930, MEM_stage_inst_dmem_n10931, MEM_stage_inst_dmem_n10932, MEM_stage_inst_dmem_n10933, MEM_stage_inst_dmem_n10934, MEM_stage_inst_dmem_n10935, MEM_stage_inst_dmem_n10936, MEM_stage_inst_dmem_n10937, MEM_stage_inst_dmem_n10938, MEM_stage_inst_dmem_n10939, MEM_stage_inst_dmem_n10940, MEM_stage_inst_dmem_n10941, MEM_stage_inst_dmem_n10942, MEM_stage_inst_dmem_n10943, MEM_stage_inst_dmem_n10944, MEM_stage_inst_dmem_n10945, MEM_stage_inst_dmem_n10946, MEM_stage_inst_dmem_n10947, MEM_stage_inst_dmem_n10948, MEM_stage_inst_dmem_n10949, MEM_stage_inst_dmem_n10950, MEM_stage_inst_dmem_n10951, MEM_stage_inst_dmem_n10952, MEM_stage_inst_dmem_n10953, MEM_stage_inst_dmem_n10954, MEM_stage_inst_dmem_n10955, MEM_stage_inst_dmem_n10956, MEM_stage_inst_dmem_n10957, MEM_stage_inst_dmem_n10958, MEM_stage_inst_dmem_n10959, MEM_stage_inst_dmem_n10960, MEM_stage_inst_dmem_n10961, MEM_stage_inst_dmem_n10962, MEM_stage_inst_dmem_n10963, MEM_stage_inst_dmem_n10964, MEM_stage_inst_dmem_n10965, MEM_stage_inst_dmem_n10966, MEM_stage_inst_dmem_n10967, MEM_stage_inst_dmem_n10968, MEM_stage_inst_dmem_n10969, MEM_stage_inst_dmem_n10970, MEM_stage_inst_dmem_n10971, MEM_stage_inst_dmem_n10972, MEM_stage_inst_dmem_n10973, MEM_stage_inst_dmem_n10974, MEM_stage_inst_dmem_n10975, MEM_stage_inst_dmem_n10976, MEM_stage_inst_dmem_n10977, MEM_stage_inst_dmem_n10978, MEM_stage_inst_dmem_n10979, MEM_stage_inst_dmem_n10980, MEM_stage_inst_dmem_n10981, MEM_stage_inst_dmem_n10982, MEM_stage_inst_dmem_n10983, MEM_stage_inst_dmem_n10984, MEM_stage_inst_dmem_n10985, MEM_stage_inst_dmem_n10986, MEM_stage_inst_dmem_n10987, MEM_stage_inst_dmem_n10988, MEM_stage_inst_dmem_n10989, MEM_stage_inst_dmem_n10990, MEM_stage_inst_dmem_n10991, MEM_stage_inst_dmem_n10992, MEM_stage_inst_dmem_n10993, MEM_stage_inst_dmem_n10994, MEM_stage_inst_dmem_n10995, MEM_stage_inst_dmem_n10996, MEM_stage_inst_dmem_n10997, MEM_stage_inst_dmem_n10998, MEM_stage_inst_dmem_n10999, MEM_stage_inst_dmem_n11000, MEM_stage_inst_dmem_n11001, MEM_stage_inst_dmem_n11002, MEM_stage_inst_dmem_n11003, MEM_stage_inst_dmem_n11004, MEM_stage_inst_dmem_n11005, MEM_stage_inst_dmem_n11006, MEM_stage_inst_dmem_n11007, MEM_stage_inst_dmem_n11008, MEM_stage_inst_dmem_n11009, MEM_stage_inst_dmem_n11010, MEM_stage_inst_dmem_n11011, MEM_stage_inst_dmem_n11012, MEM_stage_inst_dmem_n11013, MEM_stage_inst_dmem_n11014, MEM_stage_inst_dmem_n11015, MEM_stage_inst_dmem_n11016, MEM_stage_inst_dmem_n11017, MEM_stage_inst_dmem_n11018, MEM_stage_inst_dmem_n11019, MEM_stage_inst_dmem_n11020, MEM_stage_inst_dmem_n11021, MEM_stage_inst_dmem_n11022, MEM_stage_inst_dmem_n11023, MEM_stage_inst_dmem_n11024, MEM_stage_inst_dmem_n11025, MEM_stage_inst_dmem_n11026, MEM_stage_inst_dmem_n11027, MEM_stage_inst_dmem_n11028, MEM_stage_inst_dmem_n11029, MEM_stage_inst_dmem_n11030, MEM_stage_inst_dmem_n11031, MEM_stage_inst_dmem_n11032, MEM_stage_inst_dmem_n11033, MEM_stage_inst_dmem_n11034, MEM_stage_inst_dmem_n11035, MEM_stage_inst_dmem_n11036, MEM_stage_inst_dmem_n11037, MEM_stage_inst_dmem_n11038, MEM_stage_inst_dmem_n11039, MEM_stage_inst_dmem_n11040, MEM_stage_inst_dmem_n11041, MEM_stage_inst_dmem_n11042, MEM_stage_inst_dmem_n11043, MEM_stage_inst_dmem_n11044, MEM_stage_inst_dmem_n11045, MEM_stage_inst_dmem_n11046, MEM_stage_inst_dmem_n11047, MEM_stage_inst_dmem_n11048, MEM_stage_inst_dmem_n11049, MEM_stage_inst_dmem_n11050, MEM_stage_inst_dmem_n11051, MEM_stage_inst_dmem_n11052, MEM_stage_inst_dmem_n11053, MEM_stage_inst_dmem_n11054, MEM_stage_inst_dmem_n11055, MEM_stage_inst_dmem_n11056, MEM_stage_inst_dmem_n11057, MEM_stage_inst_dmem_n11058, MEM_stage_inst_dmem_n11059, MEM_stage_inst_dmem_n11060, MEM_stage_inst_dmem_n11061, MEM_stage_inst_dmem_n11062, MEM_stage_inst_dmem_n11063, MEM_stage_inst_dmem_n11064, MEM_stage_inst_dmem_n11065, MEM_stage_inst_dmem_n11066, MEM_stage_inst_dmem_n11067, MEM_stage_inst_dmem_n11068, MEM_stage_inst_dmem_n11069, MEM_stage_inst_dmem_n11070, MEM_stage_inst_dmem_n11071, MEM_stage_inst_dmem_n11072, MEM_stage_inst_dmem_n11073, MEM_stage_inst_dmem_n11074, MEM_stage_inst_dmem_n11075, MEM_stage_inst_dmem_n11076, MEM_stage_inst_dmem_n11077, MEM_stage_inst_dmem_n11078, MEM_stage_inst_dmem_n11079, MEM_stage_inst_dmem_n11080, MEM_stage_inst_dmem_n11081, MEM_stage_inst_dmem_n11082, MEM_stage_inst_dmem_n11083, MEM_stage_inst_dmem_n11084, MEM_stage_inst_dmem_n11085, MEM_stage_inst_dmem_n11086, MEM_stage_inst_dmem_n11087, MEM_stage_inst_dmem_n11088, MEM_stage_inst_dmem_n11089, MEM_stage_inst_dmem_n11090, MEM_stage_inst_dmem_n11091, MEM_stage_inst_dmem_n11092, MEM_stage_inst_dmem_n11093, MEM_stage_inst_dmem_n11094, MEM_stage_inst_dmem_n11095, MEM_stage_inst_dmem_n11096, MEM_stage_inst_dmem_n11097, MEM_stage_inst_dmem_n11098, MEM_stage_inst_dmem_n11099, MEM_stage_inst_dmem_n11100, MEM_stage_inst_dmem_n11101, MEM_stage_inst_dmem_n11102, MEM_stage_inst_dmem_n11103, MEM_stage_inst_dmem_n11104, MEM_stage_inst_dmem_n11105, MEM_stage_inst_dmem_n11106, MEM_stage_inst_dmem_n11107, MEM_stage_inst_dmem_n11108, MEM_stage_inst_dmem_n11109, MEM_stage_inst_dmem_n11110, MEM_stage_inst_dmem_n11111, MEM_stage_inst_dmem_n11112, MEM_stage_inst_dmem_n11113, MEM_stage_inst_dmem_n11114, MEM_stage_inst_dmem_n11115, MEM_stage_inst_dmem_n11116, MEM_stage_inst_dmem_n11117, MEM_stage_inst_dmem_n11118, MEM_stage_inst_dmem_n11119, MEM_stage_inst_dmem_n11120, MEM_stage_inst_dmem_n11121, MEM_stage_inst_dmem_n11122, MEM_stage_inst_dmem_n11123, MEM_stage_inst_dmem_n11124, MEM_stage_inst_dmem_n11125, MEM_stage_inst_dmem_n11126, MEM_stage_inst_dmem_n11127, MEM_stage_inst_dmem_n11128, MEM_stage_inst_dmem_n11129, MEM_stage_inst_dmem_n11130, MEM_stage_inst_dmem_n11131, MEM_stage_inst_dmem_n11132, MEM_stage_inst_dmem_n11133, MEM_stage_inst_dmem_n11134, MEM_stage_inst_dmem_n11135, MEM_stage_inst_dmem_n11136, MEM_stage_inst_dmem_n11137, MEM_stage_inst_dmem_n11138, MEM_stage_inst_dmem_n11139, MEM_stage_inst_dmem_n11140, MEM_stage_inst_dmem_n11141, MEM_stage_inst_dmem_n11142, MEM_stage_inst_dmem_n11143, MEM_stage_inst_dmem_n11144, MEM_stage_inst_dmem_n11145, MEM_stage_inst_dmem_n11146, MEM_stage_inst_dmem_n11147, MEM_stage_inst_dmem_n11148, MEM_stage_inst_dmem_n11149, MEM_stage_inst_dmem_n11150, MEM_stage_inst_dmem_n11151, MEM_stage_inst_dmem_n11152, MEM_stage_inst_dmem_n11153, MEM_stage_inst_dmem_n11154, MEM_stage_inst_dmem_n11155, MEM_stage_inst_dmem_n11156, MEM_stage_inst_dmem_n11157, MEM_stage_inst_dmem_n11158, MEM_stage_inst_dmem_n11159, MEM_stage_inst_dmem_n11160, MEM_stage_inst_dmem_n11161, MEM_stage_inst_dmem_n11162, MEM_stage_inst_dmem_n11163, MEM_stage_inst_dmem_n11164, MEM_stage_inst_dmem_n11165, MEM_stage_inst_dmem_n11166, MEM_stage_inst_dmem_n11167, MEM_stage_inst_dmem_n11168, MEM_stage_inst_dmem_n11169, MEM_stage_inst_dmem_n11170, MEM_stage_inst_dmem_n11171, MEM_stage_inst_dmem_n11172, MEM_stage_inst_dmem_n11173, MEM_stage_inst_dmem_n11174, MEM_stage_inst_dmem_n11175, MEM_stage_inst_dmem_n11176, MEM_stage_inst_dmem_n11177, MEM_stage_inst_dmem_n11178, MEM_stage_inst_dmem_n11179, MEM_stage_inst_dmem_n11180, MEM_stage_inst_dmem_n11181, MEM_stage_inst_dmem_n11182, MEM_stage_inst_dmem_n11183, MEM_stage_inst_dmem_n11184, MEM_stage_inst_dmem_n11185, MEM_stage_inst_dmem_n11186, MEM_stage_inst_dmem_n11187, MEM_stage_inst_dmem_n11188, MEM_stage_inst_dmem_n11189, MEM_stage_inst_dmem_n11190, MEM_stage_inst_dmem_n11191, MEM_stage_inst_dmem_n11192, MEM_stage_inst_dmem_n11193, MEM_stage_inst_dmem_n11194, MEM_stage_inst_dmem_n11195, MEM_stage_inst_dmem_n11196, MEM_stage_inst_dmem_n11197, MEM_stage_inst_dmem_n11198, MEM_stage_inst_dmem_n11199, MEM_stage_inst_dmem_n11200, MEM_stage_inst_dmem_n11201, MEM_stage_inst_dmem_n11202, MEM_stage_inst_dmem_n11203, MEM_stage_inst_dmem_n11204, MEM_stage_inst_dmem_n11205, MEM_stage_inst_dmem_n11206, MEM_stage_inst_dmem_n11207, MEM_stage_inst_dmem_n11208, MEM_stage_inst_dmem_n11209, MEM_stage_inst_dmem_n11210, MEM_stage_inst_dmem_n11211, MEM_stage_inst_dmem_n11212, MEM_stage_inst_dmem_n11213, MEM_stage_inst_dmem_n11214, MEM_stage_inst_dmem_n11215, MEM_stage_inst_dmem_n11216, MEM_stage_inst_dmem_n11217, MEM_stage_inst_dmem_n11218, MEM_stage_inst_dmem_n11219, MEM_stage_inst_dmem_n11220, MEM_stage_inst_dmem_n11221, MEM_stage_inst_dmem_n11222, MEM_stage_inst_dmem_n11223, MEM_stage_inst_dmem_n11224, MEM_stage_inst_dmem_n11225, MEM_stage_inst_dmem_n11226, MEM_stage_inst_dmem_n11227, MEM_stage_inst_dmem_n11228, MEM_stage_inst_dmem_n11229, MEM_stage_inst_dmem_n11230, MEM_stage_inst_dmem_n11231, MEM_stage_inst_dmem_n11232, MEM_stage_inst_dmem_n11233, MEM_stage_inst_dmem_n11234, MEM_stage_inst_dmem_n11235, MEM_stage_inst_dmem_n11236, MEM_stage_inst_dmem_n11237, MEM_stage_inst_dmem_n11238, MEM_stage_inst_dmem_n11239, MEM_stage_inst_dmem_n11240, MEM_stage_inst_dmem_n11241, MEM_stage_inst_dmem_n11242, MEM_stage_inst_dmem_n11243, MEM_stage_inst_dmem_n11244, MEM_stage_inst_dmem_n11245, MEM_stage_inst_dmem_n11246, MEM_stage_inst_dmem_n11247, MEM_stage_inst_dmem_n11248, MEM_stage_inst_dmem_n11249, MEM_stage_inst_dmem_n11250, MEM_stage_inst_dmem_n11251, MEM_stage_inst_dmem_n11252, MEM_stage_inst_dmem_n11253, MEM_stage_inst_dmem_n11254, MEM_stage_inst_dmem_n11255, MEM_stage_inst_dmem_n11256, MEM_stage_inst_dmem_n11257, MEM_stage_inst_dmem_n11258, MEM_stage_inst_dmem_n11259, MEM_stage_inst_dmem_n11260, MEM_stage_inst_dmem_n11261, MEM_stage_inst_dmem_n11262, MEM_stage_inst_dmem_n11263, MEM_stage_inst_dmem_n11264, MEM_stage_inst_dmem_n11265, MEM_stage_inst_dmem_n11266, MEM_stage_inst_dmem_n11267, MEM_stage_inst_dmem_n11268, MEM_stage_inst_dmem_n11269, MEM_stage_inst_dmem_n11270, MEM_stage_inst_dmem_n11271, MEM_stage_inst_dmem_n11272, MEM_stage_inst_dmem_n11273, MEM_stage_inst_dmem_n11274, MEM_stage_inst_dmem_n11275, MEM_stage_inst_dmem_n11276, MEM_stage_inst_dmem_n11277, MEM_stage_inst_dmem_n11278, MEM_stage_inst_dmem_n11279, MEM_stage_inst_dmem_n11280, MEM_stage_inst_dmem_n11281, MEM_stage_inst_dmem_n11282, MEM_stage_inst_dmem_n11283, MEM_stage_inst_dmem_n11284, MEM_stage_inst_dmem_n11285, MEM_stage_inst_dmem_n11286, MEM_stage_inst_dmem_n11287, MEM_stage_inst_dmem_n11288, MEM_stage_inst_dmem_n11289, MEM_stage_inst_dmem_n11290, MEM_stage_inst_dmem_n11291, MEM_stage_inst_dmem_n11292, MEM_stage_inst_dmem_n11293, MEM_stage_inst_dmem_n11294, MEM_stage_inst_dmem_n11295, MEM_stage_inst_dmem_n11296, MEM_stage_inst_dmem_n11297, MEM_stage_inst_dmem_n11298, MEM_stage_inst_dmem_n11299, MEM_stage_inst_dmem_n11300, MEM_stage_inst_dmem_n11301, MEM_stage_inst_dmem_n11302, MEM_stage_inst_dmem_n11303, MEM_stage_inst_dmem_n11304, MEM_stage_inst_dmem_n11305, MEM_stage_inst_dmem_n11306, MEM_stage_inst_dmem_n11307, MEM_stage_inst_dmem_n11308, MEM_stage_inst_dmem_n11309, MEM_stage_inst_dmem_n11310, MEM_stage_inst_dmem_n11311, MEM_stage_inst_dmem_n11312, MEM_stage_inst_dmem_n11313, MEM_stage_inst_dmem_n11314, MEM_stage_inst_dmem_n11315, MEM_stage_inst_dmem_n11316, MEM_stage_inst_dmem_n11317, MEM_stage_inst_dmem_n11318, MEM_stage_inst_dmem_n11319, MEM_stage_inst_dmem_n11320, MEM_stage_inst_dmem_n11321, MEM_stage_inst_dmem_n11322, MEM_stage_inst_dmem_n11323, MEM_stage_inst_dmem_n11324, MEM_stage_inst_dmem_n11325, MEM_stage_inst_dmem_n11326, MEM_stage_inst_dmem_n11327, MEM_stage_inst_dmem_n11328, MEM_stage_inst_dmem_n11329, MEM_stage_inst_dmem_n11330, MEM_stage_inst_dmem_n11331, MEM_stage_inst_dmem_n11332, MEM_stage_inst_dmem_n11333, MEM_stage_inst_dmem_n11334, MEM_stage_inst_dmem_n11335, MEM_stage_inst_dmem_n11336, MEM_stage_inst_dmem_n11337, MEM_stage_inst_dmem_n11338, MEM_stage_inst_dmem_n11339, MEM_stage_inst_dmem_n11340, MEM_stage_inst_dmem_n11341, MEM_stage_inst_dmem_n11342, MEM_stage_inst_dmem_n11343, MEM_stage_inst_dmem_n11344, MEM_stage_inst_dmem_n11345, MEM_stage_inst_dmem_n11346, MEM_stage_inst_dmem_n11347, MEM_stage_inst_dmem_n11348, MEM_stage_inst_dmem_n11349, MEM_stage_inst_dmem_n11350, MEM_stage_inst_dmem_n11351, MEM_stage_inst_dmem_n11352, MEM_stage_inst_dmem_n11353, MEM_stage_inst_dmem_n11354, MEM_stage_inst_dmem_n11355, MEM_stage_inst_dmem_n11356, MEM_stage_inst_dmem_n11357, MEM_stage_inst_dmem_n11358, MEM_stage_inst_dmem_n11359, MEM_stage_inst_dmem_n11360, MEM_stage_inst_dmem_n11361, MEM_stage_inst_dmem_n11362, MEM_stage_inst_dmem_n11363, MEM_stage_inst_dmem_n11364, MEM_stage_inst_dmem_n11365, MEM_stage_inst_dmem_n11366, MEM_stage_inst_dmem_n11367, MEM_stage_inst_dmem_n11368, MEM_stage_inst_dmem_n11369, MEM_stage_inst_dmem_n11370, MEM_stage_inst_dmem_n11371, MEM_stage_inst_dmem_n11372, MEM_stage_inst_dmem_n11373, MEM_stage_inst_dmem_n11374, MEM_stage_inst_dmem_n11375, MEM_stage_inst_dmem_n11376, MEM_stage_inst_dmem_n11377, MEM_stage_inst_dmem_n11378, MEM_stage_inst_dmem_n11379, MEM_stage_inst_dmem_n11380, MEM_stage_inst_dmem_n11381, MEM_stage_inst_dmem_n11382, MEM_stage_inst_dmem_n11383, MEM_stage_inst_dmem_n11384, MEM_stage_inst_dmem_n11385, MEM_stage_inst_dmem_n11386, MEM_stage_inst_dmem_n11387, MEM_stage_inst_dmem_n11388, MEM_stage_inst_dmem_n11389, MEM_stage_inst_dmem_n11390, MEM_stage_inst_dmem_n11391, MEM_stage_inst_dmem_n11392, MEM_stage_inst_dmem_n11393, MEM_stage_inst_dmem_n11394, MEM_stage_inst_dmem_n11395, MEM_stage_inst_dmem_n11396, MEM_stage_inst_dmem_n11397, MEM_stage_inst_dmem_n11398, MEM_stage_inst_dmem_n11399, MEM_stage_inst_dmem_n11400, MEM_stage_inst_dmem_n11401, MEM_stage_inst_dmem_n11402, MEM_stage_inst_dmem_n11403, MEM_stage_inst_dmem_n11404, MEM_stage_inst_dmem_n11405, MEM_stage_inst_dmem_n11406, MEM_stage_inst_dmem_n11407, MEM_stage_inst_dmem_n11408, MEM_stage_inst_dmem_n11409, MEM_stage_inst_dmem_n11410, MEM_stage_inst_dmem_n11411, MEM_stage_inst_dmem_n11412, MEM_stage_inst_dmem_n11413, MEM_stage_inst_dmem_n11414, MEM_stage_inst_dmem_n11415, MEM_stage_inst_dmem_n11416, MEM_stage_inst_dmem_n11417, MEM_stage_inst_dmem_n11418, MEM_stage_inst_dmem_n11419, MEM_stage_inst_dmem_n11420, MEM_stage_inst_dmem_n11421, MEM_stage_inst_dmem_n11422, MEM_stage_inst_dmem_n11423, MEM_stage_inst_dmem_n11424, MEM_stage_inst_dmem_n11425, MEM_stage_inst_dmem_n11426, MEM_stage_inst_dmem_n11427, MEM_stage_inst_dmem_n11428, MEM_stage_inst_dmem_n11429, MEM_stage_inst_dmem_n11430, MEM_stage_inst_dmem_n11431, MEM_stage_inst_dmem_n11432, MEM_stage_inst_dmem_n11433, MEM_stage_inst_dmem_n11434, MEM_stage_inst_dmem_n11435, MEM_stage_inst_dmem_n11436, MEM_stage_inst_dmem_n11437, MEM_stage_inst_dmem_n11438, MEM_stage_inst_dmem_n11439, MEM_stage_inst_dmem_n11440, MEM_stage_inst_dmem_n11441, MEM_stage_inst_dmem_n11442, MEM_stage_inst_dmem_n11443, MEM_stage_inst_dmem_n11444, MEM_stage_inst_dmem_n11445, MEM_stage_inst_dmem_n11446, MEM_stage_inst_dmem_n11447, MEM_stage_inst_dmem_n11448, MEM_stage_inst_dmem_n11449, MEM_stage_inst_dmem_n11450, MEM_stage_inst_dmem_n11451, MEM_stage_inst_dmem_n11452, MEM_stage_inst_dmem_n11453, MEM_stage_inst_dmem_n11454, MEM_stage_inst_dmem_n11455, MEM_stage_inst_dmem_n11456, MEM_stage_inst_dmem_n11457, MEM_stage_inst_dmem_n11458, MEM_stage_inst_dmem_n11459, MEM_stage_inst_dmem_n11460, MEM_stage_inst_dmem_n11461, MEM_stage_inst_dmem_n11462, MEM_stage_inst_dmem_n11463, MEM_stage_inst_dmem_n11464, MEM_stage_inst_dmem_n11465, MEM_stage_inst_dmem_n11466, MEM_stage_inst_dmem_n11467, MEM_stage_inst_dmem_n11468, MEM_stage_inst_dmem_n11469, MEM_stage_inst_dmem_n11470, MEM_stage_inst_dmem_n11471, MEM_stage_inst_dmem_n11472, MEM_stage_inst_dmem_n11473, MEM_stage_inst_dmem_n11474, MEM_stage_inst_dmem_n11475, MEM_stage_inst_dmem_n11476, MEM_stage_inst_dmem_n11477, MEM_stage_inst_dmem_n11478, MEM_stage_inst_dmem_n11479, MEM_stage_inst_dmem_n11480, MEM_stage_inst_dmem_n11481, MEM_stage_inst_dmem_n11482, MEM_stage_inst_dmem_n11483, MEM_stage_inst_dmem_n11484, MEM_stage_inst_dmem_n11485, MEM_stage_inst_dmem_n11486, MEM_stage_inst_dmem_n11487, MEM_stage_inst_dmem_n11488, MEM_stage_inst_dmem_n11489, MEM_stage_inst_dmem_n11490, MEM_stage_inst_dmem_n11491, MEM_stage_inst_dmem_n11492, MEM_stage_inst_dmem_n11493, MEM_stage_inst_dmem_n11494, MEM_stage_inst_dmem_n11495, MEM_stage_inst_dmem_n11496, MEM_stage_inst_dmem_n11497, MEM_stage_inst_dmem_n11498, MEM_stage_inst_dmem_n11499, MEM_stage_inst_dmem_n11500, MEM_stage_inst_dmem_n11501, MEM_stage_inst_dmem_n11502, MEM_stage_inst_dmem_n11503, MEM_stage_inst_dmem_n11504, MEM_stage_inst_dmem_n11505, MEM_stage_inst_dmem_n11506, MEM_stage_inst_dmem_n11507, MEM_stage_inst_dmem_n11508, MEM_stage_inst_dmem_n11509, MEM_stage_inst_dmem_n11510, MEM_stage_inst_dmem_n11511, MEM_stage_inst_dmem_n11512, MEM_stage_inst_dmem_n11513, MEM_stage_inst_dmem_n11514, MEM_stage_inst_dmem_n11515, MEM_stage_inst_dmem_n11516, MEM_stage_inst_dmem_n11517, MEM_stage_inst_dmem_n11518, MEM_stage_inst_dmem_n11519, MEM_stage_inst_dmem_n11520, MEM_stage_inst_dmem_n11521, MEM_stage_inst_dmem_n11522, MEM_stage_inst_dmem_n11523, MEM_stage_inst_dmem_n11524, MEM_stage_inst_dmem_n11525, MEM_stage_inst_dmem_n11526, MEM_stage_inst_dmem_n11527, MEM_stage_inst_dmem_n11528, MEM_stage_inst_dmem_n11529, MEM_stage_inst_dmem_n11530, MEM_stage_inst_dmem_n11531, MEM_stage_inst_dmem_n11532, MEM_stage_inst_dmem_n11533, MEM_stage_inst_dmem_n11534, MEM_stage_inst_dmem_n11535, MEM_stage_inst_dmem_n11536, MEM_stage_inst_dmem_n11537, MEM_stage_inst_dmem_n11538, MEM_stage_inst_dmem_n11539, MEM_stage_inst_dmem_n11540, MEM_stage_inst_dmem_n11541, MEM_stage_inst_dmem_n11542, MEM_stage_inst_dmem_n11543, MEM_stage_inst_dmem_n11544, MEM_stage_inst_dmem_n11545, MEM_stage_inst_dmem_n11546, MEM_stage_inst_dmem_n11547, MEM_stage_inst_dmem_n11548, MEM_stage_inst_dmem_n11549, MEM_stage_inst_dmem_n11550, MEM_stage_inst_dmem_n11551, MEM_stage_inst_dmem_n11552, MEM_stage_inst_dmem_n11553, MEM_stage_inst_dmem_n11554, MEM_stage_inst_dmem_n11555, MEM_stage_inst_dmem_n11556, MEM_stage_inst_dmem_n11557, MEM_stage_inst_dmem_n11558, MEM_stage_inst_dmem_n11559, MEM_stage_inst_dmem_n11560, MEM_stage_inst_dmem_n11561, MEM_stage_inst_dmem_n11562, MEM_stage_inst_dmem_n11563, MEM_stage_inst_dmem_n11564, MEM_stage_inst_dmem_n11565, MEM_stage_inst_dmem_n11566, MEM_stage_inst_dmem_n11567, MEM_stage_inst_dmem_n11568, MEM_stage_inst_dmem_n11569, MEM_stage_inst_dmem_n11570, MEM_stage_inst_dmem_n11571, MEM_stage_inst_dmem_n11572, MEM_stage_inst_dmem_n11573, MEM_stage_inst_dmem_n11574, MEM_stage_inst_dmem_n11575, MEM_stage_inst_dmem_n11576, MEM_stage_inst_dmem_n11577, MEM_stage_inst_dmem_n11578, MEM_stage_inst_dmem_n11579, MEM_stage_inst_dmem_n11580, MEM_stage_inst_dmem_n11581, MEM_stage_inst_dmem_n11582, MEM_stage_inst_dmem_n11583, MEM_stage_inst_dmem_n11584, MEM_stage_inst_dmem_n11585, MEM_stage_inst_dmem_n11586, MEM_stage_inst_dmem_n11587, MEM_stage_inst_dmem_n11588, MEM_stage_inst_dmem_n11589, MEM_stage_inst_dmem_n11590, MEM_stage_inst_dmem_n11591, MEM_stage_inst_dmem_n11592, MEM_stage_inst_dmem_n11593, MEM_stage_inst_dmem_n11594, MEM_stage_inst_dmem_n11595, MEM_stage_inst_dmem_n11596, MEM_stage_inst_dmem_n11597, MEM_stage_inst_dmem_n11598, MEM_stage_inst_dmem_n11599, MEM_stage_inst_dmem_n11600, MEM_stage_inst_dmem_n11601, MEM_stage_inst_dmem_n11602, MEM_stage_inst_dmem_n11603, MEM_stage_inst_dmem_n11604, MEM_stage_inst_dmem_n11605, MEM_stage_inst_dmem_n11606, MEM_stage_inst_dmem_n11607, MEM_stage_inst_dmem_n11608, MEM_stage_inst_dmem_n11609, MEM_stage_inst_dmem_n11610, MEM_stage_inst_dmem_n11611, MEM_stage_inst_dmem_n11612, MEM_stage_inst_dmem_n11613, MEM_stage_inst_dmem_n11614, MEM_stage_inst_dmem_n11615, MEM_stage_inst_dmem_n11616, MEM_stage_inst_dmem_n11617, MEM_stage_inst_dmem_n11618, MEM_stage_inst_dmem_n11619, MEM_stage_inst_dmem_n11620, MEM_stage_inst_dmem_n11621, MEM_stage_inst_dmem_n11622, MEM_stage_inst_dmem_n11623, MEM_stage_inst_dmem_n11624, MEM_stage_inst_dmem_n11625, MEM_stage_inst_dmem_n11626, MEM_stage_inst_dmem_n11627, MEM_stage_inst_dmem_n11628, MEM_stage_inst_dmem_n11629, MEM_stage_inst_dmem_n11630, MEM_stage_inst_dmem_n11631, MEM_stage_inst_dmem_n11632, MEM_stage_inst_dmem_n11633, MEM_stage_inst_dmem_n11634, MEM_stage_inst_dmem_n11635, MEM_stage_inst_dmem_n11636, MEM_stage_inst_dmem_n11637, MEM_stage_inst_dmem_n11638, MEM_stage_inst_dmem_n11639, MEM_stage_inst_dmem_n11640, MEM_stage_inst_dmem_n11641, MEM_stage_inst_dmem_n11642, MEM_stage_inst_dmem_n11643, MEM_stage_inst_dmem_n11644, MEM_stage_inst_dmem_n11645, MEM_stage_inst_dmem_n11646, MEM_stage_inst_dmem_n11647, MEM_stage_inst_dmem_n11648, MEM_stage_inst_dmem_n11649, MEM_stage_inst_dmem_n11650, MEM_stage_inst_dmem_n11651, MEM_stage_inst_dmem_n11652, MEM_stage_inst_dmem_n11653, MEM_stage_inst_dmem_n11654, MEM_stage_inst_dmem_n11655, MEM_stage_inst_dmem_n11656, MEM_stage_inst_dmem_n11657, MEM_stage_inst_dmem_n11658, MEM_stage_inst_dmem_n11659, MEM_stage_inst_dmem_n11660, MEM_stage_inst_dmem_n11661, MEM_stage_inst_dmem_n11662, MEM_stage_inst_dmem_n11663, MEM_stage_inst_dmem_n11664, MEM_stage_inst_dmem_n11665, MEM_stage_inst_dmem_n11666, MEM_stage_inst_dmem_n11667, MEM_stage_inst_dmem_n11668, MEM_stage_inst_dmem_n11669, MEM_stage_inst_dmem_n11670, MEM_stage_inst_dmem_n11671, MEM_stage_inst_dmem_n11672, MEM_stage_inst_dmem_n11673, MEM_stage_inst_dmem_n11674, MEM_stage_inst_dmem_n11675, MEM_stage_inst_dmem_n11676, MEM_stage_inst_dmem_n11677, MEM_stage_inst_dmem_n11678, MEM_stage_inst_dmem_n11679, MEM_stage_inst_dmem_n11680, MEM_stage_inst_dmem_n11681, MEM_stage_inst_dmem_n11682, MEM_stage_inst_dmem_n11683, MEM_stage_inst_dmem_n11684, MEM_stage_inst_dmem_n11685, MEM_stage_inst_dmem_n11686, MEM_stage_inst_dmem_n11687, MEM_stage_inst_dmem_n11688, MEM_stage_inst_dmem_n11689, MEM_stage_inst_dmem_n11690, MEM_stage_inst_dmem_n11691, MEM_stage_inst_dmem_n11692, MEM_stage_inst_dmem_n11693, MEM_stage_inst_dmem_n11694, MEM_stage_inst_dmem_n11695, MEM_stage_inst_dmem_n11696, MEM_stage_inst_dmem_n11697, MEM_stage_inst_dmem_n11698, MEM_stage_inst_dmem_n11699, MEM_stage_inst_dmem_n11700, MEM_stage_inst_dmem_n11701, MEM_stage_inst_dmem_n11702, MEM_stage_inst_dmem_n11703, MEM_stage_inst_dmem_n11704, MEM_stage_inst_dmem_n11705, MEM_stage_inst_dmem_n11706, MEM_stage_inst_dmem_n11707, MEM_stage_inst_dmem_n11708, MEM_stage_inst_dmem_n11709, MEM_stage_inst_dmem_n11710, MEM_stage_inst_dmem_n11711, MEM_stage_inst_dmem_n11712, MEM_stage_inst_dmem_n11713, MEM_stage_inst_dmem_n11714, MEM_stage_inst_dmem_n11715, MEM_stage_inst_dmem_n11716, MEM_stage_inst_dmem_n11717, MEM_stage_inst_dmem_n11718, MEM_stage_inst_dmem_n11719, MEM_stage_inst_dmem_n11720, MEM_stage_inst_dmem_n11721, MEM_stage_inst_dmem_n11722, MEM_stage_inst_dmem_n11723, MEM_stage_inst_dmem_n11724, MEM_stage_inst_dmem_n11725, MEM_stage_inst_dmem_n11726, MEM_stage_inst_dmem_n11727, MEM_stage_inst_dmem_n11728, MEM_stage_inst_dmem_n11729, MEM_stage_inst_dmem_n11730, MEM_stage_inst_dmem_n11731, MEM_stage_inst_dmem_n11732, MEM_stage_inst_dmem_n11733, MEM_stage_inst_dmem_n11734, MEM_stage_inst_dmem_n11735, MEM_stage_inst_dmem_n11736, MEM_stage_inst_dmem_n11737, MEM_stage_inst_dmem_n11738, MEM_stage_inst_dmem_n11739, MEM_stage_inst_dmem_n11740, MEM_stage_inst_dmem_n11741, MEM_stage_inst_dmem_n11742, MEM_stage_inst_dmem_n11743, MEM_stage_inst_dmem_n11744, MEM_stage_inst_dmem_n11745, MEM_stage_inst_dmem_n11746, MEM_stage_inst_dmem_n11747, MEM_stage_inst_dmem_n11748, MEM_stage_inst_dmem_n11749, MEM_stage_inst_dmem_n11750, MEM_stage_inst_dmem_n11751, MEM_stage_inst_dmem_n11752, MEM_stage_inst_dmem_n11753, MEM_stage_inst_dmem_n11754, MEM_stage_inst_dmem_n11755, MEM_stage_inst_dmem_n11756, MEM_stage_inst_dmem_n11757, MEM_stage_inst_dmem_n11758, MEM_stage_inst_dmem_n11759, MEM_stage_inst_dmem_n11760, MEM_stage_inst_dmem_n11761, MEM_stage_inst_dmem_n11762, MEM_stage_inst_dmem_n11763, MEM_stage_inst_dmem_n11764, MEM_stage_inst_dmem_n11765, MEM_stage_inst_dmem_n11766, MEM_stage_inst_dmem_n11767, MEM_stage_inst_dmem_n11768, MEM_stage_inst_dmem_n11769, MEM_stage_inst_dmem_n11770, MEM_stage_inst_dmem_n11771, MEM_stage_inst_dmem_n11772, MEM_stage_inst_dmem_n11773, MEM_stage_inst_dmem_n11774, MEM_stage_inst_dmem_n11775, MEM_stage_inst_dmem_n11776, MEM_stage_inst_dmem_n11777, MEM_stage_inst_dmem_n11778, MEM_stage_inst_dmem_n11779, MEM_stage_inst_dmem_n11780, MEM_stage_inst_dmem_n11781, MEM_stage_inst_dmem_n11782, MEM_stage_inst_dmem_n11783, MEM_stage_inst_dmem_n11784, MEM_stage_inst_dmem_n11785, MEM_stage_inst_dmem_n11786, MEM_stage_inst_dmem_n11787, MEM_stage_inst_dmem_n11788, MEM_stage_inst_dmem_n11789, MEM_stage_inst_dmem_n11790, MEM_stage_inst_dmem_n11791, MEM_stage_inst_dmem_n11792, MEM_stage_inst_dmem_n11793, MEM_stage_inst_dmem_n11794, MEM_stage_inst_dmem_n11795, MEM_stage_inst_dmem_n11796, MEM_stage_inst_dmem_n11797, MEM_stage_inst_dmem_n11798, MEM_stage_inst_dmem_n11799, MEM_stage_inst_dmem_n11800, MEM_stage_inst_dmem_n11801, MEM_stage_inst_dmem_n11802, MEM_stage_inst_dmem_n11803, MEM_stage_inst_dmem_n11804, MEM_stage_inst_dmem_n11805, MEM_stage_inst_dmem_n11806, MEM_stage_inst_dmem_n11807, MEM_stage_inst_dmem_n11808, MEM_stage_inst_dmem_n11809, MEM_stage_inst_dmem_n11810, MEM_stage_inst_dmem_n11811, MEM_stage_inst_dmem_n11812, MEM_stage_inst_dmem_n11813, MEM_stage_inst_dmem_n11814, MEM_stage_inst_dmem_n11815, MEM_stage_inst_dmem_n11816, MEM_stage_inst_dmem_n11817, MEM_stage_inst_dmem_n11818, MEM_stage_inst_dmem_n11819, MEM_stage_inst_dmem_n11820, MEM_stage_inst_dmem_n11821, MEM_stage_inst_dmem_n11822, MEM_stage_inst_dmem_n11823, MEM_stage_inst_dmem_n11824, MEM_stage_inst_dmem_n11825, MEM_stage_inst_dmem_n11826, MEM_stage_inst_dmem_n11827, MEM_stage_inst_dmem_n11828, MEM_stage_inst_dmem_n11829, MEM_stage_inst_dmem_n11830, MEM_stage_inst_dmem_n11831, MEM_stage_inst_dmem_n11832, MEM_stage_inst_dmem_n11833, MEM_stage_inst_dmem_n11834, MEM_stage_inst_dmem_n11835, MEM_stage_inst_dmem_n11836, MEM_stage_inst_dmem_n11837, MEM_stage_inst_dmem_n11838, MEM_stage_inst_dmem_n11839, MEM_stage_inst_dmem_n11840, MEM_stage_inst_dmem_n11841, MEM_stage_inst_dmem_n11842, MEM_stage_inst_dmem_n11843, MEM_stage_inst_dmem_n11844, MEM_stage_inst_dmem_n11845, MEM_stage_inst_dmem_n11846, MEM_stage_inst_dmem_n11847, MEM_stage_inst_dmem_n11848, MEM_stage_inst_dmem_n11849, MEM_stage_inst_dmem_n11850, MEM_stage_inst_dmem_n11851, MEM_stage_inst_dmem_n11852, MEM_stage_inst_dmem_n11853, MEM_stage_inst_dmem_n11854, MEM_stage_inst_dmem_n11855, MEM_stage_inst_dmem_n11856, MEM_stage_inst_dmem_n11857, MEM_stage_inst_dmem_n11858, MEM_stage_inst_dmem_n11859, MEM_stage_inst_dmem_n11860, MEM_stage_inst_dmem_n11861, MEM_stage_inst_dmem_n11862, MEM_stage_inst_dmem_n11863, MEM_stage_inst_dmem_n11864, MEM_stage_inst_dmem_n11865, MEM_stage_inst_dmem_n11866, MEM_stage_inst_dmem_n11867, MEM_stage_inst_dmem_n11868, MEM_stage_inst_dmem_n11869, MEM_stage_inst_dmem_n11870, MEM_stage_inst_dmem_n11871, MEM_stage_inst_dmem_n11872, MEM_stage_inst_dmem_n11873, MEM_stage_inst_dmem_n11874, MEM_stage_inst_dmem_n11875, MEM_stage_inst_dmem_n11876, MEM_stage_inst_dmem_n11877, MEM_stage_inst_dmem_n11878, MEM_stage_inst_dmem_n11879, MEM_stage_inst_dmem_n11880, MEM_stage_inst_dmem_n11881, MEM_stage_inst_dmem_n11882, MEM_stage_inst_dmem_n11883, MEM_stage_inst_dmem_n11884, MEM_stage_inst_dmem_n11885, MEM_stage_inst_dmem_n11886, MEM_stage_inst_dmem_n11887, MEM_stage_inst_dmem_n11888, MEM_stage_inst_dmem_n11889, MEM_stage_inst_dmem_n11890, MEM_stage_inst_dmem_n11891, MEM_stage_inst_dmem_n11892, MEM_stage_inst_dmem_n11893, MEM_stage_inst_dmem_n11894, MEM_stage_inst_dmem_n11895, MEM_stage_inst_dmem_n11896, MEM_stage_inst_dmem_n11897, MEM_stage_inst_dmem_n11898, MEM_stage_inst_dmem_n11899, MEM_stage_inst_dmem_n11900, MEM_stage_inst_dmem_n11901, MEM_stage_inst_dmem_n11902, MEM_stage_inst_dmem_n11903, MEM_stage_inst_dmem_n11904, MEM_stage_inst_dmem_n11905, MEM_stage_inst_dmem_n11906, MEM_stage_inst_dmem_n11907, MEM_stage_inst_dmem_n11908, MEM_stage_inst_dmem_n11909, MEM_stage_inst_dmem_n11910, MEM_stage_inst_dmem_n11911, MEM_stage_inst_dmem_n11912, MEM_stage_inst_dmem_n11913, MEM_stage_inst_dmem_n11914, MEM_stage_inst_dmem_n11915, MEM_stage_inst_dmem_n11916, MEM_stage_inst_dmem_n11917, MEM_stage_inst_dmem_n11918, MEM_stage_inst_dmem_n11919, MEM_stage_inst_dmem_n11920, MEM_stage_inst_dmem_n11921, MEM_stage_inst_dmem_n11922, MEM_stage_inst_dmem_n11923, MEM_stage_inst_dmem_n11924, MEM_stage_inst_dmem_n11925, MEM_stage_inst_dmem_n11926, MEM_stage_inst_dmem_n11927, MEM_stage_inst_dmem_n11928, MEM_stage_inst_dmem_n11929, MEM_stage_inst_dmem_n11930, MEM_stage_inst_dmem_n11931, MEM_stage_inst_dmem_n11932, MEM_stage_inst_dmem_n11933, MEM_stage_inst_dmem_n11934, MEM_stage_inst_dmem_n11935, MEM_stage_inst_dmem_n11936, MEM_stage_inst_dmem_n11937, MEM_stage_inst_dmem_n11938, MEM_stage_inst_dmem_n11939, MEM_stage_inst_dmem_n11940, MEM_stage_inst_dmem_n11941, MEM_stage_inst_dmem_n11942, MEM_stage_inst_dmem_n11943, MEM_stage_inst_dmem_n11944, MEM_stage_inst_dmem_n11945, MEM_stage_inst_dmem_n11946, MEM_stage_inst_dmem_n11947, MEM_stage_inst_dmem_n11948, MEM_stage_inst_dmem_n11949, MEM_stage_inst_dmem_n11950, MEM_stage_inst_dmem_n11951, MEM_stage_inst_dmem_n11952, MEM_stage_inst_dmem_n11953, MEM_stage_inst_dmem_n11954, MEM_stage_inst_dmem_n11955, MEM_stage_inst_dmem_n11956, MEM_stage_inst_dmem_n11957, MEM_stage_inst_dmem_n11958, MEM_stage_inst_dmem_n11959, MEM_stage_inst_dmem_n11960, MEM_stage_inst_dmem_n11961, MEM_stage_inst_dmem_n11962, MEM_stage_inst_dmem_n11963, MEM_stage_inst_dmem_n11964, MEM_stage_inst_dmem_n11965, MEM_stage_inst_dmem_n11966, MEM_stage_inst_dmem_n11967, MEM_stage_inst_dmem_n11968, MEM_stage_inst_dmem_n11969, MEM_stage_inst_dmem_n11970, MEM_stage_inst_dmem_n11971, MEM_stage_inst_dmem_n11972, MEM_stage_inst_dmem_n11973, MEM_stage_inst_dmem_n11974, MEM_stage_inst_dmem_n11975, MEM_stage_inst_dmem_n11976, MEM_stage_inst_dmem_n11977, MEM_stage_inst_dmem_n11978, MEM_stage_inst_dmem_n11979, MEM_stage_inst_dmem_n11980, MEM_stage_inst_dmem_n11981, MEM_stage_inst_dmem_n11982, MEM_stage_inst_dmem_n11983, MEM_stage_inst_dmem_n11984, MEM_stage_inst_dmem_n11985, MEM_stage_inst_dmem_n11986, MEM_stage_inst_dmem_n11987, MEM_stage_inst_dmem_n11988, MEM_stage_inst_dmem_n11989, MEM_stage_inst_dmem_n11990, MEM_stage_inst_dmem_n11991, MEM_stage_inst_dmem_n11992, MEM_stage_inst_dmem_n11993, MEM_stage_inst_dmem_n11994, MEM_stage_inst_dmem_n11995, MEM_stage_inst_dmem_n11996, MEM_stage_inst_dmem_n11997, MEM_stage_inst_dmem_n11998, MEM_stage_inst_dmem_n11999, MEM_stage_inst_dmem_n12000, MEM_stage_inst_dmem_n12001, MEM_stage_inst_dmem_n12002, MEM_stage_inst_dmem_n12003, MEM_stage_inst_dmem_n12004, MEM_stage_inst_dmem_n12005, MEM_stage_inst_dmem_n12006, MEM_stage_inst_dmem_n12007, MEM_stage_inst_dmem_n12008, MEM_stage_inst_dmem_n12009, MEM_stage_inst_dmem_n12010, MEM_stage_inst_dmem_n12011, MEM_stage_inst_dmem_n12012, MEM_stage_inst_dmem_n12013, MEM_stage_inst_dmem_n12014, MEM_stage_inst_dmem_n12015, MEM_stage_inst_dmem_n12016, MEM_stage_inst_dmem_n12017, MEM_stage_inst_dmem_n12018, MEM_stage_inst_dmem_n12019, MEM_stage_inst_dmem_n12020, MEM_stage_inst_dmem_n12021, MEM_stage_inst_dmem_n12022, MEM_stage_inst_dmem_n12023, MEM_stage_inst_dmem_n12024, MEM_stage_inst_dmem_n12025, MEM_stage_inst_dmem_n12026, MEM_stage_inst_dmem_n12027, MEM_stage_inst_dmem_n12028, MEM_stage_inst_dmem_n12029, MEM_stage_inst_dmem_n12030, MEM_stage_inst_dmem_n12031, MEM_stage_inst_dmem_n12032, MEM_stage_inst_dmem_n12033, MEM_stage_inst_dmem_n12034, MEM_stage_inst_dmem_n12035, MEM_stage_inst_dmem_n12036, MEM_stage_inst_dmem_n12037, MEM_stage_inst_dmem_n12038, MEM_stage_inst_dmem_n12039, MEM_stage_inst_dmem_n12040, MEM_stage_inst_dmem_n12041, MEM_stage_inst_dmem_n12042, MEM_stage_inst_dmem_n12043, MEM_stage_inst_dmem_n12044, MEM_stage_inst_dmem_n12045, MEM_stage_inst_dmem_n12046, MEM_stage_inst_dmem_n12047, MEM_stage_inst_dmem_n12048, MEM_stage_inst_dmem_n12049, MEM_stage_inst_dmem_n12050, MEM_stage_inst_dmem_n12051, MEM_stage_inst_dmem_n12052, MEM_stage_inst_dmem_n12053, MEM_stage_inst_dmem_n12054, MEM_stage_inst_dmem_n12055, MEM_stage_inst_dmem_n12056, MEM_stage_inst_dmem_n12057, MEM_stage_inst_dmem_n12058, MEM_stage_inst_dmem_n12059, MEM_stage_inst_dmem_n12060, MEM_stage_inst_dmem_n12061, MEM_stage_inst_dmem_n12062, MEM_stage_inst_dmem_n12063, MEM_stage_inst_dmem_n12064, MEM_stage_inst_dmem_n12065, MEM_stage_inst_dmem_n12066, MEM_stage_inst_dmem_n12067, MEM_stage_inst_dmem_n12068, MEM_stage_inst_dmem_n12069, MEM_stage_inst_dmem_n12070, MEM_stage_inst_dmem_n12071, MEM_stage_inst_dmem_n12072, MEM_stage_inst_dmem_n12073, MEM_stage_inst_dmem_n12074, MEM_stage_inst_dmem_n12075, MEM_stage_inst_dmem_n12076, MEM_stage_inst_dmem_n12077, MEM_stage_inst_dmem_n12078, MEM_stage_inst_dmem_n12079, MEM_stage_inst_dmem_n12080, MEM_stage_inst_dmem_n12081, MEM_stage_inst_dmem_n12082, MEM_stage_inst_dmem_n12083, MEM_stage_inst_dmem_n12084, MEM_stage_inst_dmem_n12085, MEM_stage_inst_dmem_n12086, MEM_stage_inst_dmem_n12087, MEM_stage_inst_dmem_n12088, MEM_stage_inst_dmem_n12089, MEM_stage_inst_dmem_n12090, MEM_stage_inst_dmem_n12091, MEM_stage_inst_dmem_n12092, MEM_stage_inst_dmem_n12093, MEM_stage_inst_dmem_n12094, MEM_stage_inst_dmem_n12095, MEM_stage_inst_dmem_n12096, MEM_stage_inst_dmem_n12097, MEM_stage_inst_dmem_n12098, MEM_stage_inst_dmem_n12099, MEM_stage_inst_dmem_n12100, MEM_stage_inst_dmem_n12101, MEM_stage_inst_dmem_n12102, MEM_stage_inst_dmem_n12103, MEM_stage_inst_dmem_n12104, MEM_stage_inst_dmem_n12105, MEM_stage_inst_dmem_n12106, MEM_stage_inst_dmem_n12107, MEM_stage_inst_dmem_n12108, MEM_stage_inst_dmem_n12109, MEM_stage_inst_dmem_n12110, MEM_stage_inst_dmem_n12111, MEM_stage_inst_dmem_n12112, MEM_stage_inst_dmem_n12113, MEM_stage_inst_dmem_n12114, MEM_stage_inst_dmem_n12115, MEM_stage_inst_dmem_n12116, MEM_stage_inst_dmem_n12117, MEM_stage_inst_dmem_n12118, MEM_stage_inst_dmem_n12119, MEM_stage_inst_dmem_n12120, MEM_stage_inst_dmem_n12121, MEM_stage_inst_dmem_n12122, MEM_stage_inst_dmem_n12123, MEM_stage_inst_dmem_n12124, MEM_stage_inst_dmem_n12125, MEM_stage_inst_dmem_n12126, MEM_stage_inst_dmem_n12127, MEM_stage_inst_dmem_n12128, MEM_stage_inst_dmem_n12129, MEM_stage_inst_dmem_n12130, MEM_stage_inst_dmem_n12131, MEM_stage_inst_dmem_n12132, MEM_stage_inst_dmem_n12133, MEM_stage_inst_dmem_n12134, MEM_stage_inst_dmem_n12135, MEM_stage_inst_dmem_n12136, MEM_stage_inst_dmem_n12137, MEM_stage_inst_dmem_n12138, MEM_stage_inst_dmem_n12139, MEM_stage_inst_dmem_n12140, MEM_stage_inst_dmem_n12141, MEM_stage_inst_dmem_n12142, MEM_stage_inst_dmem_n12143, MEM_stage_inst_dmem_n12144, MEM_stage_inst_dmem_n12145, MEM_stage_inst_dmem_n12146, MEM_stage_inst_dmem_n12147, MEM_stage_inst_dmem_n12148, MEM_stage_inst_dmem_n12149, MEM_stage_inst_dmem_n12150, MEM_stage_inst_dmem_n12151, MEM_stage_inst_dmem_n12152, MEM_stage_inst_dmem_n12153, MEM_stage_inst_dmem_n12154, MEM_stage_inst_dmem_n12155, MEM_stage_inst_dmem_n12156, MEM_stage_inst_dmem_n12157, MEM_stage_inst_dmem_n12158, MEM_stage_inst_dmem_n12159, MEM_stage_inst_dmem_n12160, MEM_stage_inst_dmem_n12161, MEM_stage_inst_dmem_n12162, MEM_stage_inst_dmem_n12163, MEM_stage_inst_dmem_n12164, MEM_stage_inst_dmem_n12165, MEM_stage_inst_dmem_n12166, MEM_stage_inst_dmem_n12167, MEM_stage_inst_dmem_n12168, MEM_stage_inst_dmem_n12169, MEM_stage_inst_dmem_n12170, MEM_stage_inst_dmem_n12171, MEM_stage_inst_dmem_n12172, MEM_stage_inst_dmem_n12173, MEM_stage_inst_dmem_n12174, MEM_stage_inst_dmem_n12175, MEM_stage_inst_dmem_n12176, MEM_stage_inst_dmem_n12177, MEM_stage_inst_dmem_n12178, MEM_stage_inst_dmem_n12179, MEM_stage_inst_dmem_n12180, MEM_stage_inst_dmem_n12181, MEM_stage_inst_dmem_n12182, MEM_stage_inst_dmem_n12183, MEM_stage_inst_dmem_n12184, MEM_stage_inst_dmem_n12185, MEM_stage_inst_dmem_n12186, MEM_stage_inst_dmem_n12187, MEM_stage_inst_dmem_n12188, MEM_stage_inst_dmem_n12189, MEM_stage_inst_dmem_n12190, MEM_stage_inst_dmem_n12191, MEM_stage_inst_dmem_n12192, MEM_stage_inst_dmem_n12193, MEM_stage_inst_dmem_n12194, MEM_stage_inst_dmem_n12195, MEM_stage_inst_dmem_n12196, MEM_stage_inst_dmem_n12197, MEM_stage_inst_dmem_n12198, MEM_stage_inst_dmem_n12199, MEM_stage_inst_dmem_n12200, MEM_stage_inst_dmem_n12201, MEM_stage_inst_dmem_n12202, MEM_stage_inst_dmem_n12203, MEM_stage_inst_dmem_n12204, MEM_stage_inst_dmem_n12205, MEM_stage_inst_dmem_n12206, MEM_stage_inst_dmem_n12207, MEM_stage_inst_dmem_n12208, MEM_stage_inst_dmem_n12209, MEM_stage_inst_dmem_n12210, MEM_stage_inst_dmem_n12211, MEM_stage_inst_dmem_n12212, MEM_stage_inst_dmem_n12213, MEM_stage_inst_dmem_n12214, MEM_stage_inst_dmem_n12215, MEM_stage_inst_dmem_n12216, MEM_stage_inst_dmem_n12217, MEM_stage_inst_dmem_n12218, MEM_stage_inst_dmem_n12219, MEM_stage_inst_dmem_n12220, MEM_stage_inst_dmem_n12221, MEM_stage_inst_dmem_n12222, MEM_stage_inst_dmem_n12223, MEM_stage_inst_dmem_n12224, MEM_stage_inst_dmem_n12225, MEM_stage_inst_dmem_n12226, MEM_stage_inst_dmem_n12227, MEM_stage_inst_dmem_n12228, MEM_stage_inst_dmem_n12229, MEM_stage_inst_dmem_n12230, MEM_stage_inst_dmem_n12231, MEM_stage_inst_dmem_n12232, MEM_stage_inst_dmem_n12233, MEM_stage_inst_dmem_n12234, MEM_stage_inst_dmem_n12235, MEM_stage_inst_dmem_n12236, MEM_stage_inst_dmem_n12237, MEM_stage_inst_dmem_n12238, MEM_stage_inst_dmem_n12239, MEM_stage_inst_dmem_n12240, MEM_stage_inst_dmem_n12241, MEM_stage_inst_dmem_n12242, MEM_stage_inst_dmem_n12243, MEM_stage_inst_dmem_n12244, MEM_stage_inst_dmem_n12245, MEM_stage_inst_dmem_n12246, MEM_stage_inst_dmem_n12247, MEM_stage_inst_dmem_n12248, MEM_stage_inst_dmem_n12249, MEM_stage_inst_dmem_n12250, MEM_stage_inst_dmem_n12251, MEM_stage_inst_dmem_n12252, MEM_stage_inst_dmem_n12253, MEM_stage_inst_dmem_n12254, MEM_stage_inst_dmem_n12255, MEM_stage_inst_dmem_n12256, MEM_stage_inst_dmem_n12257, MEM_stage_inst_dmem_n12258, MEM_stage_inst_dmem_n12259, MEM_stage_inst_dmem_n12260, MEM_stage_inst_dmem_n12261, MEM_stage_inst_dmem_n12262, MEM_stage_inst_dmem_n12263, MEM_stage_inst_dmem_n12264, MEM_stage_inst_dmem_n12265, MEM_stage_inst_dmem_n12266, MEM_stage_inst_dmem_n12267, MEM_stage_inst_dmem_n12268, MEM_stage_inst_dmem_n12269, MEM_stage_inst_dmem_n12270, MEM_stage_inst_dmem_n12271, MEM_stage_inst_dmem_n12272, MEM_stage_inst_dmem_n12273, MEM_stage_inst_dmem_n12274, MEM_stage_inst_dmem_n12275, MEM_stage_inst_dmem_n12276, MEM_stage_inst_dmem_n12277, MEM_stage_inst_dmem_n12278, MEM_stage_inst_dmem_n12279, MEM_stage_inst_dmem_n12280, MEM_stage_inst_dmem_n12281, MEM_stage_inst_dmem_n12282, MEM_stage_inst_dmem_n12283, MEM_stage_inst_dmem_n12284, MEM_stage_inst_dmem_n12285, MEM_stage_inst_dmem_n12286, MEM_stage_inst_dmem_n12287, MEM_stage_inst_dmem_n12288, MEM_stage_inst_dmem_n12289, MEM_stage_inst_dmem_n12290, MEM_stage_inst_dmem_n12291, MEM_stage_inst_dmem_n12292, MEM_stage_inst_dmem_n12293, MEM_stage_inst_dmem_n12294, MEM_stage_inst_dmem_n12295, MEM_stage_inst_dmem_n12296, MEM_stage_inst_dmem_n12297, MEM_stage_inst_dmem_n12298, MEM_stage_inst_dmem_n12299, MEM_stage_inst_dmem_n12300, MEM_stage_inst_dmem_n12301, MEM_stage_inst_dmem_n12302, MEM_stage_inst_dmem_n12303, MEM_stage_inst_dmem_n12304, MEM_stage_inst_dmem_n12305, MEM_stage_inst_dmem_n12306, MEM_stage_inst_dmem_n12307, MEM_stage_inst_dmem_n12308, MEM_stage_inst_dmem_n12309, MEM_stage_inst_dmem_n12310, MEM_stage_inst_dmem_n12311, MEM_stage_inst_dmem_n12312, MEM_stage_inst_dmem_n12313, MEM_stage_inst_dmem_n12314, MEM_stage_inst_dmem_n12315, MEM_stage_inst_dmem_n12316, MEM_stage_inst_dmem_n12317, MEM_stage_inst_dmem_n12318, MEM_stage_inst_dmem_n12319, MEM_stage_inst_dmem_n12320, MEM_stage_inst_dmem_n12321, MEM_stage_inst_dmem_n12322, MEM_stage_inst_dmem_n12323, MEM_stage_inst_dmem_n12324, MEM_stage_inst_dmem_n12325, MEM_stage_inst_dmem_n12326, MEM_stage_inst_dmem_n12327, MEM_stage_inst_dmem_n12328, MEM_stage_inst_dmem_n12329, MEM_stage_inst_dmem_n12330, MEM_stage_inst_dmem_n12331, MEM_stage_inst_dmem_n12332, MEM_stage_inst_dmem_n12333, MEM_stage_inst_dmem_n12334, MEM_stage_inst_dmem_n12335, MEM_stage_inst_dmem_n12336, MEM_stage_inst_dmem_n12337, MEM_stage_inst_dmem_n12338, MEM_stage_inst_dmem_n12339, MEM_stage_inst_dmem_n12340, MEM_stage_inst_dmem_n12341, MEM_stage_inst_dmem_n12342, MEM_stage_inst_dmem_n12343, MEM_stage_inst_dmem_n12344, MEM_stage_inst_dmem_n12345, MEM_stage_inst_dmem_n12346, MEM_stage_inst_dmem_n12347, MEM_stage_inst_dmem_n12348, MEM_stage_inst_dmem_n12349, MEM_stage_inst_dmem_n12350, MEM_stage_inst_dmem_n12351, MEM_stage_inst_dmem_n12352, MEM_stage_inst_dmem_n12353, MEM_stage_inst_dmem_n12354, MEM_stage_inst_dmem_n12355, MEM_stage_inst_dmem_n12356, MEM_stage_inst_dmem_n12357, MEM_stage_inst_dmem_n12358, MEM_stage_inst_dmem_n12359, MEM_stage_inst_dmem_n12360, MEM_stage_inst_dmem_n12361, MEM_stage_inst_dmem_n12362, MEM_stage_inst_dmem_n12363, MEM_stage_inst_dmem_n12364, MEM_stage_inst_dmem_n12365, MEM_stage_inst_dmem_n12366, MEM_stage_inst_dmem_n12367, MEM_stage_inst_dmem_n12368, MEM_stage_inst_dmem_n12369, MEM_stage_inst_dmem_n12370, MEM_stage_inst_dmem_n12371, MEM_stage_inst_dmem_n12372, MEM_stage_inst_dmem_n12373, MEM_stage_inst_dmem_n12374, MEM_stage_inst_dmem_n12375, MEM_stage_inst_dmem_n12376, MEM_stage_inst_dmem_n12377, MEM_stage_inst_dmem_n12378, MEM_stage_inst_dmem_n12379, MEM_stage_inst_dmem_n12380, MEM_stage_inst_dmem_n12381, MEM_stage_inst_dmem_n12382, MEM_stage_inst_dmem_n12383, MEM_stage_inst_dmem_n12384, MEM_stage_inst_dmem_n12385, MEM_stage_inst_dmem_n12386, MEM_stage_inst_dmem_n12387, MEM_stage_inst_dmem_n12388, MEM_stage_inst_dmem_n12389, MEM_stage_inst_dmem_n12390, MEM_stage_inst_dmem_n12391, MEM_stage_inst_dmem_n12392, MEM_stage_inst_dmem_n12393, MEM_stage_inst_dmem_n12394, MEM_stage_inst_dmem_n12395, MEM_stage_inst_dmem_n12396, MEM_stage_inst_dmem_n12397, MEM_stage_inst_dmem_n12398, MEM_stage_inst_dmem_n12399, MEM_stage_inst_dmem_n12400, MEM_stage_inst_dmem_n12401, MEM_stage_inst_dmem_n12402, MEM_stage_inst_dmem_n12403, MEM_stage_inst_dmem_n12404, MEM_stage_inst_dmem_n12405, MEM_stage_inst_dmem_n12406, MEM_stage_inst_dmem_n12407, MEM_stage_inst_dmem_n12408, MEM_stage_inst_dmem_n12409, MEM_stage_inst_dmem_n12410, MEM_stage_inst_dmem_n12411, MEM_stage_inst_dmem_n12412, MEM_stage_inst_dmem_n12413, MEM_stage_inst_dmem_n12414, MEM_stage_inst_dmem_n12415, MEM_stage_inst_dmem_n12416, MEM_stage_inst_dmem_n12417, MEM_stage_inst_dmem_n12418, MEM_stage_inst_dmem_n12419, MEM_stage_inst_dmem_n12420, MEM_stage_inst_dmem_n12421, MEM_stage_inst_dmem_n12422, MEM_stage_inst_dmem_n12423, MEM_stage_inst_dmem_n12424, MEM_stage_inst_dmem_n12425, MEM_stage_inst_dmem_n12426, MEM_stage_inst_dmem_n12427, MEM_stage_inst_dmem_n12428, MEM_stage_inst_dmem_n12429, MEM_stage_inst_dmem_n12430, MEM_stage_inst_dmem_n12431, MEM_stage_inst_dmem_n12432, MEM_stage_inst_dmem_n12433, MEM_stage_inst_dmem_n12434, MEM_stage_inst_dmem_n12435, MEM_stage_inst_dmem_n12436, MEM_stage_inst_dmem_n12437, MEM_stage_inst_dmem_n12438, MEM_stage_inst_dmem_n12439, MEM_stage_inst_dmem_n12440, MEM_stage_inst_dmem_n12441, MEM_stage_inst_dmem_n12442, MEM_stage_inst_dmem_n12443, MEM_stage_inst_dmem_n12444, MEM_stage_inst_dmem_n12445, MEM_stage_inst_dmem_n12446, MEM_stage_inst_dmem_n12447, MEM_stage_inst_dmem_n12448, MEM_stage_inst_dmem_n12449, MEM_stage_inst_dmem_n12450, MEM_stage_inst_dmem_n12451, MEM_stage_inst_dmem_n12452, MEM_stage_inst_dmem_n12453, MEM_stage_inst_dmem_n12454, MEM_stage_inst_dmem_n12455, MEM_stage_inst_dmem_n12456, MEM_stage_inst_dmem_n12457, MEM_stage_inst_dmem_n12458, MEM_stage_inst_dmem_n12459, MEM_stage_inst_dmem_n12460, MEM_stage_inst_dmem_n12461, MEM_stage_inst_dmem_n12462, MEM_stage_inst_dmem_n12463, MEM_stage_inst_dmem_n12464, MEM_stage_inst_dmem_n12465, MEM_stage_inst_dmem_n12466, MEM_stage_inst_dmem_n12467, MEM_stage_inst_dmem_n12468, MEM_stage_inst_dmem_n12469, MEM_stage_inst_dmem_n12470, MEM_stage_inst_dmem_n12471, MEM_stage_inst_dmem_n12472, MEM_stage_inst_dmem_n12473, MEM_stage_inst_dmem_n12474, MEM_stage_inst_dmem_n12475, MEM_stage_inst_dmem_n12476, MEM_stage_inst_dmem_n12477, MEM_stage_inst_dmem_n12478, MEM_stage_inst_dmem_n12479, MEM_stage_inst_dmem_n12480, MEM_stage_inst_dmem_n12481, MEM_stage_inst_dmem_n12482, MEM_stage_inst_dmem_n12483, MEM_stage_inst_dmem_n12484, MEM_stage_inst_dmem_n12485, MEM_stage_inst_dmem_n12486, MEM_stage_inst_dmem_n12487, MEM_stage_inst_dmem_n12488, MEM_stage_inst_dmem_n12489, MEM_stage_inst_dmem_n12490, MEM_stage_inst_dmem_n12491, MEM_stage_inst_dmem_n12492, MEM_stage_inst_dmem_n12493, MEM_stage_inst_dmem_n12494, MEM_stage_inst_dmem_n12495, MEM_stage_inst_dmem_n12496, MEM_stage_inst_dmem_n12497, MEM_stage_inst_dmem_n12498, MEM_stage_inst_dmem_n12499, MEM_stage_inst_dmem_n12500, MEM_stage_inst_dmem_n12501, MEM_stage_inst_dmem_n12502, MEM_stage_inst_dmem_n12503, MEM_stage_inst_dmem_n12504, MEM_stage_inst_dmem_n12505, MEM_stage_inst_dmem_n12506, MEM_stage_inst_dmem_n12507, MEM_stage_inst_dmem_n12508, MEM_stage_inst_dmem_n12509, MEM_stage_inst_dmem_n12510, MEM_stage_inst_dmem_n12511, MEM_stage_inst_dmem_n12512, MEM_stage_inst_dmem_n12513, MEM_stage_inst_dmem_n12514, MEM_stage_inst_dmem_n12515, MEM_stage_inst_dmem_n12516, MEM_stage_inst_dmem_n12517, MEM_stage_inst_dmem_n12518, MEM_stage_inst_dmem_n12519, MEM_stage_inst_dmem_n12520, MEM_stage_inst_dmem_n12521, MEM_stage_inst_dmem_n12522, MEM_stage_inst_dmem_n12523, MEM_stage_inst_dmem_n12524, MEM_stage_inst_dmem_n12525, MEM_stage_inst_dmem_n12526, MEM_stage_inst_dmem_n12527, MEM_stage_inst_dmem_n12528, MEM_stage_inst_dmem_n12529, MEM_stage_inst_dmem_n12530, MEM_stage_inst_dmem_n12531, MEM_stage_inst_dmem_n12532, MEM_stage_inst_dmem_n12533, MEM_stage_inst_dmem_n12534, MEM_stage_inst_dmem_n12535, MEM_stage_inst_dmem_n12536, MEM_stage_inst_dmem_n12537, MEM_stage_inst_dmem_n12538, MEM_stage_inst_dmem_n12539, MEM_stage_inst_dmem_n12540, MEM_stage_inst_dmem_n12541, MEM_stage_inst_dmem_n12542, MEM_stage_inst_dmem_n12543, MEM_stage_inst_dmem_n12544, MEM_stage_inst_dmem_n12545, MEM_stage_inst_dmem_n12546, MEM_stage_inst_dmem_n12547, MEM_stage_inst_dmem_n12548, MEM_stage_inst_dmem_n12549, MEM_stage_inst_dmem_n12550, MEM_stage_inst_dmem_n12551, MEM_stage_inst_dmem_n12552, MEM_stage_inst_dmem_n12553, MEM_stage_inst_dmem_n12554, MEM_stage_inst_dmem_n12555, MEM_stage_inst_dmem_n12556, MEM_stage_inst_dmem_n12557, MEM_stage_inst_dmem_n12558, MEM_stage_inst_dmem_n12559, MEM_stage_inst_dmem_n12560, MEM_stage_inst_dmem_n12561, MEM_stage_inst_dmem_n12562, MEM_stage_inst_dmem_n12563, MEM_stage_inst_dmem_n12564, MEM_stage_inst_dmem_n12565, MEM_stage_inst_dmem_n12566, MEM_stage_inst_dmem_n12567, MEM_stage_inst_dmem_n12568, MEM_stage_inst_dmem_n12569, MEM_stage_inst_dmem_n12570, MEM_stage_inst_dmem_n12571, MEM_stage_inst_dmem_n12572, MEM_stage_inst_dmem_n12573, MEM_stage_inst_dmem_n12574, MEM_stage_inst_dmem_n12575, MEM_stage_inst_dmem_n12576, MEM_stage_inst_dmem_n12577, MEM_stage_inst_dmem_n12578, MEM_stage_inst_dmem_n12579, MEM_stage_inst_dmem_n12580, MEM_stage_inst_dmem_n12581, MEM_stage_inst_dmem_n12582, MEM_stage_inst_dmem_n12583, MEM_stage_inst_dmem_n12584, MEM_stage_inst_dmem_n12585, MEM_stage_inst_dmem_n12586, MEM_stage_inst_dmem_n12587, MEM_stage_inst_dmem_n12588, MEM_stage_inst_dmem_n12589, MEM_stage_inst_dmem_n12590, MEM_stage_inst_dmem_n12591, MEM_stage_inst_dmem_n12592, MEM_stage_inst_dmem_n12593, MEM_stage_inst_dmem_n12594, MEM_stage_inst_dmem_n12595, MEM_stage_inst_dmem_n12596, MEM_stage_inst_dmem_n12597, MEM_stage_inst_dmem_n12598, MEM_stage_inst_dmem_n12599, MEM_stage_inst_dmem_n12600, MEM_stage_inst_dmem_n12601, MEM_stage_inst_dmem_n12602, MEM_stage_inst_dmem_n12603, MEM_stage_inst_dmem_n12604, MEM_stage_inst_dmem_n12605, MEM_stage_inst_dmem_n12606, MEM_stage_inst_dmem_n12607, MEM_stage_inst_dmem_n12608, MEM_stage_inst_dmem_n12609, MEM_stage_inst_dmem_n12610, MEM_stage_inst_dmem_n12611, MEM_stage_inst_dmem_n12612, MEM_stage_inst_dmem_n12613, MEM_stage_inst_dmem_n12614, MEM_stage_inst_dmem_n12615, MEM_stage_inst_dmem_n12616, MEM_stage_inst_dmem_n12617, MEM_stage_inst_dmem_n12618, MEM_stage_inst_dmem_n12619, MEM_stage_inst_dmem_n12620, MEM_stage_inst_dmem_n12621, MEM_stage_inst_dmem_n12622, MEM_stage_inst_dmem_n12623, MEM_stage_inst_dmem_n12624, MEM_stage_inst_dmem_n12625, MEM_stage_inst_dmem_n12626, MEM_stage_inst_dmem_n12627, MEM_stage_inst_dmem_n12628, MEM_stage_inst_dmem_n12629, MEM_stage_inst_dmem_n12630, MEM_stage_inst_dmem_n12631, MEM_stage_inst_dmem_n12632, MEM_stage_inst_dmem_n12633, MEM_stage_inst_dmem_n12634, MEM_stage_inst_dmem_n12635, MEM_stage_inst_dmem_n12636, MEM_stage_inst_dmem_n12637, MEM_stage_inst_dmem_n12638, MEM_stage_inst_dmem_n12639, MEM_stage_inst_dmem_n12640, MEM_stage_inst_dmem_n12641, MEM_stage_inst_dmem_n12642, MEM_stage_inst_dmem_n12643, MEM_stage_inst_dmem_n12644, MEM_stage_inst_dmem_n12645, MEM_stage_inst_dmem_n12646, MEM_stage_inst_dmem_n12647, MEM_stage_inst_dmem_n12648, MEM_stage_inst_dmem_n12649, MEM_stage_inst_dmem_n12650, MEM_stage_inst_dmem_n12651, MEM_stage_inst_dmem_n12652, MEM_stage_inst_dmem_n12653, MEM_stage_inst_dmem_n12654, MEM_stage_inst_dmem_n12655, MEM_stage_inst_dmem_n12656, MEM_stage_inst_dmem_n12657, MEM_stage_inst_dmem_n12658, MEM_stage_inst_dmem_n12659, MEM_stage_inst_dmem_n12660, MEM_stage_inst_dmem_n12661, MEM_stage_inst_dmem_n12662, MEM_stage_inst_dmem_n12663, MEM_stage_inst_dmem_n12664, MEM_stage_inst_dmem_n12665, MEM_stage_inst_dmem_n12666, MEM_stage_inst_dmem_n12667, MEM_stage_inst_dmem_n12668, MEM_stage_inst_dmem_n12669, MEM_stage_inst_dmem_n12670, MEM_stage_inst_dmem_n12671, MEM_stage_inst_dmem_n12672, MEM_stage_inst_dmem_n12673, MEM_stage_inst_dmem_n12674, MEM_stage_inst_dmem_n12675, MEM_stage_inst_dmem_n12676, MEM_stage_inst_dmem_n12677, MEM_stage_inst_dmem_n12678, MEM_stage_inst_dmem_n12679, MEM_stage_inst_dmem_n12680, MEM_stage_inst_dmem_n12681, MEM_stage_inst_dmem_n12682, MEM_stage_inst_dmem_n12683, MEM_stage_inst_dmem_n12684, MEM_stage_inst_dmem_n12685, MEM_stage_inst_dmem_n12686, MEM_stage_inst_dmem_n12687, MEM_stage_inst_dmem_n12688, MEM_stage_inst_dmem_n12689, MEM_stage_inst_dmem_n12690, MEM_stage_inst_dmem_n12691, MEM_stage_inst_dmem_n12692, MEM_stage_inst_dmem_n12693, MEM_stage_inst_dmem_n12694, MEM_stage_inst_dmem_n12695, MEM_stage_inst_dmem_n12696, MEM_stage_inst_dmem_n12697, MEM_stage_inst_dmem_n12698, MEM_stage_inst_dmem_n12699, MEM_stage_inst_dmem_n12700, MEM_stage_inst_dmem_n12701, MEM_stage_inst_dmem_n12702, MEM_stage_inst_dmem_n12703, MEM_stage_inst_dmem_n12704, MEM_stage_inst_dmem_n12705, MEM_stage_inst_dmem_n12706, MEM_stage_inst_dmem_n12707, MEM_stage_inst_dmem_n12708, MEM_stage_inst_dmem_n12709, MEM_stage_inst_dmem_n12710, MEM_stage_inst_dmem_n12711, MEM_stage_inst_dmem_n12712, MEM_stage_inst_dmem_n12713, MEM_stage_inst_dmem_n12714, MEM_stage_inst_dmem_n12715, MEM_stage_inst_dmem_n12716, MEM_stage_inst_dmem_n12717, MEM_stage_inst_dmem_n12718, MEM_stage_inst_dmem_n12719, MEM_stage_inst_dmem_n12720, MEM_stage_inst_dmem_n12721, MEM_stage_inst_dmem_n12722, MEM_stage_inst_dmem_n12723, MEM_stage_inst_dmem_n12724, MEM_stage_inst_dmem_n12725, MEM_stage_inst_dmem_n12726, MEM_stage_inst_dmem_n12727, MEM_stage_inst_dmem_n12728, MEM_stage_inst_dmem_n12729, MEM_stage_inst_dmem_n12730, MEM_stage_inst_dmem_n12731, MEM_stage_inst_dmem_n12732, MEM_stage_inst_dmem_n12733, MEM_stage_inst_dmem_n12734, MEM_stage_inst_dmem_n12735, MEM_stage_inst_dmem_n12736, MEM_stage_inst_dmem_n12737, MEM_stage_inst_dmem_n12738, MEM_stage_inst_dmem_n12739, MEM_stage_inst_dmem_n12740, MEM_stage_inst_dmem_n12741, MEM_stage_inst_dmem_n12742, MEM_stage_inst_dmem_n12743, MEM_stage_inst_dmem_n12744, MEM_stage_inst_dmem_n12745, MEM_stage_inst_dmem_n12746, MEM_stage_inst_dmem_n12747, MEM_stage_inst_dmem_n12748, MEM_stage_inst_dmem_n12749, MEM_stage_inst_dmem_n12750, MEM_stage_inst_dmem_n12751, MEM_stage_inst_dmem_n12752, MEM_stage_inst_dmem_n12753, MEM_stage_inst_dmem_n12754, MEM_stage_inst_dmem_n12755, MEM_stage_inst_dmem_n12756, MEM_stage_inst_dmem_n12757, MEM_stage_inst_dmem_n12758, MEM_stage_inst_dmem_n12759, MEM_stage_inst_dmem_n12760, MEM_stage_inst_dmem_n12761, MEM_stage_inst_dmem_n12762, MEM_stage_inst_dmem_n12763, MEM_stage_inst_dmem_n12764, MEM_stage_inst_dmem_n12765, MEM_stage_inst_dmem_n12766, MEM_stage_inst_dmem_n12767, MEM_stage_inst_dmem_n12768, MEM_stage_inst_dmem_n12769, MEM_stage_inst_dmem_n12770, MEM_stage_inst_dmem_n12771, MEM_stage_inst_dmem_n12772, MEM_stage_inst_dmem_n12773, MEM_stage_inst_dmem_n12774, MEM_stage_inst_dmem_n12775, MEM_stage_inst_dmem_n12776, MEM_stage_inst_dmem_n12777, MEM_stage_inst_dmem_n12778, MEM_stage_inst_dmem_n12779, MEM_stage_inst_dmem_n12780, MEM_stage_inst_dmem_n12781, MEM_stage_inst_dmem_n12782, MEM_stage_inst_dmem_n12783, MEM_stage_inst_dmem_n12784, MEM_stage_inst_dmem_n12785, MEM_stage_inst_dmem_n12786, MEM_stage_inst_dmem_n12787, MEM_stage_inst_dmem_n12788, MEM_stage_inst_dmem_n12789, MEM_stage_inst_dmem_n12790, MEM_stage_inst_dmem_n12791, MEM_stage_inst_dmem_n12792, MEM_stage_inst_dmem_n12793, MEM_stage_inst_dmem_n12794, MEM_stage_inst_dmem_n12795, MEM_stage_inst_dmem_n12796, MEM_stage_inst_dmem_n12797, MEM_stage_inst_dmem_n12798, MEM_stage_inst_dmem_n12799, MEM_stage_inst_dmem_n12800, MEM_stage_inst_dmem_n12801, MEM_stage_inst_dmem_n12802, MEM_stage_inst_dmem_n12803, MEM_stage_inst_dmem_n12804, MEM_stage_inst_dmem_n12805, MEM_stage_inst_dmem_n12806, MEM_stage_inst_dmem_n12807, MEM_stage_inst_dmem_n12808, MEM_stage_inst_dmem_n12809, MEM_stage_inst_dmem_n12810, MEM_stage_inst_dmem_n12811, MEM_stage_inst_dmem_n12812, MEM_stage_inst_dmem_n12813, MEM_stage_inst_dmem_n12814, MEM_stage_inst_dmem_n12815, MEM_stage_inst_dmem_n12816, MEM_stage_inst_dmem_n12817, MEM_stage_inst_dmem_n12818, MEM_stage_inst_dmem_n12819, MEM_stage_inst_dmem_n12820, MEM_stage_inst_dmem_n12821, MEM_stage_inst_dmem_n12822, MEM_stage_inst_dmem_n12823, MEM_stage_inst_dmem_n12824, MEM_stage_inst_dmem_n12825, MEM_stage_inst_dmem_n12826, MEM_stage_inst_dmem_n12827, MEM_stage_inst_dmem_n12828, MEM_stage_inst_dmem_n12829, MEM_stage_inst_dmem_n12830, MEM_stage_inst_dmem_n12831, MEM_stage_inst_dmem_n12832, MEM_stage_inst_dmem_n12833, MEM_stage_inst_dmem_n12834, MEM_stage_inst_dmem_n12835, MEM_stage_inst_dmem_n12836, MEM_stage_inst_dmem_n12837, MEM_stage_inst_dmem_n12838, MEM_stage_inst_dmem_n12839, MEM_stage_inst_dmem_n12840, MEM_stage_inst_dmem_n12841, MEM_stage_inst_dmem_n12842, MEM_stage_inst_dmem_n12843, MEM_stage_inst_dmem_n12844, MEM_stage_inst_dmem_n12845, MEM_stage_inst_dmem_n12846, MEM_stage_inst_dmem_n12847, MEM_stage_inst_dmem_n12848, MEM_stage_inst_dmem_n12849, MEM_stage_inst_dmem_n12850, MEM_stage_inst_dmem_n12851, MEM_stage_inst_dmem_n12852, MEM_stage_inst_dmem_n12853, MEM_stage_inst_dmem_n12854, MEM_stage_inst_dmem_n12855, MEM_stage_inst_dmem_n12856, MEM_stage_inst_dmem_n12857, MEM_stage_inst_dmem_n12858;
wire MEM_stage_inst_mem_read_data_15, MEM_stage_inst_mem_read_data_14, MEM_stage_inst_mem_read_data_13, MEM_stage_inst_mem_read_data_12, MEM_stage_inst_mem_read_data_11, MEM_stage_inst_mem_read_data_10, MEM_stage_inst_mem_read_data_9, MEM_stage_inst_mem_read_data_8, MEM_stage_inst_mem_read_data_7, MEM_stage_inst_mem_read_data_6, MEM_stage_inst_mem_read_data_5, MEM_stage_inst_mem_read_data_4, MEM_stage_inst_mem_read_data_3, MEM_stage_inst_mem_read_data_2, MEM_stage_inst_mem_read_data_1, MEM_stage_inst_mem_read_data_0, n1740, n1742, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, MEM_stage_inst_dmem_n21508, MEM_stage_inst_dmem_n21507, MEM_stage_inst_dmem_n21506, MEM_stage_inst_dmem_n21505, MEM_stage_inst_dmem_n21503, MEM_stage_inst_dmem_n21502, MEM_stage_inst_dmem_n21501, MEM_stage_inst_dmem_n21500, MEM_stage_inst_dmem_n21499, MEM_stage_inst_dmem_n21498, MEM_stage_inst_dmem_n21497, MEM_stage_inst_dmem_n21496, MEM_stage_inst_dmem_n21495, MEM_stage_inst_dmem_n21494, MEM_stage_inst_dmem_n21493, MEM_stage_inst_dmem_n21492, MEM_stage_inst_dmem_n21491, MEM_stage_inst_dmem_n21490, MEM_stage_inst_dmem_n21489, MEM_stage_inst_dmem_n21488, MEM_stage_inst_dmem_n21487, MEM_stage_inst_dmem_n21486, MEM_stage_inst_dmem_n21485, MEM_stage_inst_dmem_n21484, MEM_stage_inst_dmem_n21483, MEM_stage_inst_dmem_n21482, MEM_stage_inst_dmem_n21481, MEM_stage_inst_dmem_n21480, MEM_stage_inst_dmem_n21479, MEM_stage_inst_dmem_n21478, MEM_stage_inst_dmem_n21477, MEM_stage_inst_dmem_n21476, MEM_stage_inst_dmem_n21475, MEM_stage_inst_dmem_n21474, MEM_stage_inst_dmem_n21473, MEM_stage_inst_dmem_n21472, MEM_stage_inst_dmem_n21471, MEM_stage_inst_dmem_n21470, MEM_stage_inst_dmem_n21469, MEM_stage_inst_dmem_n21468, MEM_stage_inst_dmem_n21467, MEM_stage_inst_dmem_n21466, MEM_stage_inst_dmem_n21465, MEM_stage_inst_dmem_n21464, MEM_stage_inst_dmem_n21463, MEM_stage_inst_dmem_n21462, MEM_stage_inst_dmem_n21461, MEM_stage_inst_dmem_n21460, MEM_stage_inst_dmem_n21459, MEM_stage_inst_dmem_n21458, MEM_stage_inst_dmem_n21457, MEM_stage_inst_dmem_n21456, MEM_stage_inst_dmem_n21455, MEM_stage_inst_dmem_n21454, MEM_stage_inst_dmem_n21453, MEM_stage_inst_dmem_n21452, MEM_stage_inst_dmem_n21451, MEM_stage_inst_dmem_n21450, MEM_stage_inst_dmem_n21449, MEM_stage_inst_dmem_n21448, MEM_stage_inst_dmem_n21447, MEM_stage_inst_dmem_n21446, MEM_stage_inst_dmem_n21445, MEM_stage_inst_dmem_n21444, MEM_stage_inst_dmem_n21443, MEM_stage_inst_dmem_n21442, MEM_stage_inst_dmem_n21441, MEM_stage_inst_dmem_n21440, MEM_stage_inst_dmem_n21439, MEM_stage_inst_dmem_n21438, MEM_stage_inst_dmem_n21437, MEM_stage_inst_dmem_n21436, MEM_stage_inst_dmem_n21435, MEM_stage_inst_dmem_n21434, MEM_stage_inst_dmem_n21433, MEM_stage_inst_dmem_n21432, MEM_stage_inst_dmem_n21431, MEM_stage_inst_dmem_n21430, MEM_stage_inst_dmem_n21429, MEM_stage_inst_dmem_n21428, MEM_stage_inst_dmem_n21427, MEM_stage_inst_dmem_n21426, MEM_stage_inst_dmem_n21425, MEM_stage_inst_dmem_n21424, MEM_stage_inst_dmem_n21423, MEM_stage_inst_dmem_n21422, MEM_stage_inst_dmem_n21421, MEM_stage_inst_dmem_n21420, MEM_stage_inst_dmem_n21419, MEM_stage_inst_dmem_n21418, MEM_stage_inst_dmem_n21417, MEM_stage_inst_dmem_n21416, MEM_stage_inst_dmem_n21415, MEM_stage_inst_dmem_n21414, MEM_stage_inst_dmem_n21413, MEM_stage_inst_dmem_n21412, MEM_stage_inst_dmem_n21411, MEM_stage_inst_dmem_n21410, MEM_stage_inst_dmem_n21409, MEM_stage_inst_dmem_n21408, MEM_stage_inst_dmem_n21407, MEM_stage_inst_dmem_n21406, MEM_stage_inst_dmem_n21405, MEM_stage_inst_dmem_n21404, MEM_stage_inst_dmem_n21403, MEM_stage_inst_dmem_n21402, MEM_stage_inst_dmem_n21401, MEM_stage_inst_dmem_n21400, MEM_stage_inst_dmem_n21399, MEM_stage_inst_dmem_n21398, MEM_stage_inst_dmem_n21397, MEM_stage_inst_dmem_n21396, MEM_stage_inst_dmem_n21395, MEM_stage_inst_dmem_n21394, MEM_stage_inst_dmem_n21393, MEM_stage_inst_dmem_n21392, MEM_stage_inst_dmem_n21391, MEM_stage_inst_dmem_n21390, MEM_stage_inst_dmem_n21389, MEM_stage_inst_dmem_n21388, MEM_stage_inst_dmem_n21387, MEM_stage_inst_dmem_n21386, MEM_stage_inst_dmem_n21385, MEM_stage_inst_dmem_n21384, MEM_stage_inst_dmem_n21383, MEM_stage_inst_dmem_n21382, MEM_stage_inst_dmem_n21381, MEM_stage_inst_dmem_n21380, MEM_stage_inst_dmem_n21379, MEM_stage_inst_dmem_n21378, MEM_stage_inst_dmem_n21377, MEM_stage_inst_dmem_n21376, MEM_stage_inst_dmem_n21375, MEM_stage_inst_dmem_n21374, MEM_stage_inst_dmem_n21373, MEM_stage_inst_dmem_n21372, MEM_stage_inst_dmem_n21371, MEM_stage_inst_dmem_n21370, MEM_stage_inst_dmem_n21369, MEM_stage_inst_dmem_n21368, MEM_stage_inst_dmem_n21367, MEM_stage_inst_dmem_n21366, MEM_stage_inst_dmem_n21365, MEM_stage_inst_dmem_n21364, MEM_stage_inst_dmem_n21363, MEM_stage_inst_dmem_n21362, MEM_stage_inst_dmem_n21361, MEM_stage_inst_dmem_n21360, MEM_stage_inst_dmem_n21359, MEM_stage_inst_dmem_n21358, MEM_stage_inst_dmem_n21357, MEM_stage_inst_dmem_n21356, MEM_stage_inst_dmem_n21355, MEM_stage_inst_dmem_n21354, MEM_stage_inst_dmem_n21353, MEM_stage_inst_dmem_n21351, MEM_stage_inst_dmem_n21350, MEM_stage_inst_dmem_n21349, MEM_stage_inst_dmem_n21348, MEM_stage_inst_dmem_n21347, MEM_stage_inst_dmem_n21346, MEM_stage_inst_dmem_n21344, MEM_stage_inst_dmem_n21343, MEM_stage_inst_dmem_n21342, MEM_stage_inst_dmem_n21341, MEM_stage_inst_dmem_n21340, MEM_stage_inst_dmem_n21339, MEM_stage_inst_dmem_n21338, MEM_stage_inst_dmem_n21337, MEM_stage_inst_dmem_n21336, MEM_stage_inst_dmem_n21335, MEM_stage_inst_dmem_n21334, MEM_stage_inst_dmem_n21333, MEM_stage_inst_dmem_n21332, MEM_stage_inst_dmem_n21331, MEM_stage_inst_dmem_n21330, MEM_stage_inst_dmem_n21329, MEM_stage_inst_dmem_n21328, MEM_stage_inst_dmem_n21327, MEM_stage_inst_dmem_n21326, MEM_stage_inst_dmem_n21325, MEM_stage_inst_dmem_n21324, MEM_stage_inst_dmem_n21323, MEM_stage_inst_dmem_n21322, MEM_stage_inst_dmem_n21321, MEM_stage_inst_dmem_n21320, MEM_stage_inst_dmem_n21319, MEM_stage_inst_dmem_n21318, MEM_stage_inst_dmem_n21317, MEM_stage_inst_dmem_n21316, MEM_stage_inst_dmem_n21315, MEM_stage_inst_dmem_n21314, MEM_stage_inst_dmem_n21313, MEM_stage_inst_dmem_n21312, MEM_stage_inst_dmem_n21311, MEM_stage_inst_dmem_n21310, MEM_stage_inst_dmem_n21309, MEM_stage_inst_dmem_n21308, MEM_stage_inst_dmem_n21307, MEM_stage_inst_dmem_n21306, MEM_stage_inst_dmem_n21305, MEM_stage_inst_dmem_n21304, MEM_stage_inst_dmem_n21303, MEM_stage_inst_dmem_n21302, MEM_stage_inst_dmem_n21301, MEM_stage_inst_dmem_n21300, MEM_stage_inst_dmem_n21299, MEM_stage_inst_dmem_n21298, MEM_stage_inst_dmem_n21297, MEM_stage_inst_dmem_n21296, MEM_stage_inst_dmem_n21295, MEM_stage_inst_dmem_n21294, MEM_stage_inst_dmem_n21293, MEM_stage_inst_dmem_n21292, MEM_stage_inst_dmem_n21291, MEM_stage_inst_dmem_n21290, MEM_stage_inst_dmem_n21289, MEM_stage_inst_dmem_n21288, MEM_stage_inst_dmem_n21287, MEM_stage_inst_dmem_n21286, MEM_stage_inst_dmem_n21285, MEM_stage_inst_dmem_n21284, MEM_stage_inst_dmem_n21283, MEM_stage_inst_dmem_n21282, MEM_stage_inst_dmem_n21281, MEM_stage_inst_dmem_n21280, MEM_stage_inst_dmem_n21279, MEM_stage_inst_dmem_n21278, MEM_stage_inst_dmem_n21277, MEM_stage_inst_dmem_n21276, MEM_stage_inst_dmem_n21275, MEM_stage_inst_dmem_n21274, MEM_stage_inst_dmem_n21273, MEM_stage_inst_dmem_n21272, MEM_stage_inst_dmem_n21271, MEM_stage_inst_dmem_n21270, MEM_stage_inst_dmem_n21269, MEM_stage_inst_dmem_n21268, MEM_stage_inst_dmem_n21267, MEM_stage_inst_dmem_n21266, MEM_stage_inst_dmem_n21265, MEM_stage_inst_dmem_n21264, MEM_stage_inst_dmem_n21263, MEM_stage_inst_dmem_n21262, MEM_stage_inst_dmem_n21261, MEM_stage_inst_dmem_n21260, MEM_stage_inst_dmem_n21259, MEM_stage_inst_dmem_n21258, MEM_stage_inst_dmem_n21257, MEM_stage_inst_dmem_n21256, MEM_stage_inst_dmem_n21255, MEM_stage_inst_dmem_n21254, MEM_stage_inst_dmem_n21253, MEM_stage_inst_dmem_n21252, MEM_stage_inst_dmem_n21251, MEM_stage_inst_dmem_n21250, MEM_stage_inst_dmem_n21249, MEM_stage_inst_dmem_n21248, MEM_stage_inst_dmem_n21247, MEM_stage_inst_dmem_n21246, MEM_stage_inst_dmem_n21245, MEM_stage_inst_dmem_n21244, MEM_stage_inst_dmem_n21243, MEM_stage_inst_dmem_n21242, MEM_stage_inst_dmem_n21241, MEM_stage_inst_dmem_n21240, MEM_stage_inst_dmem_n21239, MEM_stage_inst_dmem_n21238, MEM_stage_inst_dmem_n21237, MEM_stage_inst_dmem_n21236, MEM_stage_inst_dmem_n21235, MEM_stage_inst_dmem_n21234, MEM_stage_inst_dmem_n21233, MEM_stage_inst_dmem_n21232, MEM_stage_inst_dmem_n21231, MEM_stage_inst_dmem_n21230, MEM_stage_inst_dmem_n21229, MEM_stage_inst_dmem_n21228, MEM_stage_inst_dmem_n21227, MEM_stage_inst_dmem_n21226, MEM_stage_inst_dmem_n21225, MEM_stage_inst_dmem_n21224, MEM_stage_inst_dmem_n21223, MEM_stage_inst_dmem_n21222, MEM_stage_inst_dmem_n21221, MEM_stage_inst_dmem_n21220, MEM_stage_inst_dmem_n21219, MEM_stage_inst_dmem_n21218, MEM_stage_inst_dmem_n21217, MEM_stage_inst_dmem_n21216, MEM_stage_inst_dmem_n21215, MEM_stage_inst_dmem_n21214, MEM_stage_inst_dmem_n21213, MEM_stage_inst_dmem_n21212, MEM_stage_inst_dmem_n21211, MEM_stage_inst_dmem_n21210, MEM_stage_inst_dmem_n21209, MEM_stage_inst_dmem_n21208, MEM_stage_inst_dmem_n21207, MEM_stage_inst_dmem_n21206, MEM_stage_inst_dmem_n21205, MEM_stage_inst_dmem_n21204, MEM_stage_inst_dmem_n21203, MEM_stage_inst_dmem_n21202, MEM_stage_inst_dmem_n21201, MEM_stage_inst_dmem_n21200, MEM_stage_inst_dmem_n21199, MEM_stage_inst_dmem_n21198, MEM_stage_inst_dmem_n21197, MEM_stage_inst_dmem_n21196, MEM_stage_inst_dmem_n21195, MEM_stage_inst_dmem_n21194, MEM_stage_inst_dmem_n21193, MEM_stage_inst_dmem_n21192, MEM_stage_inst_dmem_n21191, MEM_stage_inst_dmem_n21190, MEM_stage_inst_dmem_n21189, MEM_stage_inst_dmem_n21188, MEM_stage_inst_dmem_n21187, MEM_stage_inst_dmem_n21186, MEM_stage_inst_dmem_n21185, MEM_stage_inst_dmem_n21184, MEM_stage_inst_dmem_n21183, MEM_stage_inst_dmem_n21182, MEM_stage_inst_dmem_n21181, MEM_stage_inst_dmem_n21180, MEM_stage_inst_dmem_n21179, MEM_stage_inst_dmem_n21178, MEM_stage_inst_dmem_n21177, MEM_stage_inst_dmem_n21176, MEM_stage_inst_dmem_n21175, MEM_stage_inst_dmem_n21174, MEM_stage_inst_dmem_n21173, MEM_stage_inst_dmem_n21172, MEM_stage_inst_dmem_n21171, MEM_stage_inst_dmem_n21170, MEM_stage_inst_dmem_n21169, MEM_stage_inst_dmem_n21168, MEM_stage_inst_dmem_n21167, MEM_stage_inst_dmem_n21166, MEM_stage_inst_dmem_n21165, MEM_stage_inst_dmem_n21164, MEM_stage_inst_dmem_n21163, MEM_stage_inst_dmem_n21162, MEM_stage_inst_dmem_n21161, MEM_stage_inst_dmem_n21160, MEM_stage_inst_dmem_n21159, MEM_stage_inst_dmem_n21158, MEM_stage_inst_dmem_n21157, MEM_stage_inst_dmem_n21156, MEM_stage_inst_dmem_n21155, MEM_stage_inst_dmem_n21154, MEM_stage_inst_dmem_n21153, MEM_stage_inst_dmem_n21152, MEM_stage_inst_dmem_n21151, MEM_stage_inst_dmem_n21150, MEM_stage_inst_dmem_n21149, MEM_stage_inst_dmem_n21148, MEM_stage_inst_dmem_n21147, MEM_stage_inst_dmem_n21146, MEM_stage_inst_dmem_n21145, MEM_stage_inst_dmem_n21144, MEM_stage_inst_dmem_n21143, MEM_stage_inst_dmem_n21142, MEM_stage_inst_dmem_n21141, MEM_stage_inst_dmem_n21140, MEM_stage_inst_dmem_n21139, MEM_stage_inst_dmem_n21138, MEM_stage_inst_dmem_n21137, MEM_stage_inst_dmem_n21136, MEM_stage_inst_dmem_n21135, MEM_stage_inst_dmem_n21134, MEM_stage_inst_dmem_n21133, MEM_stage_inst_dmem_n21132, MEM_stage_inst_dmem_n21131, MEM_stage_inst_dmem_n21130, MEM_stage_inst_dmem_n21129, MEM_stage_inst_dmem_n21128, MEM_stage_inst_dmem_n21127, MEM_stage_inst_dmem_n21126, MEM_stage_inst_dmem_n21125, MEM_stage_inst_dmem_n21124, MEM_stage_inst_dmem_n21123, MEM_stage_inst_dmem_n21122, MEM_stage_inst_dmem_n21121, MEM_stage_inst_dmem_n21120, MEM_stage_inst_dmem_n21119, MEM_stage_inst_dmem_n21118, MEM_stage_inst_dmem_n21117, MEM_stage_inst_dmem_n21116, MEM_stage_inst_dmem_n21115, MEM_stage_inst_dmem_n21114, MEM_stage_inst_dmem_n21113, MEM_stage_inst_dmem_n21112, MEM_stage_inst_dmem_n21111, MEM_stage_inst_dmem_n21110, MEM_stage_inst_dmem_n21109, MEM_stage_inst_dmem_n21108, MEM_stage_inst_dmem_n21107, MEM_stage_inst_dmem_n21106, MEM_stage_inst_dmem_n21105, MEM_stage_inst_dmem_n21104, MEM_stage_inst_dmem_n21103, MEM_stage_inst_dmem_n21102, MEM_stage_inst_dmem_n21101, MEM_stage_inst_dmem_n21100, MEM_stage_inst_dmem_n21099, MEM_stage_inst_dmem_n21098, MEM_stage_inst_dmem_n21097, MEM_stage_inst_dmem_n21096, MEM_stage_inst_dmem_n21095, MEM_stage_inst_dmem_n21094, MEM_stage_inst_dmem_n21093, MEM_stage_inst_dmem_n21092, MEM_stage_inst_dmem_n21091, MEM_stage_inst_dmem_n21090, MEM_stage_inst_dmem_n21089, MEM_stage_inst_dmem_n21088, MEM_stage_inst_dmem_n21087, MEM_stage_inst_dmem_n21086, MEM_stage_inst_dmem_n21085, MEM_stage_inst_dmem_n21084, MEM_stage_inst_dmem_n21083, MEM_stage_inst_dmem_n21082, MEM_stage_inst_dmem_n21081, MEM_stage_inst_dmem_n21080, MEM_stage_inst_dmem_n21079, MEM_stage_inst_dmem_n21078, MEM_stage_inst_dmem_n21077, MEM_stage_inst_dmem_n21076, MEM_stage_inst_dmem_n21075, MEM_stage_inst_dmem_n21074, MEM_stage_inst_dmem_n21073, MEM_stage_inst_dmem_n21072, MEM_stage_inst_dmem_n21071, MEM_stage_inst_dmem_n21070, MEM_stage_inst_dmem_n21069, MEM_stage_inst_dmem_n21068, MEM_stage_inst_dmem_n21067, MEM_stage_inst_dmem_n21066, MEM_stage_inst_dmem_n21065, MEM_stage_inst_dmem_n21064, MEM_stage_inst_dmem_n21063, MEM_stage_inst_dmem_n21062, MEM_stage_inst_dmem_n21061, MEM_stage_inst_dmem_n21060, MEM_stage_inst_dmem_n21059, MEM_stage_inst_dmem_n21058, MEM_stage_inst_dmem_n21057, MEM_stage_inst_dmem_n21056, MEM_stage_inst_dmem_n21055, MEM_stage_inst_dmem_n21054, MEM_stage_inst_dmem_n21053, MEM_stage_inst_dmem_n21052, MEM_stage_inst_dmem_n21051, MEM_stage_inst_dmem_n21050, MEM_stage_inst_dmem_n21049, MEM_stage_inst_dmem_n21048, MEM_stage_inst_dmem_n21047, MEM_stage_inst_dmem_n21046, MEM_stage_inst_dmem_n21045, MEM_stage_inst_dmem_n21044, MEM_stage_inst_dmem_n21043, MEM_stage_inst_dmem_n21042, MEM_stage_inst_dmem_n21041, MEM_stage_inst_dmem_n21040, MEM_stage_inst_dmem_n21039, MEM_stage_inst_dmem_n21038, MEM_stage_inst_dmem_n21037, MEM_stage_inst_dmem_n21036, MEM_stage_inst_dmem_n21035, MEM_stage_inst_dmem_n21034, MEM_stage_inst_dmem_n21033, MEM_stage_inst_dmem_n21032, MEM_stage_inst_dmem_n21031, MEM_stage_inst_dmem_n21030, MEM_stage_inst_dmem_n21029, MEM_stage_inst_dmem_n21028, MEM_stage_inst_dmem_n21027, MEM_stage_inst_dmem_n21026, MEM_stage_inst_dmem_n21025, MEM_stage_inst_dmem_n21024, MEM_stage_inst_dmem_n21023, MEM_stage_inst_dmem_n21022, MEM_stage_inst_dmem_n21021, MEM_stage_inst_dmem_n21020, MEM_stage_inst_dmem_n21019, MEM_stage_inst_dmem_n21018, MEM_stage_inst_dmem_n21017, MEM_stage_inst_dmem_n21016, MEM_stage_inst_dmem_n21015, MEM_stage_inst_dmem_n21014, MEM_stage_inst_dmem_n21013, MEM_stage_inst_dmem_n21012, MEM_stage_inst_dmem_n21011, MEM_stage_inst_dmem_n21010, MEM_stage_inst_dmem_n21009, MEM_stage_inst_dmem_n21008, MEM_stage_inst_dmem_n21007, MEM_stage_inst_dmem_n21006, MEM_stage_inst_dmem_n21005, MEM_stage_inst_dmem_n21004, MEM_stage_inst_dmem_n21003, MEM_stage_inst_dmem_n21002, MEM_stage_inst_dmem_n21001, MEM_stage_inst_dmem_n21000, MEM_stage_inst_dmem_n20999, MEM_stage_inst_dmem_n20998, MEM_stage_inst_dmem_n20997, MEM_stage_inst_dmem_n20996, MEM_stage_inst_dmem_n20995, MEM_stage_inst_dmem_n20994, MEM_stage_inst_dmem_n20993, MEM_stage_inst_dmem_n20992, MEM_stage_inst_dmem_n20991, MEM_stage_inst_dmem_n20990, MEM_stage_inst_dmem_n20989, MEM_stage_inst_dmem_n20988, MEM_stage_inst_dmem_n20987, MEM_stage_inst_dmem_n20986, MEM_stage_inst_dmem_n20985, MEM_stage_inst_dmem_n20984, MEM_stage_inst_dmem_n20983, MEM_stage_inst_dmem_n20982, MEM_stage_inst_dmem_n20981, MEM_stage_inst_dmem_n20980, MEM_stage_inst_dmem_n20979, MEM_stage_inst_dmem_n20978, MEM_stage_inst_dmem_n20977, MEM_stage_inst_dmem_n20976, MEM_stage_inst_dmem_n20975, MEM_stage_inst_dmem_n20974, MEM_stage_inst_dmem_n20973, MEM_stage_inst_dmem_n20972, MEM_stage_inst_dmem_n20971, MEM_stage_inst_dmem_n20970, MEM_stage_inst_dmem_n20969, MEM_stage_inst_dmem_n20968, MEM_stage_inst_dmem_n20967, MEM_stage_inst_dmem_n20966, MEM_stage_inst_dmem_n20965, MEM_stage_inst_dmem_n20964, MEM_stage_inst_dmem_n20963, MEM_stage_inst_dmem_n20962, MEM_stage_inst_dmem_n20961, MEM_stage_inst_dmem_n20960, MEM_stage_inst_dmem_n20959, MEM_stage_inst_dmem_n20958, MEM_stage_inst_dmem_n20957, MEM_stage_inst_dmem_n20956, MEM_stage_inst_dmem_n20955, MEM_stage_inst_dmem_n20954, MEM_stage_inst_dmem_n20953, MEM_stage_inst_dmem_n20952, MEM_stage_inst_dmem_n20951, MEM_stage_inst_dmem_n20950, MEM_stage_inst_dmem_n20949, MEM_stage_inst_dmem_n20948, MEM_stage_inst_dmem_n20947, MEM_stage_inst_dmem_n20946, MEM_stage_inst_dmem_n20945, MEM_stage_inst_dmem_n20944, MEM_stage_inst_dmem_n20943, MEM_stage_inst_dmem_n20942, MEM_stage_inst_dmem_n20941, MEM_stage_inst_dmem_n20940, MEM_stage_inst_dmem_n20939, MEM_stage_inst_dmem_n20938, MEM_stage_inst_dmem_n20937, MEM_stage_inst_dmem_n20936, MEM_stage_inst_dmem_n20935, MEM_stage_inst_dmem_n20934, MEM_stage_inst_dmem_n20933, MEM_stage_inst_dmem_n20932, MEM_stage_inst_dmem_n20931, MEM_stage_inst_dmem_n20930, MEM_stage_inst_dmem_n20929, MEM_stage_inst_dmem_n20928, MEM_stage_inst_dmem_n20927, MEM_stage_inst_dmem_n20926, MEM_stage_inst_dmem_n20925, MEM_stage_inst_dmem_n20924, MEM_stage_inst_dmem_n20923, MEM_stage_inst_dmem_n20922, MEM_stage_inst_dmem_n20921, MEM_stage_inst_dmem_n20920, MEM_stage_inst_dmem_n20918, MEM_stage_inst_dmem_n20917, MEM_stage_inst_dmem_n20916, MEM_stage_inst_dmem_n20915, MEM_stage_inst_dmem_n20914, MEM_stage_inst_dmem_n20913, MEM_stage_inst_dmem_n20912, MEM_stage_inst_dmem_n20911, MEM_stage_inst_dmem_n20910, MEM_stage_inst_dmem_n20909, MEM_stage_inst_dmem_n20908, MEM_stage_inst_dmem_n20907, MEM_stage_inst_dmem_n20906, MEM_stage_inst_dmem_n20905, MEM_stage_inst_dmem_n20904, MEM_stage_inst_dmem_n20903, MEM_stage_inst_dmem_n20902, MEM_stage_inst_dmem_n20901, MEM_stage_inst_dmem_n20900, MEM_stage_inst_dmem_n20899, MEM_stage_inst_dmem_n20898, MEM_stage_inst_dmem_n20897, MEM_stage_inst_dmem_n20896, MEM_stage_inst_dmem_n20895, MEM_stage_inst_dmem_n20894, MEM_stage_inst_dmem_n20893, MEM_stage_inst_dmem_n20892, MEM_stage_inst_dmem_n20891, MEM_stage_inst_dmem_n20890, MEM_stage_inst_dmem_n20889, MEM_stage_inst_dmem_n20888, MEM_stage_inst_dmem_n20887, MEM_stage_inst_dmem_n20886, MEM_stage_inst_dmem_n20885, MEM_stage_inst_dmem_n20884, MEM_stage_inst_dmem_n20883, MEM_stage_inst_dmem_n20882, MEM_stage_inst_dmem_n20881, MEM_stage_inst_dmem_n20880, MEM_stage_inst_dmem_n20879, MEM_stage_inst_dmem_n20878, MEM_stage_inst_dmem_n20877, MEM_stage_inst_dmem_n20876, MEM_stage_inst_dmem_n20875, MEM_stage_inst_dmem_n20874, MEM_stage_inst_dmem_n20873, MEM_stage_inst_dmem_n20872, MEM_stage_inst_dmem_n20871, MEM_stage_inst_dmem_n20870, MEM_stage_inst_dmem_n20869, MEM_stage_inst_dmem_n20868, MEM_stage_inst_dmem_n20867, MEM_stage_inst_dmem_n20866, MEM_stage_inst_dmem_n20865, MEM_stage_inst_dmem_n20864, MEM_stage_inst_dmem_n20863, MEM_stage_inst_dmem_n20862, MEM_stage_inst_dmem_n20861, MEM_stage_inst_dmem_n20860, MEM_stage_inst_dmem_n20859, MEM_stage_inst_dmem_n20858, MEM_stage_inst_dmem_n20857, MEM_stage_inst_dmem_n20856, MEM_stage_inst_dmem_n20855, MEM_stage_inst_dmem_n20854, MEM_stage_inst_dmem_n20853, MEM_stage_inst_dmem_n20852, MEM_stage_inst_dmem_n20851, MEM_stage_inst_dmem_n20850, MEM_stage_inst_dmem_n20849, MEM_stage_inst_dmem_n20848, MEM_stage_inst_dmem_n20847, MEM_stage_inst_dmem_n20846, MEM_stage_inst_dmem_n20845, MEM_stage_inst_dmem_n20844, MEM_stage_inst_dmem_n20843, MEM_stage_inst_dmem_n20842, MEM_stage_inst_dmem_n20841, MEM_stage_inst_dmem_n20840, MEM_stage_inst_dmem_n20839, MEM_stage_inst_dmem_n20838, MEM_stage_inst_dmem_n20837, MEM_stage_inst_dmem_n20836, MEM_stage_inst_dmem_n20835, MEM_stage_inst_dmem_n20834, MEM_stage_inst_dmem_n20833, MEM_stage_inst_dmem_n20832, MEM_stage_inst_dmem_n20831, MEM_stage_inst_dmem_n20830, MEM_stage_inst_dmem_n20829, MEM_stage_inst_dmem_n20828, MEM_stage_inst_dmem_n20827, MEM_stage_inst_dmem_n20826, MEM_stage_inst_dmem_n20825, MEM_stage_inst_dmem_n20824, MEM_stage_inst_dmem_n20823, MEM_stage_inst_dmem_n20822, MEM_stage_inst_dmem_n20821, MEM_stage_inst_dmem_n20820, MEM_stage_inst_dmem_n20819, MEM_stage_inst_dmem_n20818, MEM_stage_inst_dmem_n20817, MEM_stage_inst_dmem_n20816, MEM_stage_inst_dmem_n20815, MEM_stage_inst_dmem_n20814, MEM_stage_inst_dmem_n20813, MEM_stage_inst_dmem_n20812, MEM_stage_inst_dmem_n20811, MEM_stage_inst_dmem_n20810, MEM_stage_inst_dmem_n20809, MEM_stage_inst_dmem_n20808, MEM_stage_inst_dmem_n20807, MEM_stage_inst_dmem_n20806, MEM_stage_inst_dmem_n20805, MEM_stage_inst_dmem_n20804, MEM_stage_inst_dmem_n20803, MEM_stage_inst_dmem_n20802, MEM_stage_inst_dmem_n20801, MEM_stage_inst_dmem_n20800, MEM_stage_inst_dmem_n20799, MEM_stage_inst_dmem_n20798, MEM_stage_inst_dmem_n20797, MEM_stage_inst_dmem_n20796, MEM_stage_inst_dmem_n20795, MEM_stage_inst_dmem_n20794, MEM_stage_inst_dmem_n20793, MEM_stage_inst_dmem_n20792, MEM_stage_inst_dmem_n20791, MEM_stage_inst_dmem_n20790, MEM_stage_inst_dmem_n20789, MEM_stage_inst_dmem_n20788, MEM_stage_inst_dmem_n20787, MEM_stage_inst_dmem_n20786, MEM_stage_inst_dmem_n20785, MEM_stage_inst_dmem_n20784, MEM_stage_inst_dmem_n20783, MEM_stage_inst_dmem_n20782, MEM_stage_inst_dmem_n20781, MEM_stage_inst_dmem_n20780, MEM_stage_inst_dmem_n20779, MEM_stage_inst_dmem_n20778, MEM_stage_inst_dmem_n20777, MEM_stage_inst_dmem_n20776, MEM_stage_inst_dmem_n20775, MEM_stage_inst_dmem_n20774, MEM_stage_inst_dmem_n20773, MEM_stage_inst_dmem_n20772, MEM_stage_inst_dmem_n20771, MEM_stage_inst_dmem_n20770, MEM_stage_inst_dmem_n20769, MEM_stage_inst_dmem_n20768, MEM_stage_inst_dmem_n20767, MEM_stage_inst_dmem_n20766, MEM_stage_inst_dmem_n20765, MEM_stage_inst_dmem_n20764, MEM_stage_inst_dmem_n20763, MEM_stage_inst_dmem_n20762, MEM_stage_inst_dmem_n20761, MEM_stage_inst_dmem_n20760, MEM_stage_inst_dmem_n20759, MEM_stage_inst_dmem_n20758, MEM_stage_inst_dmem_n20757, MEM_stage_inst_dmem_n20756, MEM_stage_inst_dmem_n20755, MEM_stage_inst_dmem_n20754, MEM_stage_inst_dmem_n20753, MEM_stage_inst_dmem_n20752, MEM_stage_inst_dmem_n20751, MEM_stage_inst_dmem_n20750, MEM_stage_inst_dmem_n20749, MEM_stage_inst_dmem_n20748, MEM_stage_inst_dmem_n20747, MEM_stage_inst_dmem_n20746, MEM_stage_inst_dmem_n20745, MEM_stage_inst_dmem_n20744, MEM_stage_inst_dmem_n20743, MEM_stage_inst_dmem_n20742, MEM_stage_inst_dmem_n20741, MEM_stage_inst_dmem_n20740, MEM_stage_inst_dmem_n20739, MEM_stage_inst_dmem_n20738, MEM_stage_inst_dmem_n20737, MEM_stage_inst_dmem_n20736, MEM_stage_inst_dmem_n20735, MEM_stage_inst_dmem_n20734, MEM_stage_inst_dmem_n20733, MEM_stage_inst_dmem_n20732, MEM_stage_inst_dmem_n20731, MEM_stage_inst_dmem_n20730, MEM_stage_inst_dmem_n20729, MEM_stage_inst_dmem_n20728, MEM_stage_inst_dmem_n20727, MEM_stage_inst_dmem_n20726, MEM_stage_inst_dmem_n20725, MEM_stage_inst_dmem_n20724, MEM_stage_inst_dmem_n20723, MEM_stage_inst_dmem_n20722, MEM_stage_inst_dmem_n20721, MEM_stage_inst_dmem_n20720, MEM_stage_inst_dmem_n20719, MEM_stage_inst_dmem_n20718, MEM_stage_inst_dmem_n20717, MEM_stage_inst_dmem_n20716, MEM_stage_inst_dmem_n20715, MEM_stage_inst_dmem_n20714, MEM_stage_inst_dmem_n20713, MEM_stage_inst_dmem_n20712, MEM_stage_inst_dmem_n20711, MEM_stage_inst_dmem_n20710, MEM_stage_inst_dmem_n20709, MEM_stage_inst_dmem_n20708, MEM_stage_inst_dmem_n20707, MEM_stage_inst_dmem_n20706, MEM_stage_inst_dmem_n20705, MEM_stage_inst_dmem_n20704, MEM_stage_inst_dmem_n20703, MEM_stage_inst_dmem_n20702, MEM_stage_inst_dmem_n20701, MEM_stage_inst_dmem_n20700, MEM_stage_inst_dmem_n20699, MEM_stage_inst_dmem_n20698, MEM_stage_inst_dmem_n20697, MEM_stage_inst_dmem_n20696, MEM_stage_inst_dmem_n20695, MEM_stage_inst_dmem_n20694, MEM_stage_inst_dmem_n20693, MEM_stage_inst_dmem_n20692, MEM_stage_inst_dmem_n20691, MEM_stage_inst_dmem_n20690, MEM_stage_inst_dmem_n20689, MEM_stage_inst_dmem_n20688, MEM_stage_inst_dmem_n20687, MEM_stage_inst_dmem_n20686, MEM_stage_inst_dmem_n20685, MEM_stage_inst_dmem_n20684, MEM_stage_inst_dmem_n20683, MEM_stage_inst_dmem_n20682, MEM_stage_inst_dmem_n20681, MEM_stage_inst_dmem_n20680, MEM_stage_inst_dmem_n20679, MEM_stage_inst_dmem_n20678, MEM_stage_inst_dmem_n20677, MEM_stage_inst_dmem_n20676, MEM_stage_inst_dmem_n20675, MEM_stage_inst_dmem_n20674, MEM_stage_inst_dmem_n20673, MEM_stage_inst_dmem_n20672, MEM_stage_inst_dmem_n20671, MEM_stage_inst_dmem_n20670, MEM_stage_inst_dmem_n20669, MEM_stage_inst_dmem_n20668, MEM_stage_inst_dmem_n20667, MEM_stage_inst_dmem_n20666, MEM_stage_inst_dmem_n20665, MEM_stage_inst_dmem_n20664, MEM_stage_inst_dmem_n20663, MEM_stage_inst_dmem_n20662, MEM_stage_inst_dmem_n20661, MEM_stage_inst_dmem_n20660, MEM_stage_inst_dmem_n20659, MEM_stage_inst_dmem_n20658, MEM_stage_inst_dmem_n20657, MEM_stage_inst_dmem_n20656, MEM_stage_inst_dmem_n20655, MEM_stage_inst_dmem_n20654, MEM_stage_inst_dmem_n20653, MEM_stage_inst_dmem_n20652, MEM_stage_inst_dmem_n20651, MEM_stage_inst_dmem_n20650, MEM_stage_inst_dmem_n20649, MEM_stage_inst_dmem_n20648, MEM_stage_inst_dmem_n20647, MEM_stage_inst_dmem_n20646, MEM_stage_inst_dmem_n20645, MEM_stage_inst_dmem_n20644, MEM_stage_inst_dmem_n20643, MEM_stage_inst_dmem_n20642, MEM_stage_inst_dmem_n20641, MEM_stage_inst_dmem_n20640, MEM_stage_inst_dmem_n20639, MEM_stage_inst_dmem_n20638, MEM_stage_inst_dmem_n20637, MEM_stage_inst_dmem_n20636, MEM_stage_inst_dmem_n20635, MEM_stage_inst_dmem_n20634, MEM_stage_inst_dmem_n20633, MEM_stage_inst_dmem_n20632, MEM_stage_inst_dmem_n20631, MEM_stage_inst_dmem_n20630, MEM_stage_inst_dmem_n20629, MEM_stage_inst_dmem_n20628, MEM_stage_inst_dmem_n20627, MEM_stage_inst_dmem_n20626, MEM_stage_inst_dmem_n20625, MEM_stage_inst_dmem_n20624, MEM_stage_inst_dmem_n20623, MEM_stage_inst_dmem_n20622, MEM_stage_inst_dmem_n20621, MEM_stage_inst_dmem_n20620, MEM_stage_inst_dmem_n20619, MEM_stage_inst_dmem_n20618, MEM_stage_inst_dmem_n20617, MEM_stage_inst_dmem_n20616, MEM_stage_inst_dmem_n20615, MEM_stage_inst_dmem_n20614, MEM_stage_inst_dmem_n20613, MEM_stage_inst_dmem_n20612, MEM_stage_inst_dmem_n20611, MEM_stage_inst_dmem_n20610, MEM_stage_inst_dmem_n20609, MEM_stage_inst_dmem_n20608, MEM_stage_inst_dmem_n20607, MEM_stage_inst_dmem_n20606, MEM_stage_inst_dmem_n20605, MEM_stage_inst_dmem_n20604, MEM_stage_inst_dmem_n20603, MEM_stage_inst_dmem_n20602, MEM_stage_inst_dmem_n20601, MEM_stage_inst_dmem_n20600, MEM_stage_inst_dmem_n20599, MEM_stage_inst_dmem_n20598, MEM_stage_inst_dmem_n20597, MEM_stage_inst_dmem_n20596, MEM_stage_inst_dmem_n20595, MEM_stage_inst_dmem_n20594, MEM_stage_inst_dmem_n20593, MEM_stage_inst_dmem_n20592, MEM_stage_inst_dmem_n20591, MEM_stage_inst_dmem_n20590, MEM_stage_inst_dmem_n20589, MEM_stage_inst_dmem_n20588, MEM_stage_inst_dmem_n20587, MEM_stage_inst_dmem_n20586, MEM_stage_inst_dmem_n20585, MEM_stage_inst_dmem_n20584, MEM_stage_inst_dmem_n20583, MEM_stage_inst_dmem_n20582, MEM_stage_inst_dmem_n20581, MEM_stage_inst_dmem_n20580, MEM_stage_inst_dmem_n20579, MEM_stage_inst_dmem_n20578, MEM_stage_inst_dmem_n20577, MEM_stage_inst_dmem_n20576, MEM_stage_inst_dmem_n20575, MEM_stage_inst_dmem_n20574, MEM_stage_inst_dmem_n20573, MEM_stage_inst_dmem_n20572, MEM_stage_inst_dmem_n20571, MEM_stage_inst_dmem_n20570, MEM_stage_inst_dmem_n20569, MEM_stage_inst_dmem_n20568, MEM_stage_inst_dmem_n20567, MEM_stage_inst_dmem_n20566, MEM_stage_inst_dmem_n20565, MEM_stage_inst_dmem_n20564, MEM_stage_inst_dmem_n20563, MEM_stage_inst_dmem_n20562, MEM_stage_inst_dmem_n20561, MEM_stage_inst_dmem_n20560, MEM_stage_inst_dmem_n20559, MEM_stage_inst_dmem_n20558, MEM_stage_inst_dmem_n20557, MEM_stage_inst_dmem_n20556, MEM_stage_inst_dmem_n20555, MEM_stage_inst_dmem_n20554, MEM_stage_inst_dmem_n20553, MEM_stage_inst_dmem_n20552, MEM_stage_inst_dmem_n20551, MEM_stage_inst_dmem_n20550, MEM_stage_inst_dmem_n20549, MEM_stage_inst_dmem_n20548, MEM_stage_inst_dmem_n20547, MEM_stage_inst_dmem_n20546, MEM_stage_inst_dmem_n20545, MEM_stage_inst_dmem_n20544, MEM_stage_inst_dmem_n20543, MEM_stage_inst_dmem_n20542, MEM_stage_inst_dmem_n20541, MEM_stage_inst_dmem_n20540, MEM_stage_inst_dmem_n20539, MEM_stage_inst_dmem_n20538, MEM_stage_inst_dmem_n20537, MEM_stage_inst_dmem_n20536, MEM_stage_inst_dmem_n20535, MEM_stage_inst_dmem_n20534, MEM_stage_inst_dmem_n20533, MEM_stage_inst_dmem_n20532, MEM_stage_inst_dmem_n20531, MEM_stage_inst_dmem_n20530, MEM_stage_inst_dmem_n20529, MEM_stage_inst_dmem_n20528, MEM_stage_inst_dmem_n20527, MEM_stage_inst_dmem_n20526, MEM_stage_inst_dmem_n20525, MEM_stage_inst_dmem_n20524, MEM_stage_inst_dmem_n20523, MEM_stage_inst_dmem_n20522, MEM_stage_inst_dmem_n20521, MEM_stage_inst_dmem_n20520, MEM_stage_inst_dmem_n20519, MEM_stage_inst_dmem_n20518, MEM_stage_inst_dmem_n20517, MEM_stage_inst_dmem_n20516, MEM_stage_inst_dmem_n20515, MEM_stage_inst_dmem_n20514, MEM_stage_inst_dmem_n20513, MEM_stage_inst_dmem_n20512, MEM_stage_inst_dmem_n20511, MEM_stage_inst_dmem_n20510, MEM_stage_inst_dmem_n20509, MEM_stage_inst_dmem_n20508, MEM_stage_inst_dmem_n20507, MEM_stage_inst_dmem_n20506, MEM_stage_inst_dmem_n20505, MEM_stage_inst_dmem_n20504, MEM_stage_inst_dmem_n20503, MEM_stage_inst_dmem_n20502, MEM_stage_inst_dmem_n20501, MEM_stage_inst_dmem_n20500, MEM_stage_inst_dmem_n20499, MEM_stage_inst_dmem_n20498, MEM_stage_inst_dmem_n20497, MEM_stage_inst_dmem_n20496, MEM_stage_inst_dmem_n20495, MEM_stage_inst_dmem_n20494, MEM_stage_inst_dmem_n20493, MEM_stage_inst_dmem_n20492, MEM_stage_inst_dmem_n20491, MEM_stage_inst_dmem_n20490, MEM_stage_inst_dmem_n20489, MEM_stage_inst_dmem_n20488, MEM_stage_inst_dmem_n20487, MEM_stage_inst_dmem_n20486, MEM_stage_inst_dmem_n20485, MEM_stage_inst_dmem_n20484, MEM_stage_inst_dmem_n20483, MEM_stage_inst_dmem_n20482, MEM_stage_inst_dmem_n20481, MEM_stage_inst_dmem_n20480, MEM_stage_inst_dmem_n20479, MEM_stage_inst_dmem_n20478, MEM_stage_inst_dmem_n20477, MEM_stage_inst_dmem_n20476, MEM_stage_inst_dmem_n20475, MEM_stage_inst_dmem_n20474, MEM_stage_inst_dmem_n20473, MEM_stage_inst_dmem_n20472, MEM_stage_inst_dmem_n20471, MEM_stage_inst_dmem_n20470, MEM_stage_inst_dmem_n20469, MEM_stage_inst_dmem_n20468, MEM_stage_inst_dmem_n20467, MEM_stage_inst_dmem_n20466, MEM_stage_inst_dmem_n20465, MEM_stage_inst_dmem_n20464, MEM_stage_inst_dmem_n20463, MEM_stage_inst_dmem_n20462, MEM_stage_inst_dmem_n20461, MEM_stage_inst_dmem_n20460, MEM_stage_inst_dmem_n20459, MEM_stage_inst_dmem_n20458, MEM_stage_inst_dmem_n20457, MEM_stage_inst_dmem_n20456, MEM_stage_inst_dmem_n20455, MEM_stage_inst_dmem_n20454, MEM_stage_inst_dmem_n20453, MEM_stage_inst_dmem_n20452, MEM_stage_inst_dmem_n20451, MEM_stage_inst_dmem_n20450, MEM_stage_inst_dmem_n20449, MEM_stage_inst_dmem_n20448, MEM_stage_inst_dmem_n20447, MEM_stage_inst_dmem_n20446, MEM_stage_inst_dmem_n20445, MEM_stage_inst_dmem_n20444, MEM_stage_inst_dmem_n20443, MEM_stage_inst_dmem_n20442, MEM_stage_inst_dmem_n20441, MEM_stage_inst_dmem_n20440, MEM_stage_inst_dmem_n20439, MEM_stage_inst_dmem_n20438, MEM_stage_inst_dmem_n20437, MEM_stage_inst_dmem_n20436, MEM_stage_inst_dmem_n20435, MEM_stage_inst_dmem_n20434, MEM_stage_inst_dmem_n20433, MEM_stage_inst_dmem_n20432, MEM_stage_inst_dmem_n20431, MEM_stage_inst_dmem_n20430, MEM_stage_inst_dmem_n20429, MEM_stage_inst_dmem_n20428, MEM_stage_inst_dmem_n20427, MEM_stage_inst_dmem_n20426, MEM_stage_inst_dmem_n20425, MEM_stage_inst_dmem_n20424, MEM_stage_inst_dmem_n20423, MEM_stage_inst_dmem_n20422, MEM_stage_inst_dmem_n20421, MEM_stage_inst_dmem_n20420, MEM_stage_inst_dmem_n20419, MEM_stage_inst_dmem_n20418, MEM_stage_inst_dmem_n20417, MEM_stage_inst_dmem_n20416, MEM_stage_inst_dmem_n20415, MEM_stage_inst_dmem_n20414, MEM_stage_inst_dmem_n20413, MEM_stage_inst_dmem_n20412, MEM_stage_inst_dmem_n20411, MEM_stage_inst_dmem_n20410, MEM_stage_inst_dmem_n20409, MEM_stage_inst_dmem_n20408, MEM_stage_inst_dmem_n20407, MEM_stage_inst_dmem_n20406, MEM_stage_inst_dmem_n20405, MEM_stage_inst_dmem_n20404, MEM_stage_inst_dmem_n20403, MEM_stage_inst_dmem_n20402, MEM_stage_inst_dmem_n20401, MEM_stage_inst_dmem_n20400, MEM_stage_inst_dmem_n20399, MEM_stage_inst_dmem_n20398, MEM_stage_inst_dmem_n20397, MEM_stage_inst_dmem_n20396, MEM_stage_inst_dmem_n20395, MEM_stage_inst_dmem_n20394, MEM_stage_inst_dmem_n20393, MEM_stage_inst_dmem_n20392, MEM_stage_inst_dmem_n20391, MEM_stage_inst_dmem_n20390, MEM_stage_inst_dmem_n20389, MEM_stage_inst_dmem_n20388, MEM_stage_inst_dmem_n20387, MEM_stage_inst_dmem_n20386, MEM_stage_inst_dmem_n20385, MEM_stage_inst_dmem_n20384, MEM_stage_inst_dmem_n20383, MEM_stage_inst_dmem_n20382, MEM_stage_inst_dmem_n20381, MEM_stage_inst_dmem_n20380, MEM_stage_inst_dmem_n20379, MEM_stage_inst_dmem_n20378, MEM_stage_inst_dmem_n20377, MEM_stage_inst_dmem_n20376, MEM_stage_inst_dmem_n20375, MEM_stage_inst_dmem_n20374, MEM_stage_inst_dmem_n20373, MEM_stage_inst_dmem_n20372, MEM_stage_inst_dmem_n20371, MEM_stage_inst_dmem_n20370, MEM_stage_inst_dmem_n20369, MEM_stage_inst_dmem_n20368, MEM_stage_inst_dmem_n20367, MEM_stage_inst_dmem_n20366, MEM_stage_inst_dmem_n20365, MEM_stage_inst_dmem_n20364, MEM_stage_inst_dmem_n20363, MEM_stage_inst_dmem_n20362, MEM_stage_inst_dmem_n20361, MEM_stage_inst_dmem_n20360, MEM_stage_inst_dmem_n20359, MEM_stage_inst_dmem_n20358, MEM_stage_inst_dmem_n20357, MEM_stage_inst_dmem_n20356, MEM_stage_inst_dmem_n20355, MEM_stage_inst_dmem_n20354, MEM_stage_inst_dmem_n20353, MEM_stage_inst_dmem_n20352, MEM_stage_inst_dmem_n20351, MEM_stage_inst_dmem_n20350, MEM_stage_inst_dmem_n20349, MEM_stage_inst_dmem_n20348, MEM_stage_inst_dmem_n20347, MEM_stage_inst_dmem_n20346, MEM_stage_inst_dmem_n20345, MEM_stage_inst_dmem_n20344, MEM_stage_inst_dmem_n20343, MEM_stage_inst_dmem_n20342, MEM_stage_inst_dmem_n20341, MEM_stage_inst_dmem_n20340, MEM_stage_inst_dmem_n20339, MEM_stage_inst_dmem_n20338, MEM_stage_inst_dmem_n20337, MEM_stage_inst_dmem_n20336, MEM_stage_inst_dmem_n20335, MEM_stage_inst_dmem_n20334, MEM_stage_inst_dmem_n20333, MEM_stage_inst_dmem_n20332, MEM_stage_inst_dmem_n20331, MEM_stage_inst_dmem_n20330, MEM_stage_inst_dmem_n20329, MEM_stage_inst_dmem_n20328, MEM_stage_inst_dmem_n20327, MEM_stage_inst_dmem_n20326, MEM_stage_inst_dmem_n20325, MEM_stage_inst_dmem_n20324, MEM_stage_inst_dmem_n20323, MEM_stage_inst_dmem_n20322, MEM_stage_inst_dmem_n20321, MEM_stage_inst_dmem_n20320, MEM_stage_inst_dmem_n20319, MEM_stage_inst_dmem_n20318, MEM_stage_inst_dmem_n20317, MEM_stage_inst_dmem_n20316, MEM_stage_inst_dmem_n20315, MEM_stage_inst_dmem_n20314, MEM_stage_inst_dmem_n20313, MEM_stage_inst_dmem_n20312, MEM_stage_inst_dmem_n20311, MEM_stage_inst_dmem_n20310, MEM_stage_inst_dmem_n20309, MEM_stage_inst_dmem_n20308, MEM_stage_inst_dmem_n20307, MEM_stage_inst_dmem_n20306, MEM_stage_inst_dmem_n20305, MEM_stage_inst_dmem_n20304, MEM_stage_inst_dmem_n20303, MEM_stage_inst_dmem_n20302, MEM_stage_inst_dmem_n20301, MEM_stage_inst_dmem_n20300, MEM_stage_inst_dmem_n20299, MEM_stage_inst_dmem_n20298, MEM_stage_inst_dmem_n20297, MEM_stage_inst_dmem_n20296, MEM_stage_inst_dmem_n20295, MEM_stage_inst_dmem_n20294, MEM_stage_inst_dmem_n20293, MEM_stage_inst_dmem_n20292, MEM_stage_inst_dmem_n20291, MEM_stage_inst_dmem_n20290, MEM_stage_inst_dmem_n20289, MEM_stage_inst_dmem_n20288, MEM_stage_inst_dmem_n20287, MEM_stage_inst_dmem_n20286, MEM_stage_inst_dmem_n20285, MEM_stage_inst_dmem_n20284, MEM_stage_inst_dmem_n20283, MEM_stage_inst_dmem_n20282, MEM_stage_inst_dmem_n20281, MEM_stage_inst_dmem_n20280, MEM_stage_inst_dmem_n20279, MEM_stage_inst_dmem_n20278, MEM_stage_inst_dmem_n20277, MEM_stage_inst_dmem_n20276, MEM_stage_inst_dmem_n20275, MEM_stage_inst_dmem_n20274, MEM_stage_inst_dmem_n20273, MEM_stage_inst_dmem_n20272, MEM_stage_inst_dmem_n20271, MEM_stage_inst_dmem_n20270, MEM_stage_inst_dmem_n20269, MEM_stage_inst_dmem_n20268, MEM_stage_inst_dmem_n20267, MEM_stage_inst_dmem_n20266, MEM_stage_inst_dmem_n20265, MEM_stage_inst_dmem_n20264, MEM_stage_inst_dmem_n20263, MEM_stage_inst_dmem_n20262, MEM_stage_inst_dmem_n20261, MEM_stage_inst_dmem_n20260, MEM_stage_inst_dmem_n20259, MEM_stage_inst_dmem_n20258, MEM_stage_inst_dmem_n20257, MEM_stage_inst_dmem_n20256, MEM_stage_inst_dmem_n20255, MEM_stage_inst_dmem_n20254, MEM_stage_inst_dmem_n20253, MEM_stage_inst_dmem_n20252, MEM_stage_inst_dmem_n20251, MEM_stage_inst_dmem_n20250, MEM_stage_inst_dmem_n20249, MEM_stage_inst_dmem_n20248, MEM_stage_inst_dmem_n20247, MEM_stage_inst_dmem_n20246, MEM_stage_inst_dmem_n20245, MEM_stage_inst_dmem_n20244, MEM_stage_inst_dmem_n20243, MEM_stage_inst_dmem_n20242, MEM_stage_inst_dmem_n20241, MEM_stage_inst_dmem_n20240, MEM_stage_inst_dmem_n20239, MEM_stage_inst_dmem_n20238, MEM_stage_inst_dmem_n20237, MEM_stage_inst_dmem_n20236, MEM_stage_inst_dmem_n20235, MEM_stage_inst_dmem_n20234, MEM_stage_inst_dmem_n20233, MEM_stage_inst_dmem_n20232, MEM_stage_inst_dmem_n20231, MEM_stage_inst_dmem_n20230, MEM_stage_inst_dmem_n20229, MEM_stage_inst_dmem_n20228, MEM_stage_inst_dmem_n20227, MEM_stage_inst_dmem_n20226, MEM_stage_inst_dmem_n20225, MEM_stage_inst_dmem_n20224, MEM_stage_inst_dmem_n20223, MEM_stage_inst_dmem_n20222, MEM_stage_inst_dmem_n20221, MEM_stage_inst_dmem_n20220, MEM_stage_inst_dmem_n20219, MEM_stage_inst_dmem_n20218, MEM_stage_inst_dmem_n20217, MEM_stage_inst_dmem_n20216, MEM_stage_inst_dmem_n20215, MEM_stage_inst_dmem_n20214, MEM_stage_inst_dmem_n20213, MEM_stage_inst_dmem_n20212, MEM_stage_inst_dmem_n20211, MEM_stage_inst_dmem_n20210, MEM_stage_inst_dmem_n20209, MEM_stage_inst_dmem_n20208, MEM_stage_inst_dmem_n20207, MEM_stage_inst_dmem_n20206, MEM_stage_inst_dmem_n20205, MEM_stage_inst_dmem_n20204, MEM_stage_inst_dmem_n20203, MEM_stage_inst_dmem_n20202, MEM_stage_inst_dmem_n20201, MEM_stage_inst_dmem_n20200, MEM_stage_inst_dmem_n20199, MEM_stage_inst_dmem_n20198, MEM_stage_inst_dmem_n20197, MEM_stage_inst_dmem_n20196, MEM_stage_inst_dmem_n20195, MEM_stage_inst_dmem_n20194, MEM_stage_inst_dmem_n20193, MEM_stage_inst_dmem_n20192, MEM_stage_inst_dmem_n20191, MEM_stage_inst_dmem_n20190, MEM_stage_inst_dmem_n20189, MEM_stage_inst_dmem_n20188, MEM_stage_inst_dmem_n20187, MEM_stage_inst_dmem_n20186, MEM_stage_inst_dmem_n20185, MEM_stage_inst_dmem_n20184, MEM_stage_inst_dmem_n20183, MEM_stage_inst_dmem_n20182, MEM_stage_inst_dmem_n20181, MEM_stage_inst_dmem_n20180, MEM_stage_inst_dmem_n20179, MEM_stage_inst_dmem_n20178, MEM_stage_inst_dmem_n20177, MEM_stage_inst_dmem_n20176, MEM_stage_inst_dmem_n20175, MEM_stage_inst_dmem_n20174, MEM_stage_inst_dmem_n20173, MEM_stage_inst_dmem_n20172, MEM_stage_inst_dmem_n20171, MEM_stage_inst_dmem_n20170, MEM_stage_inst_dmem_n20169, MEM_stage_inst_dmem_n20168, MEM_stage_inst_dmem_n20167, MEM_stage_inst_dmem_n20166, MEM_stage_inst_dmem_n20165, MEM_stage_inst_dmem_n20164, MEM_stage_inst_dmem_n20163, MEM_stage_inst_dmem_n20162, MEM_stage_inst_dmem_n20161, MEM_stage_inst_dmem_n20160, MEM_stage_inst_dmem_n20159, MEM_stage_inst_dmem_n20158, MEM_stage_inst_dmem_n20157, MEM_stage_inst_dmem_n20156, MEM_stage_inst_dmem_n20155, MEM_stage_inst_dmem_n20154, MEM_stage_inst_dmem_n20153, MEM_stage_inst_dmem_n20152, MEM_stage_inst_dmem_n20151, MEM_stage_inst_dmem_n20150, MEM_stage_inst_dmem_n20149, MEM_stage_inst_dmem_n20148, MEM_stage_inst_dmem_n20147, MEM_stage_inst_dmem_n20146, MEM_stage_inst_dmem_n20145, MEM_stage_inst_dmem_n20144, MEM_stage_inst_dmem_n20143, MEM_stage_inst_dmem_n20142, MEM_stage_inst_dmem_n20141, MEM_stage_inst_dmem_n20140, MEM_stage_inst_dmem_n20139, MEM_stage_inst_dmem_n20138, MEM_stage_inst_dmem_n20137, MEM_stage_inst_dmem_n20136, MEM_stage_inst_dmem_n20135, MEM_stage_inst_dmem_n20134, MEM_stage_inst_dmem_n20133, MEM_stage_inst_dmem_n20132, MEM_stage_inst_dmem_n20131, MEM_stage_inst_dmem_n20130, MEM_stage_inst_dmem_n20129, MEM_stage_inst_dmem_n20128, MEM_stage_inst_dmem_n20127, MEM_stage_inst_dmem_n20126, MEM_stage_inst_dmem_n20125, MEM_stage_inst_dmem_n20124, MEM_stage_inst_dmem_n20123, MEM_stage_inst_dmem_n20122, MEM_stage_inst_dmem_n20121, MEM_stage_inst_dmem_n20120, MEM_stage_inst_dmem_n20119, MEM_stage_inst_dmem_n20118, MEM_stage_inst_dmem_n20117, MEM_stage_inst_dmem_n20116, MEM_stage_inst_dmem_n20115, MEM_stage_inst_dmem_n20114, MEM_stage_inst_dmem_n20113, MEM_stage_inst_dmem_n20112, MEM_stage_inst_dmem_n20111, MEM_stage_inst_dmem_n20110, MEM_stage_inst_dmem_n20109, MEM_stage_inst_dmem_n20108, MEM_stage_inst_dmem_n20107, MEM_stage_inst_dmem_n20106, MEM_stage_inst_dmem_n20105, MEM_stage_inst_dmem_n20104, MEM_stage_inst_dmem_n20103, MEM_stage_inst_dmem_n20102, MEM_stage_inst_dmem_n20101, MEM_stage_inst_dmem_n20100, MEM_stage_inst_dmem_n20099, MEM_stage_inst_dmem_n20098, MEM_stage_inst_dmem_n20097, MEM_stage_inst_dmem_n20096, MEM_stage_inst_dmem_n20095, MEM_stage_inst_dmem_n20094, MEM_stage_inst_dmem_n20093, MEM_stage_inst_dmem_n20092, MEM_stage_inst_dmem_n20091, MEM_stage_inst_dmem_n20090, MEM_stage_inst_dmem_n20089, MEM_stage_inst_dmem_n20088, MEM_stage_inst_dmem_n20087, MEM_stage_inst_dmem_n20086, MEM_stage_inst_dmem_n20085, MEM_stage_inst_dmem_n20084, MEM_stage_inst_dmem_n20083, MEM_stage_inst_dmem_n20082, MEM_stage_inst_dmem_n20081, MEM_stage_inst_dmem_n20080, MEM_stage_inst_dmem_n20079, MEM_stage_inst_dmem_n20078, MEM_stage_inst_dmem_n20077, MEM_stage_inst_dmem_n20076, MEM_stage_inst_dmem_n20075, MEM_stage_inst_dmem_n20074, MEM_stage_inst_dmem_n20073, MEM_stage_inst_dmem_n20072, MEM_stage_inst_dmem_n20071, MEM_stage_inst_dmem_n20070, MEM_stage_inst_dmem_n20069, MEM_stage_inst_dmem_n20068, MEM_stage_inst_dmem_n20067, MEM_stage_inst_dmem_n20066, MEM_stage_inst_dmem_n20065, MEM_stage_inst_dmem_n20064, MEM_stage_inst_dmem_n20063, MEM_stage_inst_dmem_n20062, MEM_stage_inst_dmem_n20061, MEM_stage_inst_dmem_n20060, MEM_stage_inst_dmem_n20059, MEM_stage_inst_dmem_n20058, MEM_stage_inst_dmem_n20057, MEM_stage_inst_dmem_n20056, MEM_stage_inst_dmem_n20055, MEM_stage_inst_dmem_n20054, MEM_stage_inst_dmem_n20053, MEM_stage_inst_dmem_n20052, MEM_stage_inst_dmem_n20051, MEM_stage_inst_dmem_n20050, MEM_stage_inst_dmem_n20049, MEM_stage_inst_dmem_n20048, MEM_stage_inst_dmem_n20047, MEM_stage_inst_dmem_n20046, MEM_stage_inst_dmem_n20045, MEM_stage_inst_dmem_n20044, MEM_stage_inst_dmem_n20043, MEM_stage_inst_dmem_n20042, MEM_stage_inst_dmem_n20041, MEM_stage_inst_dmem_n20040, MEM_stage_inst_dmem_n20039, MEM_stage_inst_dmem_n20038, MEM_stage_inst_dmem_n20037, MEM_stage_inst_dmem_n20036, MEM_stage_inst_dmem_n20035, MEM_stage_inst_dmem_n20034, MEM_stage_inst_dmem_n20033, MEM_stage_inst_dmem_n20032, MEM_stage_inst_dmem_n20031, MEM_stage_inst_dmem_n20030, MEM_stage_inst_dmem_n20029, MEM_stage_inst_dmem_n20028, MEM_stage_inst_dmem_n20027, MEM_stage_inst_dmem_n20026, MEM_stage_inst_dmem_n20025, MEM_stage_inst_dmem_n20024, MEM_stage_inst_dmem_n20023, MEM_stage_inst_dmem_n20022, MEM_stage_inst_dmem_n20021, MEM_stage_inst_dmem_n20020, MEM_stage_inst_dmem_n20019, MEM_stage_inst_dmem_n20018, MEM_stage_inst_dmem_n20017, MEM_stage_inst_dmem_n20016, MEM_stage_inst_dmem_n20015, MEM_stage_inst_dmem_n20014, MEM_stage_inst_dmem_n20013, MEM_stage_inst_dmem_n20012, MEM_stage_inst_dmem_n20011, MEM_stage_inst_dmem_n20010, MEM_stage_inst_dmem_n20009, MEM_stage_inst_dmem_n20008, MEM_stage_inst_dmem_n20007, MEM_stage_inst_dmem_n20006, MEM_stage_inst_dmem_n20005, MEM_stage_inst_dmem_n20004, MEM_stage_inst_dmem_n20003, MEM_stage_inst_dmem_n20002, MEM_stage_inst_dmem_n20001, MEM_stage_inst_dmem_n20000, MEM_stage_inst_dmem_n19999, MEM_stage_inst_dmem_n19998, MEM_stage_inst_dmem_n19997, MEM_stage_inst_dmem_n19996, MEM_stage_inst_dmem_n19995, MEM_stage_inst_dmem_n19994, MEM_stage_inst_dmem_n19993, MEM_stage_inst_dmem_n19992, MEM_stage_inst_dmem_n19991, MEM_stage_inst_dmem_n19990, MEM_stage_inst_dmem_n19989, MEM_stage_inst_dmem_n19988, MEM_stage_inst_dmem_n19987, MEM_stage_inst_dmem_n19986, MEM_stage_inst_dmem_n19985, MEM_stage_inst_dmem_n19984, MEM_stage_inst_dmem_n19983, MEM_stage_inst_dmem_n19982, MEM_stage_inst_dmem_n19981, MEM_stage_inst_dmem_n19980, MEM_stage_inst_dmem_n19979, MEM_stage_inst_dmem_n19978, MEM_stage_inst_dmem_n19977, MEM_stage_inst_dmem_n19976, MEM_stage_inst_dmem_n19975, MEM_stage_inst_dmem_n19974, MEM_stage_inst_dmem_n19973, MEM_stage_inst_dmem_n19972, MEM_stage_inst_dmem_n19971, MEM_stage_inst_dmem_n19970, MEM_stage_inst_dmem_n19969, MEM_stage_inst_dmem_n19968, MEM_stage_inst_dmem_n19967, MEM_stage_inst_dmem_n19966, MEM_stage_inst_dmem_n19965, MEM_stage_inst_dmem_n19964, MEM_stage_inst_dmem_n19963, MEM_stage_inst_dmem_n19962, MEM_stage_inst_dmem_n19961, MEM_stage_inst_dmem_n19960, MEM_stage_inst_dmem_n19959, MEM_stage_inst_dmem_n19958, MEM_stage_inst_dmem_n19957, MEM_stage_inst_dmem_n19956, MEM_stage_inst_dmem_n19955, MEM_stage_inst_dmem_n19954, MEM_stage_inst_dmem_n19953, MEM_stage_inst_dmem_n19952, MEM_stage_inst_dmem_n19951, MEM_stage_inst_dmem_n19950, MEM_stage_inst_dmem_n19949, MEM_stage_inst_dmem_n19948, MEM_stage_inst_dmem_n19947, MEM_stage_inst_dmem_n19946, MEM_stage_inst_dmem_n19945, MEM_stage_inst_dmem_n19944, MEM_stage_inst_dmem_n19943, MEM_stage_inst_dmem_n19942, MEM_stage_inst_dmem_n19941, MEM_stage_inst_dmem_n19940, MEM_stage_inst_dmem_n19939, MEM_stage_inst_dmem_n19938, MEM_stage_inst_dmem_n19937, MEM_stage_inst_dmem_n19936, MEM_stage_inst_dmem_n19935, MEM_stage_inst_dmem_n19934, MEM_stage_inst_dmem_n19933, MEM_stage_inst_dmem_n19932, MEM_stage_inst_dmem_n19931, MEM_stage_inst_dmem_n19930, MEM_stage_inst_dmem_n19929, MEM_stage_inst_dmem_n19928, MEM_stage_inst_dmem_n19927, MEM_stage_inst_dmem_n19926, MEM_stage_inst_dmem_n19925, MEM_stage_inst_dmem_n19924, MEM_stage_inst_dmem_n19923, MEM_stage_inst_dmem_n19922, MEM_stage_inst_dmem_n19921, MEM_stage_inst_dmem_n19920, MEM_stage_inst_dmem_n19919, MEM_stage_inst_dmem_n19918, MEM_stage_inst_dmem_n19917, MEM_stage_inst_dmem_n19916, MEM_stage_inst_dmem_n19915, MEM_stage_inst_dmem_n19914, MEM_stage_inst_dmem_n19913, MEM_stage_inst_dmem_n19912, MEM_stage_inst_dmem_n19911, MEM_stage_inst_dmem_n19910, MEM_stage_inst_dmem_n19909, MEM_stage_inst_dmem_n19908, MEM_stage_inst_dmem_n19907, MEM_stage_inst_dmem_n19906, MEM_stage_inst_dmem_n19905, MEM_stage_inst_dmem_n19904, MEM_stage_inst_dmem_n19903, MEM_stage_inst_dmem_n19902, MEM_stage_inst_dmem_n19901, MEM_stage_inst_dmem_n19900, MEM_stage_inst_dmem_n19899, MEM_stage_inst_dmem_n19898, MEM_stage_inst_dmem_n19897, MEM_stage_inst_dmem_n19896, MEM_stage_inst_dmem_n19895, MEM_stage_inst_dmem_n19894, MEM_stage_inst_dmem_n19893, MEM_stage_inst_dmem_n19892, MEM_stage_inst_dmem_n19891, MEM_stage_inst_dmem_n19890, MEM_stage_inst_dmem_n19889, MEM_stage_inst_dmem_n19888, MEM_stage_inst_dmem_n19887, MEM_stage_inst_dmem_n19886, MEM_stage_inst_dmem_n19885, MEM_stage_inst_dmem_n19884, MEM_stage_inst_dmem_n19883, MEM_stage_inst_dmem_n19882, MEM_stage_inst_dmem_n19881, MEM_stage_inst_dmem_n19880, MEM_stage_inst_dmem_n19879, MEM_stage_inst_dmem_n19878, MEM_stage_inst_dmem_n19877, MEM_stage_inst_dmem_n19876, MEM_stage_inst_dmem_n19875, MEM_stage_inst_dmem_n19874, MEM_stage_inst_dmem_n19873, MEM_stage_inst_dmem_n19872, MEM_stage_inst_dmem_n19871, MEM_stage_inst_dmem_n19870, MEM_stage_inst_dmem_n19869, MEM_stage_inst_dmem_n19868, MEM_stage_inst_dmem_n19867, MEM_stage_inst_dmem_n19866, MEM_stage_inst_dmem_n19865, MEM_stage_inst_dmem_n19864, MEM_stage_inst_dmem_n19863, MEM_stage_inst_dmem_n19862, MEM_stage_inst_dmem_n19861, MEM_stage_inst_dmem_n19860, MEM_stage_inst_dmem_n19859, MEM_stage_inst_dmem_n19858, MEM_stage_inst_dmem_n19857, MEM_stage_inst_dmem_n19856, MEM_stage_inst_dmem_n19855, MEM_stage_inst_dmem_n19854, MEM_stage_inst_dmem_n19853, MEM_stage_inst_dmem_n19852, MEM_stage_inst_dmem_n19851, MEM_stage_inst_dmem_n19850, MEM_stage_inst_dmem_n19849, MEM_stage_inst_dmem_n19848, MEM_stage_inst_dmem_n19847, MEM_stage_inst_dmem_n19846, MEM_stage_inst_dmem_n19845, MEM_stage_inst_dmem_n19844, MEM_stage_inst_dmem_n19843, MEM_stage_inst_dmem_n19842, MEM_stage_inst_dmem_n19841, MEM_stage_inst_dmem_n19840, MEM_stage_inst_dmem_n19839, MEM_stage_inst_dmem_n19838, MEM_stage_inst_dmem_n19837, MEM_stage_inst_dmem_n19836, MEM_stage_inst_dmem_n19835, MEM_stage_inst_dmem_n19834, MEM_stage_inst_dmem_n19833, MEM_stage_inst_dmem_n19832, MEM_stage_inst_dmem_n19831, MEM_stage_inst_dmem_n19830, MEM_stage_inst_dmem_n19829, MEM_stage_inst_dmem_n19828, MEM_stage_inst_dmem_n19827, MEM_stage_inst_dmem_n19826, MEM_stage_inst_dmem_n19825, MEM_stage_inst_dmem_n19824, MEM_stage_inst_dmem_n19823, MEM_stage_inst_dmem_n19822, MEM_stage_inst_dmem_n19821, MEM_stage_inst_dmem_n19820, MEM_stage_inst_dmem_n19819, MEM_stage_inst_dmem_n19818, MEM_stage_inst_dmem_n19817, MEM_stage_inst_dmem_n19816, MEM_stage_inst_dmem_n19815, MEM_stage_inst_dmem_n19814, MEM_stage_inst_dmem_n19813, MEM_stage_inst_dmem_n19812, MEM_stage_inst_dmem_n19811, MEM_stage_inst_dmem_n19810, MEM_stage_inst_dmem_n19809, MEM_stage_inst_dmem_n19808, MEM_stage_inst_dmem_n19807, MEM_stage_inst_dmem_n19806, MEM_stage_inst_dmem_n19805, MEM_stage_inst_dmem_n19804, MEM_stage_inst_dmem_n19803, MEM_stage_inst_dmem_n19802, MEM_stage_inst_dmem_n19801, MEM_stage_inst_dmem_n19800, MEM_stage_inst_dmem_n19799, MEM_stage_inst_dmem_n19798, MEM_stage_inst_dmem_n19797, MEM_stage_inst_dmem_n19796, MEM_stage_inst_dmem_n19795, MEM_stage_inst_dmem_n19794, MEM_stage_inst_dmem_n19793, MEM_stage_inst_dmem_n19792, MEM_stage_inst_dmem_n19791, MEM_stage_inst_dmem_n19790, MEM_stage_inst_dmem_n19789, MEM_stage_inst_dmem_n19788, MEM_stage_inst_dmem_n19787, MEM_stage_inst_dmem_n19786, MEM_stage_inst_dmem_n19785, MEM_stage_inst_dmem_n19784, MEM_stage_inst_dmem_n19783, MEM_stage_inst_dmem_n19782, MEM_stage_inst_dmem_n19781, MEM_stage_inst_dmem_n19780, MEM_stage_inst_dmem_n19779, MEM_stage_inst_dmem_n19778, MEM_stage_inst_dmem_n19777, MEM_stage_inst_dmem_n19776, MEM_stage_inst_dmem_n19775, MEM_stage_inst_dmem_n19774, MEM_stage_inst_dmem_n19773, MEM_stage_inst_dmem_n19772, MEM_stage_inst_dmem_n19771, MEM_stage_inst_dmem_n19770, MEM_stage_inst_dmem_n19769, MEM_stage_inst_dmem_n19768, MEM_stage_inst_dmem_n19767, MEM_stage_inst_dmem_n19766, MEM_stage_inst_dmem_n19765, MEM_stage_inst_dmem_n19764, MEM_stage_inst_dmem_n19763, MEM_stage_inst_dmem_n19762, MEM_stage_inst_dmem_n19761, MEM_stage_inst_dmem_n19760, MEM_stage_inst_dmem_n19759, MEM_stage_inst_dmem_n19758, MEM_stage_inst_dmem_n19757, MEM_stage_inst_dmem_n19756, MEM_stage_inst_dmem_n19755, MEM_stage_inst_dmem_n19754, MEM_stage_inst_dmem_n19753, MEM_stage_inst_dmem_n19752, MEM_stage_inst_dmem_n19751, MEM_stage_inst_dmem_n19750, MEM_stage_inst_dmem_n19749, MEM_stage_inst_dmem_n19748, MEM_stage_inst_dmem_n19747, MEM_stage_inst_dmem_n19746, MEM_stage_inst_dmem_n19745, MEM_stage_inst_dmem_n19744, MEM_stage_inst_dmem_n19743, MEM_stage_inst_dmem_n19742, MEM_stage_inst_dmem_n19741, MEM_stage_inst_dmem_n19740, MEM_stage_inst_dmem_n19739, MEM_stage_inst_dmem_n19738, MEM_stage_inst_dmem_n19737, MEM_stage_inst_dmem_n19736, MEM_stage_inst_dmem_n19735, MEM_stage_inst_dmem_n19734, MEM_stage_inst_dmem_n19733, MEM_stage_inst_dmem_n19732, MEM_stage_inst_dmem_n19731, MEM_stage_inst_dmem_n19730, MEM_stage_inst_dmem_n19729, MEM_stage_inst_dmem_n19728, MEM_stage_inst_dmem_n19727, MEM_stage_inst_dmem_n19726, MEM_stage_inst_dmem_n19725, MEM_stage_inst_dmem_n19724, MEM_stage_inst_dmem_n19723, MEM_stage_inst_dmem_n19722, MEM_stage_inst_dmem_n19721, MEM_stage_inst_dmem_n19720, MEM_stage_inst_dmem_n19719, MEM_stage_inst_dmem_n19718, MEM_stage_inst_dmem_n19717, MEM_stage_inst_dmem_n19716, MEM_stage_inst_dmem_n19715, MEM_stage_inst_dmem_n19714, MEM_stage_inst_dmem_n19713, MEM_stage_inst_dmem_n19712, MEM_stage_inst_dmem_n19711, MEM_stage_inst_dmem_n19710, MEM_stage_inst_dmem_n19709, MEM_stage_inst_dmem_n19708, MEM_stage_inst_dmem_n19707, MEM_stage_inst_dmem_n19706, MEM_stage_inst_dmem_n19705, MEM_stage_inst_dmem_n19704, MEM_stage_inst_dmem_n19703, MEM_stage_inst_dmem_n19702, MEM_stage_inst_dmem_n19701, MEM_stage_inst_dmem_n19700, MEM_stage_inst_dmem_n19699, MEM_stage_inst_dmem_n19698, MEM_stage_inst_dmem_n19697, MEM_stage_inst_dmem_n19696, MEM_stage_inst_dmem_n19695, MEM_stage_inst_dmem_n19694, MEM_stage_inst_dmem_n19693, MEM_stage_inst_dmem_n19692, MEM_stage_inst_dmem_n19691, MEM_stage_inst_dmem_n19690, MEM_stage_inst_dmem_n19689, MEM_stage_inst_dmem_n19688, MEM_stage_inst_dmem_n19687, MEM_stage_inst_dmem_n19686, MEM_stage_inst_dmem_n19685, MEM_stage_inst_dmem_n19684, MEM_stage_inst_dmem_n19683, MEM_stage_inst_dmem_n19682, MEM_stage_inst_dmem_n19681, MEM_stage_inst_dmem_n19680, MEM_stage_inst_dmem_n19679, MEM_stage_inst_dmem_n19678, MEM_stage_inst_dmem_n19677, MEM_stage_inst_dmem_n19676, MEM_stage_inst_dmem_n19675, MEM_stage_inst_dmem_n19674, MEM_stage_inst_dmem_n19673, MEM_stage_inst_dmem_n19672, MEM_stage_inst_dmem_n19671, MEM_stage_inst_dmem_n19670, MEM_stage_inst_dmem_n19669, MEM_stage_inst_dmem_n19668, MEM_stage_inst_dmem_n19667, MEM_stage_inst_dmem_n19666, MEM_stage_inst_dmem_n19665, MEM_stage_inst_dmem_n19664, MEM_stage_inst_dmem_n19663, MEM_stage_inst_dmem_n19662, MEM_stage_inst_dmem_n19661, MEM_stage_inst_dmem_n19660, MEM_stage_inst_dmem_n19659, MEM_stage_inst_dmem_n19658, MEM_stage_inst_dmem_n19657, MEM_stage_inst_dmem_n19656, MEM_stage_inst_dmem_n19655, MEM_stage_inst_dmem_n19654, MEM_stage_inst_dmem_n19653, MEM_stage_inst_dmem_n19652, MEM_stage_inst_dmem_n19651, MEM_stage_inst_dmem_n19650, MEM_stage_inst_dmem_n19649, MEM_stage_inst_dmem_n19648, MEM_stage_inst_dmem_n19647, MEM_stage_inst_dmem_n19646, MEM_stage_inst_dmem_n19645, MEM_stage_inst_dmem_n19644, MEM_stage_inst_dmem_n19643, MEM_stage_inst_dmem_n19642, MEM_stage_inst_dmem_n19641, MEM_stage_inst_dmem_n19640, MEM_stage_inst_dmem_n19639, MEM_stage_inst_dmem_n19638, MEM_stage_inst_dmem_n19637, MEM_stage_inst_dmem_n19636, MEM_stage_inst_dmem_n19635, MEM_stage_inst_dmem_n19634, MEM_stage_inst_dmem_n19633, MEM_stage_inst_dmem_n19632, MEM_stage_inst_dmem_n19631, MEM_stage_inst_dmem_n19630, MEM_stage_inst_dmem_n19629, MEM_stage_inst_dmem_n19628, MEM_stage_inst_dmem_n19627, MEM_stage_inst_dmem_n19626, MEM_stage_inst_dmem_n19625, MEM_stage_inst_dmem_n19624, MEM_stage_inst_dmem_n19623, MEM_stage_inst_dmem_n19622, MEM_stage_inst_dmem_n19621, MEM_stage_inst_dmem_n19620, MEM_stage_inst_dmem_n19619, MEM_stage_inst_dmem_n19618, MEM_stage_inst_dmem_n19617, MEM_stage_inst_dmem_n19616, MEM_stage_inst_dmem_n19615, MEM_stage_inst_dmem_n19614, MEM_stage_inst_dmem_n19613, MEM_stage_inst_dmem_n19612, MEM_stage_inst_dmem_n19611, MEM_stage_inst_dmem_n19610, MEM_stage_inst_dmem_n19609, MEM_stage_inst_dmem_n19608, MEM_stage_inst_dmem_n19607, MEM_stage_inst_dmem_n19606, MEM_stage_inst_dmem_n19605, MEM_stage_inst_dmem_n19604, MEM_stage_inst_dmem_n19603, MEM_stage_inst_dmem_n19602, MEM_stage_inst_dmem_n19601, MEM_stage_inst_dmem_n19600, MEM_stage_inst_dmem_n19599, MEM_stage_inst_dmem_n19598, MEM_stage_inst_dmem_n19597, MEM_stage_inst_dmem_n19596, MEM_stage_inst_dmem_n19595, MEM_stage_inst_dmem_n19594, MEM_stage_inst_dmem_n19593, MEM_stage_inst_dmem_n19592, MEM_stage_inst_dmem_n19591, MEM_stage_inst_dmem_n19590, MEM_stage_inst_dmem_n19589, MEM_stage_inst_dmem_n19588, MEM_stage_inst_dmem_n19587, MEM_stage_inst_dmem_n19586, MEM_stage_inst_dmem_n19585, MEM_stage_inst_dmem_n19584, MEM_stage_inst_dmem_n19583, MEM_stage_inst_dmem_n19582, MEM_stage_inst_dmem_n19581, MEM_stage_inst_dmem_n19580, MEM_stage_inst_dmem_n19579, MEM_stage_inst_dmem_n19578, MEM_stage_inst_dmem_n19577, MEM_stage_inst_dmem_n19576, MEM_stage_inst_dmem_n19575, MEM_stage_inst_dmem_n19574, MEM_stage_inst_dmem_n19573, MEM_stage_inst_dmem_n19572, MEM_stage_inst_dmem_n19571, MEM_stage_inst_dmem_n19570, MEM_stage_inst_dmem_n19569, MEM_stage_inst_dmem_n19568, MEM_stage_inst_dmem_n19567, MEM_stage_inst_dmem_n19566, MEM_stage_inst_dmem_n19565, MEM_stage_inst_dmem_n19564, MEM_stage_inst_dmem_n19563, MEM_stage_inst_dmem_n19562, MEM_stage_inst_dmem_n19561, MEM_stage_inst_dmem_n19560, MEM_stage_inst_dmem_n19559, MEM_stage_inst_dmem_n19558, MEM_stage_inst_dmem_n19557, MEM_stage_inst_dmem_n19556, MEM_stage_inst_dmem_n19555, MEM_stage_inst_dmem_n19554, MEM_stage_inst_dmem_n19553, MEM_stage_inst_dmem_n19552, MEM_stage_inst_dmem_n19551, MEM_stage_inst_dmem_n19550, MEM_stage_inst_dmem_n19549, MEM_stage_inst_dmem_n19548, MEM_stage_inst_dmem_n19547, MEM_stage_inst_dmem_n19546, MEM_stage_inst_dmem_n19545, MEM_stage_inst_dmem_n19544, MEM_stage_inst_dmem_n19543, MEM_stage_inst_dmem_n19542, MEM_stage_inst_dmem_n19541, MEM_stage_inst_dmem_n19540, MEM_stage_inst_dmem_n19539, MEM_stage_inst_dmem_n19538, MEM_stage_inst_dmem_n19537, MEM_stage_inst_dmem_n19536, MEM_stage_inst_dmem_n19535, MEM_stage_inst_dmem_n19534, MEM_stage_inst_dmem_n19533, MEM_stage_inst_dmem_n19532, MEM_stage_inst_dmem_n19531, MEM_stage_inst_dmem_n19530, MEM_stage_inst_dmem_n19529, MEM_stage_inst_dmem_n19528, MEM_stage_inst_dmem_n19527, MEM_stage_inst_dmem_n19526, MEM_stage_inst_dmem_n19525, MEM_stage_inst_dmem_n19524, MEM_stage_inst_dmem_n19523, MEM_stage_inst_dmem_n19522, MEM_stage_inst_dmem_n19521, MEM_stage_inst_dmem_n19520, MEM_stage_inst_dmem_n19519, MEM_stage_inst_dmem_n19518, MEM_stage_inst_dmem_n19517, MEM_stage_inst_dmem_n19516, MEM_stage_inst_dmem_n19515, MEM_stage_inst_dmem_n19514, MEM_stage_inst_dmem_n19513, MEM_stage_inst_dmem_n19512, MEM_stage_inst_dmem_n19511, MEM_stage_inst_dmem_n19510, MEM_stage_inst_dmem_n19509, MEM_stage_inst_dmem_n19508, MEM_stage_inst_dmem_n19507, MEM_stage_inst_dmem_n19506, MEM_stage_inst_dmem_n19505, MEM_stage_inst_dmem_n19504, MEM_stage_inst_dmem_n19503, MEM_stage_inst_dmem_n19502, MEM_stage_inst_dmem_n19501, MEM_stage_inst_dmem_n19500, MEM_stage_inst_dmem_n19499, MEM_stage_inst_dmem_n19498, MEM_stage_inst_dmem_n19497, MEM_stage_inst_dmem_n19496, MEM_stage_inst_dmem_n19495, MEM_stage_inst_dmem_n19494, MEM_stage_inst_dmem_n19493, MEM_stage_inst_dmem_n19492, MEM_stage_inst_dmem_n19491, MEM_stage_inst_dmem_n19490, MEM_stage_inst_dmem_n19489, MEM_stage_inst_dmem_n19488, MEM_stage_inst_dmem_n19487, MEM_stage_inst_dmem_n19486, MEM_stage_inst_dmem_n19485, MEM_stage_inst_dmem_n19484, MEM_stage_inst_dmem_n19483, MEM_stage_inst_dmem_n19482, MEM_stage_inst_dmem_n19481, MEM_stage_inst_dmem_n19480, MEM_stage_inst_dmem_n19479, MEM_stage_inst_dmem_n19478, MEM_stage_inst_dmem_n19477, MEM_stage_inst_dmem_n19476, MEM_stage_inst_dmem_n19475, MEM_stage_inst_dmem_n19474, MEM_stage_inst_dmem_n19473, MEM_stage_inst_dmem_n19472, MEM_stage_inst_dmem_n19471, MEM_stage_inst_dmem_n19470, MEM_stage_inst_dmem_n19469, MEM_stage_inst_dmem_n19468, MEM_stage_inst_dmem_n19467, MEM_stage_inst_dmem_n19466, MEM_stage_inst_dmem_n19465, MEM_stage_inst_dmem_n19464, MEM_stage_inst_dmem_n19463, MEM_stage_inst_dmem_n19462, MEM_stage_inst_dmem_n19461, MEM_stage_inst_dmem_n19460, MEM_stage_inst_dmem_n19459, MEM_stage_inst_dmem_n19458, MEM_stage_inst_dmem_n19457, MEM_stage_inst_dmem_n19456, MEM_stage_inst_dmem_n19455, MEM_stage_inst_dmem_n19454, MEM_stage_inst_dmem_n19453, MEM_stage_inst_dmem_n19452, MEM_stage_inst_dmem_n19451, MEM_stage_inst_dmem_n19450, MEM_stage_inst_dmem_n19449, MEM_stage_inst_dmem_n19448, MEM_stage_inst_dmem_n19447, MEM_stage_inst_dmem_n19446, MEM_stage_inst_dmem_n19445, MEM_stage_inst_dmem_n19444, MEM_stage_inst_dmem_n19443, MEM_stage_inst_dmem_n19442, MEM_stage_inst_dmem_n19441, MEM_stage_inst_dmem_n19440, MEM_stage_inst_dmem_n19439, MEM_stage_inst_dmem_n19438, MEM_stage_inst_dmem_n19437, MEM_stage_inst_dmem_n19436, MEM_stage_inst_dmem_n19435, MEM_stage_inst_dmem_n19434, MEM_stage_inst_dmem_n19433, MEM_stage_inst_dmem_n19432, MEM_stage_inst_dmem_n19431, MEM_stage_inst_dmem_n19430, MEM_stage_inst_dmem_n19429, MEM_stage_inst_dmem_n19428, MEM_stage_inst_dmem_n19427, MEM_stage_inst_dmem_n19426, MEM_stage_inst_dmem_n19425, MEM_stage_inst_dmem_n19424, MEM_stage_inst_dmem_n19423, MEM_stage_inst_dmem_n19422, MEM_stage_inst_dmem_n19421, MEM_stage_inst_dmem_n19420, MEM_stage_inst_dmem_n19419, MEM_stage_inst_dmem_n19418, MEM_stage_inst_dmem_n19417, MEM_stage_inst_dmem_n19416, MEM_stage_inst_dmem_n19415, MEM_stage_inst_dmem_n19414, MEM_stage_inst_dmem_n19413, MEM_stage_inst_dmem_n19412, MEM_stage_inst_dmem_n19411, MEM_stage_inst_dmem_n19410, MEM_stage_inst_dmem_n19409, MEM_stage_inst_dmem_n19408, MEM_stage_inst_dmem_n19407, MEM_stage_inst_dmem_n19406, MEM_stage_inst_dmem_n19405, MEM_stage_inst_dmem_n19404, MEM_stage_inst_dmem_n19403, MEM_stage_inst_dmem_n19402, MEM_stage_inst_dmem_n19401, MEM_stage_inst_dmem_n19400, MEM_stage_inst_dmem_n19399, MEM_stage_inst_dmem_n19398, MEM_stage_inst_dmem_n19397, MEM_stage_inst_dmem_n19396, MEM_stage_inst_dmem_n19395, MEM_stage_inst_dmem_n19394, MEM_stage_inst_dmem_n19393, MEM_stage_inst_dmem_n19392, MEM_stage_inst_dmem_n19391, MEM_stage_inst_dmem_n19390, MEM_stage_inst_dmem_n19389, MEM_stage_inst_dmem_n19388, MEM_stage_inst_dmem_n19387, MEM_stage_inst_dmem_n19386, MEM_stage_inst_dmem_n19385, MEM_stage_inst_dmem_n19384, MEM_stage_inst_dmem_n19383, MEM_stage_inst_dmem_n19382, MEM_stage_inst_dmem_n19381, MEM_stage_inst_dmem_n19380, MEM_stage_inst_dmem_n19379, MEM_stage_inst_dmem_n19378, MEM_stage_inst_dmem_n19377, MEM_stage_inst_dmem_n19376, MEM_stage_inst_dmem_n19375, MEM_stage_inst_dmem_n19374, MEM_stage_inst_dmem_n19373, MEM_stage_inst_dmem_n19372, MEM_stage_inst_dmem_n19371, MEM_stage_inst_dmem_n19370, MEM_stage_inst_dmem_n19369, MEM_stage_inst_dmem_n19368, MEM_stage_inst_dmem_n19367, MEM_stage_inst_dmem_n19366, MEM_stage_inst_dmem_n19365, MEM_stage_inst_dmem_n19364, MEM_stage_inst_dmem_n19363, MEM_stage_inst_dmem_n19362, MEM_stage_inst_dmem_n19361, MEM_stage_inst_dmem_n19360, MEM_stage_inst_dmem_n19359, MEM_stage_inst_dmem_n19358, MEM_stage_inst_dmem_n19357, MEM_stage_inst_dmem_n19356, MEM_stage_inst_dmem_n19355, MEM_stage_inst_dmem_n19354, MEM_stage_inst_dmem_n19353, MEM_stage_inst_dmem_n19352, MEM_stage_inst_dmem_n19351, MEM_stage_inst_dmem_n19350, MEM_stage_inst_dmem_n19349, MEM_stage_inst_dmem_n19348, MEM_stage_inst_dmem_n19347, MEM_stage_inst_dmem_n19346, MEM_stage_inst_dmem_n19345, MEM_stage_inst_dmem_n19344, MEM_stage_inst_dmem_n19343, MEM_stage_inst_dmem_n19342, MEM_stage_inst_dmem_n19341, MEM_stage_inst_dmem_n19340, MEM_stage_inst_dmem_n19339, MEM_stage_inst_dmem_n19338, MEM_stage_inst_dmem_n19337, MEM_stage_inst_dmem_n19336, MEM_stage_inst_dmem_n19335, MEM_stage_inst_dmem_n19334, MEM_stage_inst_dmem_n19333, MEM_stage_inst_dmem_n19332, MEM_stage_inst_dmem_n19331, MEM_stage_inst_dmem_n19330, MEM_stage_inst_dmem_n19329, MEM_stage_inst_dmem_n19328, MEM_stage_inst_dmem_n19327, MEM_stage_inst_dmem_n19326, MEM_stage_inst_dmem_n19325, MEM_stage_inst_dmem_n19324, MEM_stage_inst_dmem_n19323, MEM_stage_inst_dmem_n19322, MEM_stage_inst_dmem_n19321, MEM_stage_inst_dmem_n19320, MEM_stage_inst_dmem_n19319, MEM_stage_inst_dmem_n19318, MEM_stage_inst_dmem_n19317, MEM_stage_inst_dmem_n19316, MEM_stage_inst_dmem_n19315, MEM_stage_inst_dmem_n19314, MEM_stage_inst_dmem_n19313, MEM_stage_inst_dmem_n19312, MEM_stage_inst_dmem_n19311, MEM_stage_inst_dmem_n19310, MEM_stage_inst_dmem_n19309, MEM_stage_inst_dmem_n19308, MEM_stage_inst_dmem_n19307, MEM_stage_inst_dmem_n19306, MEM_stage_inst_dmem_n19305, MEM_stage_inst_dmem_n19304, MEM_stage_inst_dmem_n19303, MEM_stage_inst_dmem_n19302, MEM_stage_inst_dmem_n19301, MEM_stage_inst_dmem_n19300, MEM_stage_inst_dmem_n19299, MEM_stage_inst_dmem_n19298, MEM_stage_inst_dmem_n19297, MEM_stage_inst_dmem_n19296, MEM_stage_inst_dmem_n19295, MEM_stage_inst_dmem_n19294, MEM_stage_inst_dmem_n19293, MEM_stage_inst_dmem_n19292, MEM_stage_inst_dmem_n19291, MEM_stage_inst_dmem_n19290, MEM_stage_inst_dmem_n19289, MEM_stage_inst_dmem_n19288, MEM_stage_inst_dmem_n19287, MEM_stage_inst_dmem_n19286, MEM_stage_inst_dmem_n19285, MEM_stage_inst_dmem_n19284, MEM_stage_inst_dmem_n19283, MEM_stage_inst_dmem_n19282, MEM_stage_inst_dmem_n19281, MEM_stage_inst_dmem_n19280, MEM_stage_inst_dmem_n19279, MEM_stage_inst_dmem_n19278, MEM_stage_inst_dmem_n19277, MEM_stage_inst_dmem_n19276, MEM_stage_inst_dmem_n19275, MEM_stage_inst_dmem_n19274, MEM_stage_inst_dmem_n19273, MEM_stage_inst_dmem_n19272, MEM_stage_inst_dmem_n19271, MEM_stage_inst_dmem_n19270, MEM_stage_inst_dmem_n19269, MEM_stage_inst_dmem_n19268, MEM_stage_inst_dmem_n19267, MEM_stage_inst_dmem_n19266, MEM_stage_inst_dmem_n19265, MEM_stage_inst_dmem_n19264, MEM_stage_inst_dmem_n19262, MEM_stage_inst_dmem_n19261, MEM_stage_inst_dmem_n19260, MEM_stage_inst_dmem_n19259, MEM_stage_inst_dmem_n19258, MEM_stage_inst_dmem_n19257, MEM_stage_inst_dmem_n19256, MEM_stage_inst_dmem_n19255, MEM_stage_inst_dmem_n19254, MEM_stage_inst_dmem_n19253, MEM_stage_inst_dmem_n19252, MEM_stage_inst_dmem_n19251, MEM_stage_inst_dmem_n19250, MEM_stage_inst_dmem_n19249, MEM_stage_inst_dmem_n19248, MEM_stage_inst_dmem_n19247, MEM_stage_inst_dmem_n19246, MEM_stage_inst_dmem_n19245, MEM_stage_inst_dmem_n19244, MEM_stage_inst_dmem_n19243, MEM_stage_inst_dmem_n19242, MEM_stage_inst_dmem_n19241, MEM_stage_inst_dmem_n19240, MEM_stage_inst_dmem_n19238, MEM_stage_inst_dmem_n19237, MEM_stage_inst_dmem_n19236, MEM_stage_inst_dmem_n19235, MEM_stage_inst_dmem_n19234, MEM_stage_inst_dmem_n19233, MEM_stage_inst_dmem_n19232, MEM_stage_inst_dmem_n19231, MEM_stage_inst_dmem_n19230, MEM_stage_inst_dmem_n19229, MEM_stage_inst_dmem_n19228, MEM_stage_inst_dmem_n19227, MEM_stage_inst_dmem_n19226, MEM_stage_inst_dmem_n19225, MEM_stage_inst_dmem_n19224, MEM_stage_inst_dmem_n19223, MEM_stage_inst_dmem_n19222, MEM_stage_inst_dmem_n19221, MEM_stage_inst_dmem_n19220, MEM_stage_inst_dmem_n19219, MEM_stage_inst_dmem_n19218, MEM_stage_inst_dmem_n19217, MEM_stage_inst_dmem_n19216, MEM_stage_inst_dmem_n19215, MEM_stage_inst_dmem_n19214, MEM_stage_inst_dmem_n19213, MEM_stage_inst_dmem_n19212, MEM_stage_inst_dmem_n19211, MEM_stage_inst_dmem_n19210, MEM_stage_inst_dmem_n19209, MEM_stage_inst_dmem_n19208, MEM_stage_inst_dmem_n19207, MEM_stage_inst_dmem_n19206, MEM_stage_inst_dmem_n19205, MEM_stage_inst_dmem_n19204, MEM_stage_inst_dmem_n19203, MEM_stage_inst_dmem_n19202, MEM_stage_inst_dmem_n19201, MEM_stage_inst_dmem_n19200, MEM_stage_inst_dmem_n19199, MEM_stage_inst_dmem_n19198, MEM_stage_inst_dmem_n19197, MEM_stage_inst_dmem_n19196, MEM_stage_inst_dmem_n19195, MEM_stage_inst_dmem_n19194, MEM_stage_inst_dmem_n19193, MEM_stage_inst_dmem_n19192, MEM_stage_inst_dmem_n19191, MEM_stage_inst_dmem_n19190, MEM_stage_inst_dmem_n19189, MEM_stage_inst_dmem_n19188, MEM_stage_inst_dmem_n19187, MEM_stage_inst_dmem_n19186, MEM_stage_inst_dmem_n19185, MEM_stage_inst_dmem_n19184, MEM_stage_inst_dmem_n19183, MEM_stage_inst_dmem_n19182, MEM_stage_inst_dmem_n19181, MEM_stage_inst_dmem_n19180, MEM_stage_inst_dmem_n19179, MEM_stage_inst_dmem_n19178, MEM_stage_inst_dmem_n19177, MEM_stage_inst_dmem_n19176, MEM_stage_inst_dmem_n19175, MEM_stage_inst_dmem_n19174, MEM_stage_inst_dmem_n19173, MEM_stage_inst_dmem_n19172, MEM_stage_inst_dmem_n19171, MEM_stage_inst_dmem_n19170, MEM_stage_inst_dmem_n19169, MEM_stage_inst_dmem_n19168, MEM_stage_inst_dmem_n19167, MEM_stage_inst_dmem_n19166, MEM_stage_inst_dmem_n19165, MEM_stage_inst_dmem_n19164, MEM_stage_inst_dmem_n19163, MEM_stage_inst_dmem_n19162, MEM_stage_inst_dmem_n19161, MEM_stage_inst_dmem_n19160, MEM_stage_inst_dmem_n19159, MEM_stage_inst_dmem_n19158, MEM_stage_inst_dmem_n19157, MEM_stage_inst_dmem_n19156, MEM_stage_inst_dmem_n19155, MEM_stage_inst_dmem_n19154, MEM_stage_inst_dmem_n19153, MEM_stage_inst_dmem_n19152, MEM_stage_inst_dmem_n19151, MEM_stage_inst_dmem_n19150, MEM_stage_inst_dmem_n19149, MEM_stage_inst_dmem_n19148, MEM_stage_inst_dmem_n19147, MEM_stage_inst_dmem_n19146, MEM_stage_inst_dmem_n19145, MEM_stage_inst_dmem_n19144, MEM_stage_inst_dmem_n19143, MEM_stage_inst_dmem_n19142, MEM_stage_inst_dmem_n19141, MEM_stage_inst_dmem_n19140, MEM_stage_inst_dmem_n19139, MEM_stage_inst_dmem_n19138, MEM_stage_inst_dmem_n19137, MEM_stage_inst_dmem_n19136, MEM_stage_inst_dmem_n19135, MEM_stage_inst_dmem_n19134, MEM_stage_inst_dmem_n19133, MEM_stage_inst_dmem_n19132, MEM_stage_inst_dmem_n19131, MEM_stage_inst_dmem_n19130, MEM_stage_inst_dmem_n19129, MEM_stage_inst_dmem_n19128, MEM_stage_inst_dmem_n19127, MEM_stage_inst_dmem_n19126, MEM_stage_inst_dmem_n19125, MEM_stage_inst_dmem_n19124, MEM_stage_inst_dmem_n19123, MEM_stage_inst_dmem_n19122, MEM_stage_inst_dmem_n19121, MEM_stage_inst_dmem_n19120, MEM_stage_inst_dmem_n19119, MEM_stage_inst_dmem_n19118, MEM_stage_inst_dmem_n19117, MEM_stage_inst_dmem_n19116, MEM_stage_inst_dmem_n19115, MEM_stage_inst_dmem_n19114, MEM_stage_inst_dmem_n19113, MEM_stage_inst_dmem_n19112, MEM_stage_inst_dmem_n19111, MEM_stage_inst_dmem_n19110, MEM_stage_inst_dmem_n19109, MEM_stage_inst_dmem_n19108, MEM_stage_inst_dmem_n19107, MEM_stage_inst_dmem_n19106, MEM_stage_inst_dmem_n19105, MEM_stage_inst_dmem_n19104, MEM_stage_inst_dmem_n19103, MEM_stage_inst_dmem_n19102, MEM_stage_inst_dmem_n19101, MEM_stage_inst_dmem_n19100, MEM_stage_inst_dmem_n19099, MEM_stage_inst_dmem_n19098, MEM_stage_inst_dmem_n19097, MEM_stage_inst_dmem_n19096, MEM_stage_inst_dmem_n19095, MEM_stage_inst_dmem_n19094, MEM_stage_inst_dmem_n19093, MEM_stage_inst_dmem_n19092, MEM_stage_inst_dmem_n19091, MEM_stage_inst_dmem_n19090, MEM_stage_inst_dmem_n19089, MEM_stage_inst_dmem_n19088, MEM_stage_inst_dmem_n19087, MEM_stage_inst_dmem_n19086, MEM_stage_inst_dmem_n19085, MEM_stage_inst_dmem_n19084, MEM_stage_inst_dmem_n19083, MEM_stage_inst_dmem_n19082, MEM_stage_inst_dmem_n19081, MEM_stage_inst_dmem_n19080, MEM_stage_inst_dmem_n19079, MEM_stage_inst_dmem_n19078, MEM_stage_inst_dmem_n19077, MEM_stage_inst_dmem_n19076, MEM_stage_inst_dmem_n19075, MEM_stage_inst_dmem_n19074, MEM_stage_inst_dmem_n19073, MEM_stage_inst_dmem_n19072, MEM_stage_inst_dmem_n19071, MEM_stage_inst_dmem_n19070, MEM_stage_inst_dmem_n19069, MEM_stage_inst_dmem_n19068, MEM_stage_inst_dmem_n19067, MEM_stage_inst_dmem_n19066, MEM_stage_inst_dmem_n19065, MEM_stage_inst_dmem_n19064, MEM_stage_inst_dmem_n19063, MEM_stage_inst_dmem_n19062, MEM_stage_inst_dmem_n19061, MEM_stage_inst_dmem_n19060, MEM_stage_inst_dmem_n19059, MEM_stage_inst_dmem_n19058, MEM_stage_inst_dmem_n19057, MEM_stage_inst_dmem_n19056, MEM_stage_inst_dmem_n19055, MEM_stage_inst_dmem_n19054, MEM_stage_inst_dmem_n19053, MEM_stage_inst_dmem_n19052, MEM_stage_inst_dmem_n19051, MEM_stage_inst_dmem_n19050, MEM_stage_inst_dmem_n19049, MEM_stage_inst_dmem_n19048, MEM_stage_inst_dmem_n19047, MEM_stage_inst_dmem_n19046, MEM_stage_inst_dmem_n19045, MEM_stage_inst_dmem_n19044, MEM_stage_inst_dmem_n19043, MEM_stage_inst_dmem_n19042, MEM_stage_inst_dmem_n19041, MEM_stage_inst_dmem_n19040, MEM_stage_inst_dmem_n19039, MEM_stage_inst_dmem_n19038, MEM_stage_inst_dmem_n19037, MEM_stage_inst_dmem_n19036, MEM_stage_inst_dmem_n19035, MEM_stage_inst_dmem_n19034, MEM_stage_inst_dmem_n19033, MEM_stage_inst_dmem_n19032, MEM_stage_inst_dmem_n19031, MEM_stage_inst_dmem_n19030, MEM_stage_inst_dmem_n19029, MEM_stage_inst_dmem_n19028, MEM_stage_inst_dmem_n19027, MEM_stage_inst_dmem_n19026, MEM_stage_inst_dmem_n19025, MEM_stage_inst_dmem_n19024, MEM_stage_inst_dmem_n19023, MEM_stage_inst_dmem_n19022, MEM_stage_inst_dmem_n19021, MEM_stage_inst_dmem_n19020, MEM_stage_inst_dmem_n19019, MEM_stage_inst_dmem_n19018, MEM_stage_inst_dmem_n19017, MEM_stage_inst_dmem_n19016, MEM_stage_inst_dmem_n19015, MEM_stage_inst_dmem_n19014, MEM_stage_inst_dmem_n19013, MEM_stage_inst_dmem_n19012, MEM_stage_inst_dmem_n19011, MEM_stage_inst_dmem_n19010, MEM_stage_inst_dmem_n19009, MEM_stage_inst_dmem_n19008, MEM_stage_inst_dmem_n19007, MEM_stage_inst_dmem_n19006, MEM_stage_inst_dmem_n19005, MEM_stage_inst_dmem_n19004, MEM_stage_inst_dmem_n19003, MEM_stage_inst_dmem_n19002, MEM_stage_inst_dmem_n19001, MEM_stage_inst_dmem_n19000, MEM_stage_inst_dmem_n18999, MEM_stage_inst_dmem_n18998, MEM_stage_inst_dmem_n18997, MEM_stage_inst_dmem_n18996, MEM_stage_inst_dmem_n18995, MEM_stage_inst_dmem_n18994, MEM_stage_inst_dmem_n18993, MEM_stage_inst_dmem_n18992, MEM_stage_inst_dmem_n18991, MEM_stage_inst_dmem_n18990, MEM_stage_inst_dmem_n18989, MEM_stage_inst_dmem_n18988, MEM_stage_inst_dmem_n18987, MEM_stage_inst_dmem_n18986, MEM_stage_inst_dmem_n18985, MEM_stage_inst_dmem_n18984, MEM_stage_inst_dmem_n18983, MEM_stage_inst_dmem_n18982, MEM_stage_inst_dmem_n18981, MEM_stage_inst_dmem_n18980, MEM_stage_inst_dmem_n18979, MEM_stage_inst_dmem_n18978, MEM_stage_inst_dmem_n18977, MEM_stage_inst_dmem_n18976, MEM_stage_inst_dmem_n18975, MEM_stage_inst_dmem_n18974, MEM_stage_inst_dmem_n18973, MEM_stage_inst_dmem_n18972, MEM_stage_inst_dmem_n18971, MEM_stage_inst_dmem_n18970, MEM_stage_inst_dmem_n18969, MEM_stage_inst_dmem_n18968, MEM_stage_inst_dmem_n18967, MEM_stage_inst_dmem_n18966, MEM_stage_inst_dmem_n18965, MEM_stage_inst_dmem_n18964, MEM_stage_inst_dmem_n18963, MEM_stage_inst_dmem_n18962, MEM_stage_inst_dmem_n18961, MEM_stage_inst_dmem_n18960, MEM_stage_inst_dmem_n18959, MEM_stage_inst_dmem_n18958, MEM_stage_inst_dmem_n18957, MEM_stage_inst_dmem_n18956, MEM_stage_inst_dmem_n18955, MEM_stage_inst_dmem_n18954, MEM_stage_inst_dmem_n18953, MEM_stage_inst_dmem_n18952, MEM_stage_inst_dmem_n18951, MEM_stage_inst_dmem_n18950, MEM_stage_inst_dmem_n18949, MEM_stage_inst_dmem_n18948, MEM_stage_inst_dmem_n18947, MEM_stage_inst_dmem_n18946, MEM_stage_inst_dmem_n18945, MEM_stage_inst_dmem_n18944, MEM_stage_inst_dmem_n18943, MEM_stage_inst_dmem_n18942, MEM_stage_inst_dmem_n18941, MEM_stage_inst_dmem_n18940, MEM_stage_inst_dmem_n18939, MEM_stage_inst_dmem_n18938, MEM_stage_inst_dmem_n18937, MEM_stage_inst_dmem_n18936, MEM_stage_inst_dmem_n18935, MEM_stage_inst_dmem_n18934, MEM_stage_inst_dmem_n18933, MEM_stage_inst_dmem_n18932, MEM_stage_inst_dmem_n18931, MEM_stage_inst_dmem_n18930, MEM_stage_inst_dmem_n18929, MEM_stage_inst_dmem_n18928, MEM_stage_inst_dmem_n18927, MEM_stage_inst_dmem_n18926, MEM_stage_inst_dmem_n18925, MEM_stage_inst_dmem_n18924, MEM_stage_inst_dmem_n18923, MEM_stage_inst_dmem_n18922, MEM_stage_inst_dmem_n18921, MEM_stage_inst_dmem_n18920, MEM_stage_inst_dmem_n18919, MEM_stage_inst_dmem_n18918, MEM_stage_inst_dmem_n18917, MEM_stage_inst_dmem_n18916, MEM_stage_inst_dmem_n18915, MEM_stage_inst_dmem_n18914, MEM_stage_inst_dmem_n18913, MEM_stage_inst_dmem_n18912, MEM_stage_inst_dmem_n18911, MEM_stage_inst_dmem_n18910, MEM_stage_inst_dmem_n18909, MEM_stage_inst_dmem_n18908, MEM_stage_inst_dmem_n18907, MEM_stage_inst_dmem_n18906, MEM_stage_inst_dmem_n18905, MEM_stage_inst_dmem_n18904, MEM_stage_inst_dmem_n18903, MEM_stage_inst_dmem_n18902, MEM_stage_inst_dmem_n18901, MEM_stage_inst_dmem_n18900, MEM_stage_inst_dmem_n18899, MEM_stage_inst_dmem_n18898, MEM_stage_inst_dmem_n18897, MEM_stage_inst_dmem_n18896, MEM_stage_inst_dmem_n18895, MEM_stage_inst_dmem_n18894, MEM_stage_inst_dmem_n18893, MEM_stage_inst_dmem_n18892, MEM_stage_inst_dmem_n18891, MEM_stage_inst_dmem_n18890, MEM_stage_inst_dmem_n18889, MEM_stage_inst_dmem_n18888, MEM_stage_inst_dmem_n18887, MEM_stage_inst_dmem_n18886, MEM_stage_inst_dmem_n18885, MEM_stage_inst_dmem_n18884, MEM_stage_inst_dmem_n18883, MEM_stage_inst_dmem_n18882, MEM_stage_inst_dmem_n18881, MEM_stage_inst_dmem_n18880, MEM_stage_inst_dmem_n18879, MEM_stage_inst_dmem_n18878, MEM_stage_inst_dmem_n18877, MEM_stage_inst_dmem_n18876, MEM_stage_inst_dmem_n18875, MEM_stage_inst_dmem_n18874, MEM_stage_inst_dmem_n18873, MEM_stage_inst_dmem_n18871, MEM_stage_inst_dmem_n18870, MEM_stage_inst_dmem_n18869, MEM_stage_inst_dmem_n18868, MEM_stage_inst_dmem_n18867, MEM_stage_inst_dmem_n18866, MEM_stage_inst_dmem_n18865, MEM_stage_inst_dmem_n18864, MEM_stage_inst_dmem_n18863, MEM_stage_inst_dmem_n18862, MEM_stage_inst_dmem_n18861, MEM_stage_inst_dmem_n18860, MEM_stage_inst_dmem_n18859, MEM_stage_inst_dmem_n18858, MEM_stage_inst_dmem_n18857, MEM_stage_inst_dmem_n18856, MEM_stage_inst_dmem_n18855, MEM_stage_inst_dmem_n18854, MEM_stage_inst_dmem_n18853, MEM_stage_inst_dmem_n18852, MEM_stage_inst_dmem_n18851, MEM_stage_inst_dmem_n18850, MEM_stage_inst_dmem_n18849, MEM_stage_inst_dmem_n18848, MEM_stage_inst_dmem_n18847, MEM_stage_inst_dmem_n18846, MEM_stage_inst_dmem_n18845, MEM_stage_inst_dmem_n18844, MEM_stage_inst_dmem_n18843, MEM_stage_inst_dmem_n18842, MEM_stage_inst_dmem_n18841, MEM_stage_inst_dmem_n18840, MEM_stage_inst_dmem_n18839, MEM_stage_inst_dmem_n18838, MEM_stage_inst_dmem_n18837, MEM_stage_inst_dmem_n18836, MEM_stage_inst_dmem_n18835, MEM_stage_inst_dmem_n18834, MEM_stage_inst_dmem_n18833, MEM_stage_inst_dmem_n18832, MEM_stage_inst_dmem_n18831, MEM_stage_inst_dmem_n18830, MEM_stage_inst_dmem_n18829, MEM_stage_inst_dmem_n18828, MEM_stage_inst_dmem_n18827, MEM_stage_inst_dmem_n18826, MEM_stage_inst_dmem_n18825, MEM_stage_inst_dmem_n18824, MEM_stage_inst_dmem_n18823, MEM_stage_inst_dmem_n18822, MEM_stage_inst_dmem_n18821, MEM_stage_inst_dmem_n18820, MEM_stage_inst_dmem_n18819, MEM_stage_inst_dmem_n18818, MEM_stage_inst_dmem_n18817, MEM_stage_inst_dmem_n18816, MEM_stage_inst_dmem_n18815, MEM_stage_inst_dmem_n18814, MEM_stage_inst_dmem_n18813, MEM_stage_inst_dmem_n18812, MEM_stage_inst_dmem_n18811, MEM_stage_inst_dmem_n18810, MEM_stage_inst_dmem_n18809, MEM_stage_inst_dmem_n18808, MEM_stage_inst_dmem_n18807, MEM_stage_inst_dmem_n18806, MEM_stage_inst_dmem_n18805, MEM_stage_inst_dmem_n18804, MEM_stage_inst_dmem_n18803, MEM_stage_inst_dmem_n18802, MEM_stage_inst_dmem_n18801, MEM_stage_inst_dmem_n18800, MEM_stage_inst_dmem_n18799, MEM_stage_inst_dmem_n18798, MEM_stage_inst_dmem_n18797, MEM_stage_inst_dmem_n18796, MEM_stage_inst_dmem_n18795, MEM_stage_inst_dmem_n18794, MEM_stage_inst_dmem_n18793, MEM_stage_inst_dmem_n18792, MEM_stage_inst_dmem_n18791, MEM_stage_inst_dmem_n18790, MEM_stage_inst_dmem_n18789, MEM_stage_inst_dmem_n18788, MEM_stage_inst_dmem_n18787, MEM_stage_inst_dmem_n18786, MEM_stage_inst_dmem_n18785, MEM_stage_inst_dmem_n18784, MEM_stage_inst_dmem_n18783, MEM_stage_inst_dmem_n18782, MEM_stage_inst_dmem_n18781, MEM_stage_inst_dmem_n18780, MEM_stage_inst_dmem_n18779, MEM_stage_inst_dmem_n18778, MEM_stage_inst_dmem_n18777, MEM_stage_inst_dmem_n18776, MEM_stage_inst_dmem_n18775, MEM_stage_inst_dmem_n18774, MEM_stage_inst_dmem_n18773, MEM_stage_inst_dmem_n18772, MEM_stage_inst_dmem_n18771, MEM_stage_inst_dmem_n18770, MEM_stage_inst_dmem_n18769, MEM_stage_inst_dmem_n18768, MEM_stage_inst_dmem_n18767, MEM_stage_inst_dmem_n18766, MEM_stage_inst_dmem_n18765, MEM_stage_inst_dmem_n18764, MEM_stage_inst_dmem_n18763, MEM_stage_inst_dmem_n18762, MEM_stage_inst_dmem_n18761, MEM_stage_inst_dmem_n18760, MEM_stage_inst_dmem_n18759, MEM_stage_inst_dmem_n18758, MEM_stage_inst_dmem_n18757, MEM_stage_inst_dmem_n18756, MEM_stage_inst_dmem_n18755, MEM_stage_inst_dmem_n18754, MEM_stage_inst_dmem_n18753, MEM_stage_inst_dmem_n18752, MEM_stage_inst_dmem_n18751, MEM_stage_inst_dmem_n18750, MEM_stage_inst_dmem_n18749, MEM_stage_inst_dmem_n18748, MEM_stage_inst_dmem_n18747, MEM_stage_inst_dmem_n18746, MEM_stage_inst_dmem_n18745, MEM_stage_inst_dmem_n18744, MEM_stage_inst_dmem_n18743, MEM_stage_inst_dmem_n18742, MEM_stage_inst_dmem_n18741, MEM_stage_inst_dmem_n18740, MEM_stage_inst_dmem_n18739, MEM_stage_inst_dmem_n18738, MEM_stage_inst_dmem_n18737, MEM_stage_inst_dmem_n18736, MEM_stage_inst_dmem_n18735, MEM_stage_inst_dmem_n18734, MEM_stage_inst_dmem_n18733, MEM_stage_inst_dmem_n18732, MEM_stage_inst_dmem_n18731, MEM_stage_inst_dmem_n18730, MEM_stage_inst_dmem_n18729, MEM_stage_inst_dmem_n18728, MEM_stage_inst_dmem_n18727, MEM_stage_inst_dmem_n18726, MEM_stage_inst_dmem_n18725, MEM_stage_inst_dmem_n18724, MEM_stage_inst_dmem_n18723, MEM_stage_inst_dmem_n18722, MEM_stage_inst_dmem_n18721, MEM_stage_inst_dmem_n18720, MEM_stage_inst_dmem_n18719, MEM_stage_inst_dmem_n18718, MEM_stage_inst_dmem_n18717, MEM_stage_inst_dmem_n18716, MEM_stage_inst_dmem_n18715, MEM_stage_inst_dmem_n18714, MEM_stage_inst_dmem_n18713, MEM_stage_inst_dmem_n18712, MEM_stage_inst_dmem_n18711, MEM_stage_inst_dmem_n18710, MEM_stage_inst_dmem_n18709, MEM_stage_inst_dmem_n18708, MEM_stage_inst_dmem_n18707, MEM_stage_inst_dmem_n18706, MEM_stage_inst_dmem_n18705, MEM_stage_inst_dmem_n18704, MEM_stage_inst_dmem_n18703, MEM_stage_inst_dmem_n18702, MEM_stage_inst_dmem_n18701, MEM_stage_inst_dmem_n18700, MEM_stage_inst_dmem_n18699, MEM_stage_inst_dmem_n18698, MEM_stage_inst_dmem_n18697, MEM_stage_inst_dmem_n18696, MEM_stage_inst_dmem_n18695, MEM_stage_inst_dmem_n18694, MEM_stage_inst_dmem_n18693, MEM_stage_inst_dmem_n18692, MEM_stage_inst_dmem_n18691, MEM_stage_inst_dmem_n18690, MEM_stage_inst_dmem_n18689, MEM_stage_inst_dmem_n18688, MEM_stage_inst_dmem_n18687, MEM_stage_inst_dmem_n18686, MEM_stage_inst_dmem_n18685, MEM_stage_inst_dmem_n18684, MEM_stage_inst_dmem_n18683, MEM_stage_inst_dmem_n18682, MEM_stage_inst_dmem_n18681, MEM_stage_inst_dmem_n18680, MEM_stage_inst_dmem_n18679, MEM_stage_inst_dmem_n18678, MEM_stage_inst_dmem_n18677, MEM_stage_inst_dmem_n18676, MEM_stage_inst_dmem_n18675, MEM_stage_inst_dmem_n18674, MEM_stage_inst_dmem_n18673, MEM_stage_inst_dmem_n18672, MEM_stage_inst_dmem_n18671, MEM_stage_inst_dmem_n18670, MEM_stage_inst_dmem_n18669, MEM_stage_inst_dmem_n18668, MEM_stage_inst_dmem_n18667, MEM_stage_inst_dmem_n18666, MEM_stage_inst_dmem_n18665, MEM_stage_inst_dmem_n18664, MEM_stage_inst_dmem_n18663, MEM_stage_inst_dmem_n18662, MEM_stage_inst_dmem_n18661, MEM_stage_inst_dmem_n18660, MEM_stage_inst_dmem_n18659, MEM_stage_inst_dmem_n18658, MEM_stage_inst_dmem_n18657, MEM_stage_inst_dmem_n18656, MEM_stage_inst_dmem_n18655, MEM_stage_inst_dmem_n18654, MEM_stage_inst_dmem_n18653, MEM_stage_inst_dmem_n18652, MEM_stage_inst_dmem_n18651, MEM_stage_inst_dmem_n18650, MEM_stage_inst_dmem_n18649, MEM_stage_inst_dmem_n18648, MEM_stage_inst_dmem_n18647, MEM_stage_inst_dmem_n18646, MEM_stage_inst_dmem_n18645, MEM_stage_inst_dmem_n18644, MEM_stage_inst_dmem_n18643, MEM_stage_inst_dmem_n18642, MEM_stage_inst_dmem_n18641, MEM_stage_inst_dmem_n18640, MEM_stage_inst_dmem_n18639, MEM_stage_inst_dmem_n18638, MEM_stage_inst_dmem_n18637, MEM_stage_inst_dmem_n18636, MEM_stage_inst_dmem_n18635, MEM_stage_inst_dmem_n18634, MEM_stage_inst_dmem_n18633, MEM_stage_inst_dmem_n18632, MEM_stage_inst_dmem_n18631, MEM_stage_inst_dmem_n18630, MEM_stage_inst_dmem_n18629, MEM_stage_inst_dmem_n18628, MEM_stage_inst_dmem_n18627, MEM_stage_inst_dmem_n18626, MEM_stage_inst_dmem_n18625, MEM_stage_inst_dmem_n18624, MEM_stage_inst_dmem_n18623, MEM_stage_inst_dmem_n18622, MEM_stage_inst_dmem_n18621, MEM_stage_inst_dmem_n18620, MEM_stage_inst_dmem_n18619, MEM_stage_inst_dmem_n18618, MEM_stage_inst_dmem_n18617, MEM_stage_inst_dmem_n18616, MEM_stage_inst_dmem_n18615, MEM_stage_inst_dmem_n18614, MEM_stage_inst_dmem_n18613, MEM_stage_inst_dmem_n18612, MEM_stage_inst_dmem_n18611, MEM_stage_inst_dmem_n18610, MEM_stage_inst_dmem_n18609, MEM_stage_inst_dmem_n18608, MEM_stage_inst_dmem_n18607, MEM_stage_inst_dmem_n18606, MEM_stage_inst_dmem_n18605, MEM_stage_inst_dmem_n18604, MEM_stage_inst_dmem_n18603, MEM_stage_inst_dmem_n18602, MEM_stage_inst_dmem_n18601, MEM_stage_inst_dmem_n18600, MEM_stage_inst_dmem_n18599, MEM_stage_inst_dmem_n18598, MEM_stage_inst_dmem_n18597, MEM_stage_inst_dmem_n18596, MEM_stage_inst_dmem_n18595, MEM_stage_inst_dmem_n18594, MEM_stage_inst_dmem_n18593, MEM_stage_inst_dmem_n18592, MEM_stage_inst_dmem_n18591, MEM_stage_inst_dmem_n18590, MEM_stage_inst_dmem_n18589, MEM_stage_inst_dmem_n18588, MEM_stage_inst_dmem_n18587, MEM_stage_inst_dmem_n18586, MEM_stage_inst_dmem_n18585, MEM_stage_inst_dmem_n18584, MEM_stage_inst_dmem_n18583, MEM_stage_inst_dmem_n18582, MEM_stage_inst_dmem_n18581, MEM_stage_inst_dmem_n18580, MEM_stage_inst_dmem_n18579, MEM_stage_inst_dmem_n18578, MEM_stage_inst_dmem_n18577, MEM_stage_inst_dmem_n18576, MEM_stage_inst_dmem_n18575, MEM_stage_inst_dmem_n18574, MEM_stage_inst_dmem_n18573, MEM_stage_inst_dmem_n18572, MEM_stage_inst_dmem_n18571, MEM_stage_inst_dmem_n18570, MEM_stage_inst_dmem_n18569, MEM_stage_inst_dmem_n18568, MEM_stage_inst_dmem_n18567, MEM_stage_inst_dmem_n18566, MEM_stage_inst_dmem_n18565, MEM_stage_inst_dmem_n18564, MEM_stage_inst_dmem_n18563, MEM_stage_inst_dmem_n18562, MEM_stage_inst_dmem_n18561, MEM_stage_inst_dmem_n18560, MEM_stage_inst_dmem_n18559, MEM_stage_inst_dmem_n18558, MEM_stage_inst_dmem_n18557, MEM_stage_inst_dmem_n18556, MEM_stage_inst_dmem_n18555, MEM_stage_inst_dmem_n18554, MEM_stage_inst_dmem_n18553, MEM_stage_inst_dmem_n18552, MEM_stage_inst_dmem_n18551, MEM_stage_inst_dmem_n18550, MEM_stage_inst_dmem_n18549, MEM_stage_inst_dmem_n18548, MEM_stage_inst_dmem_n18547, MEM_stage_inst_dmem_n18546, MEM_stage_inst_dmem_n18545, MEM_stage_inst_dmem_n18544, MEM_stage_inst_dmem_n18543, MEM_stage_inst_dmem_n18542, MEM_stage_inst_dmem_n18541, MEM_stage_inst_dmem_n18540, MEM_stage_inst_dmem_n18539, MEM_stage_inst_dmem_n18538, MEM_stage_inst_dmem_n18537, MEM_stage_inst_dmem_n18536, MEM_stage_inst_dmem_n18535, MEM_stage_inst_dmem_n18534, MEM_stage_inst_dmem_n18533, MEM_stage_inst_dmem_n18532, MEM_stage_inst_dmem_n18531, MEM_stage_inst_dmem_n18530, MEM_stage_inst_dmem_n18529, MEM_stage_inst_dmem_n18528, MEM_stage_inst_dmem_n18527, MEM_stage_inst_dmem_n18526, MEM_stage_inst_dmem_n18525, MEM_stage_inst_dmem_n18524, MEM_stage_inst_dmem_n18523, MEM_stage_inst_dmem_n18522, MEM_stage_inst_dmem_n18521, MEM_stage_inst_dmem_n18520, MEM_stage_inst_dmem_n18519, MEM_stage_inst_dmem_n18518, MEM_stage_inst_dmem_n18517, MEM_stage_inst_dmem_n18516, MEM_stage_inst_dmem_n18515, MEM_stage_inst_dmem_n18514, MEM_stage_inst_dmem_n18513, MEM_stage_inst_dmem_n18512, MEM_stage_inst_dmem_n18511, MEM_stage_inst_dmem_n18510, MEM_stage_inst_dmem_n18509, MEM_stage_inst_dmem_n18508, MEM_stage_inst_dmem_n18507, MEM_stage_inst_dmem_n18506, MEM_stage_inst_dmem_n18505, MEM_stage_inst_dmem_n18504, MEM_stage_inst_dmem_n18503, MEM_stage_inst_dmem_n18502, MEM_stage_inst_dmem_n18501, MEM_stage_inst_dmem_n18500, MEM_stage_inst_dmem_n18499, MEM_stage_inst_dmem_n18498, MEM_stage_inst_dmem_n18497, MEM_stage_inst_dmem_n18496, MEM_stage_inst_dmem_n18495, MEM_stage_inst_dmem_n18494, MEM_stage_inst_dmem_n18493, MEM_stage_inst_dmem_n18492, MEM_stage_inst_dmem_n18491, MEM_stage_inst_dmem_n18490, MEM_stage_inst_dmem_n18489, MEM_stage_inst_dmem_n18488, MEM_stage_inst_dmem_n18487, MEM_stage_inst_dmem_n18486, MEM_stage_inst_dmem_n18485, MEM_stage_inst_dmem_n18484, MEM_stage_inst_dmem_n18483, MEM_stage_inst_dmem_n18482, MEM_stage_inst_dmem_n18481, MEM_stage_inst_dmem_n18480, MEM_stage_inst_dmem_n18479, MEM_stage_inst_dmem_n18478, MEM_stage_inst_dmem_n18477, MEM_stage_inst_dmem_n18476, MEM_stage_inst_dmem_n18475, MEM_stage_inst_dmem_n18474, MEM_stage_inst_dmem_n18473, MEM_stage_inst_dmem_n18472, MEM_stage_inst_dmem_n18471, MEM_stage_inst_dmem_n18470, MEM_stage_inst_dmem_n18469, MEM_stage_inst_dmem_n18468, MEM_stage_inst_dmem_n18467, MEM_stage_inst_dmem_n18466, MEM_stage_inst_dmem_n18465, MEM_stage_inst_dmem_n18464, MEM_stage_inst_dmem_n18463, MEM_stage_inst_dmem_n18462, MEM_stage_inst_dmem_n18461, MEM_stage_inst_dmem_n18460, MEM_stage_inst_dmem_n18459, MEM_stage_inst_dmem_n18458, MEM_stage_inst_dmem_n18457, MEM_stage_inst_dmem_n18456, MEM_stage_inst_dmem_n18455, MEM_stage_inst_dmem_n18454, MEM_stage_inst_dmem_n18453, MEM_stage_inst_dmem_n18452, MEM_stage_inst_dmem_n18451, MEM_stage_inst_dmem_n18450, MEM_stage_inst_dmem_n18449, MEM_stage_inst_dmem_n18448, MEM_stage_inst_dmem_n18447, MEM_stage_inst_dmem_n18446, MEM_stage_inst_dmem_n18445, MEM_stage_inst_dmem_n18444, MEM_stage_inst_dmem_n18443, MEM_stage_inst_dmem_n18442, MEM_stage_inst_dmem_n18441, MEM_stage_inst_dmem_n18440, MEM_stage_inst_dmem_n18439, MEM_stage_inst_dmem_n18438, MEM_stage_inst_dmem_n18437, MEM_stage_inst_dmem_n18436, MEM_stage_inst_dmem_n18435, MEM_stage_inst_dmem_n18434, MEM_stage_inst_dmem_n18433, MEM_stage_inst_dmem_n18432, MEM_stage_inst_dmem_n18431, MEM_stage_inst_dmem_n18430, MEM_stage_inst_dmem_n18429, MEM_stage_inst_dmem_n18428, MEM_stage_inst_dmem_n18427, MEM_stage_inst_dmem_n18426, MEM_stage_inst_dmem_n18425, MEM_stage_inst_dmem_n18424, MEM_stage_inst_dmem_n18423, MEM_stage_inst_dmem_n18422, MEM_stage_inst_dmem_n18421, MEM_stage_inst_dmem_n18420, MEM_stage_inst_dmem_n18419, MEM_stage_inst_dmem_n18418, MEM_stage_inst_dmem_n18417, MEM_stage_inst_dmem_n18416, MEM_stage_inst_dmem_n18415, MEM_stage_inst_dmem_n18414, MEM_stage_inst_dmem_n18413, MEM_stage_inst_dmem_n18412, MEM_stage_inst_dmem_n18411, MEM_stage_inst_dmem_n18410, MEM_stage_inst_dmem_n18409, MEM_stage_inst_dmem_n18408, MEM_stage_inst_dmem_n18407, MEM_stage_inst_dmem_n18406, MEM_stage_inst_dmem_n18405, MEM_stage_inst_dmem_n18404, MEM_stage_inst_dmem_n18403, MEM_stage_inst_dmem_n18402, MEM_stage_inst_dmem_n18401, MEM_stage_inst_dmem_n18400, MEM_stage_inst_dmem_n18399, MEM_stage_inst_dmem_n18398, MEM_stage_inst_dmem_n18397, MEM_stage_inst_dmem_n18396, MEM_stage_inst_dmem_n18395, MEM_stage_inst_dmem_n18394, MEM_stage_inst_dmem_n18393, MEM_stage_inst_dmem_n18392, MEM_stage_inst_dmem_n18391, MEM_stage_inst_dmem_n18390, MEM_stage_inst_dmem_n18389, MEM_stage_inst_dmem_n18388, MEM_stage_inst_dmem_n18387, MEM_stage_inst_dmem_n18386, MEM_stage_inst_dmem_n18385, MEM_stage_inst_dmem_n18384, MEM_stage_inst_dmem_n18383, MEM_stage_inst_dmem_n18382, MEM_stage_inst_dmem_n18381, MEM_stage_inst_dmem_n18380, MEM_stage_inst_dmem_n18379, MEM_stage_inst_dmem_n18378, MEM_stage_inst_dmem_n18377, MEM_stage_inst_dmem_n18376, MEM_stage_inst_dmem_n18375, MEM_stage_inst_dmem_n18374, MEM_stage_inst_dmem_n18373, MEM_stage_inst_dmem_n18372, MEM_stage_inst_dmem_n18371, MEM_stage_inst_dmem_n18370, MEM_stage_inst_dmem_n18369, MEM_stage_inst_dmem_n18368, MEM_stage_inst_dmem_n18367, MEM_stage_inst_dmem_n18366, MEM_stage_inst_dmem_n18365, MEM_stage_inst_dmem_n18364, MEM_stage_inst_dmem_n18363, MEM_stage_inst_dmem_n18362, MEM_stage_inst_dmem_n18361, MEM_stage_inst_dmem_n18360, MEM_stage_inst_dmem_n18359, MEM_stage_inst_dmem_n18358, MEM_stage_inst_dmem_n18357, MEM_stage_inst_dmem_n18356, MEM_stage_inst_dmem_n18355, MEM_stage_inst_dmem_n18354, MEM_stage_inst_dmem_n18353, MEM_stage_inst_dmem_n18352, MEM_stage_inst_dmem_n18351, MEM_stage_inst_dmem_n18350, MEM_stage_inst_dmem_n18349, MEM_stage_inst_dmem_n18348, MEM_stage_inst_dmem_n18347, MEM_stage_inst_dmem_n18346, MEM_stage_inst_dmem_n18345, MEM_stage_inst_dmem_n18344, MEM_stage_inst_dmem_n18343, MEM_stage_inst_dmem_n18342, MEM_stage_inst_dmem_n18341, MEM_stage_inst_dmem_n18340, MEM_stage_inst_dmem_n18339, MEM_stage_inst_dmem_n18338, MEM_stage_inst_dmem_n18337, MEM_stage_inst_dmem_n18336, MEM_stage_inst_dmem_n18335, MEM_stage_inst_dmem_n18334, MEM_stage_inst_dmem_n18333, MEM_stage_inst_dmem_n18332, MEM_stage_inst_dmem_n18331, MEM_stage_inst_dmem_n18330, MEM_stage_inst_dmem_n18329, MEM_stage_inst_dmem_n18328, MEM_stage_inst_dmem_n18327, MEM_stage_inst_dmem_n18326, MEM_stage_inst_dmem_n18325, MEM_stage_inst_dmem_n18324, MEM_stage_inst_dmem_n18323, MEM_stage_inst_dmem_n18322, MEM_stage_inst_dmem_n18321, MEM_stage_inst_dmem_n18320, MEM_stage_inst_dmem_n18319, MEM_stage_inst_dmem_n18318, MEM_stage_inst_dmem_n18317, MEM_stage_inst_dmem_n18316, MEM_stage_inst_dmem_n18315, MEM_stage_inst_dmem_n18314, MEM_stage_inst_dmem_n18313, MEM_stage_inst_dmem_n18312, MEM_stage_inst_dmem_n18311, MEM_stage_inst_dmem_n18310, MEM_stage_inst_dmem_n18309, MEM_stage_inst_dmem_n18308, MEM_stage_inst_dmem_n18307, MEM_stage_inst_dmem_n18306, MEM_stage_inst_dmem_n18305, MEM_stage_inst_dmem_n18304, MEM_stage_inst_dmem_n18303, MEM_stage_inst_dmem_n18302, MEM_stage_inst_dmem_n18301, MEM_stage_inst_dmem_n18300, MEM_stage_inst_dmem_n18299, MEM_stage_inst_dmem_n18298, MEM_stage_inst_dmem_n18297, MEM_stage_inst_dmem_n18296, MEM_stage_inst_dmem_n18295, MEM_stage_inst_dmem_n18294, MEM_stage_inst_dmem_n18293, MEM_stage_inst_dmem_n18292, MEM_stage_inst_dmem_n18291, MEM_stage_inst_dmem_n18290, MEM_stage_inst_dmem_n18289, MEM_stage_inst_dmem_n18288, MEM_stage_inst_dmem_n18287, MEM_stage_inst_dmem_n18286, MEM_stage_inst_dmem_n18285, MEM_stage_inst_dmem_n18284, MEM_stage_inst_dmem_n18283, MEM_stage_inst_dmem_n18282, MEM_stage_inst_dmem_n18281, MEM_stage_inst_dmem_n18280, MEM_stage_inst_dmem_n18279, MEM_stage_inst_dmem_n18278, MEM_stage_inst_dmem_n18277, MEM_stage_inst_dmem_n18276, MEM_stage_inst_dmem_n18275, MEM_stage_inst_dmem_n18274, MEM_stage_inst_dmem_n18273, MEM_stage_inst_dmem_n18272, MEM_stage_inst_dmem_n18271, MEM_stage_inst_dmem_n18270, MEM_stage_inst_dmem_n18269, MEM_stage_inst_dmem_n18268, MEM_stage_inst_dmem_n18267, MEM_stage_inst_dmem_n18266, MEM_stage_inst_dmem_n18265, MEM_stage_inst_dmem_n18264, MEM_stage_inst_dmem_n18263, MEM_stage_inst_dmem_n18262, MEM_stage_inst_dmem_n18261, MEM_stage_inst_dmem_n18260, MEM_stage_inst_dmem_n18259, MEM_stage_inst_dmem_n18258, MEM_stage_inst_dmem_n18257, MEM_stage_inst_dmem_n18256, MEM_stage_inst_dmem_n18255, MEM_stage_inst_dmem_n18254, MEM_stage_inst_dmem_n18253, MEM_stage_inst_dmem_n18252, MEM_stage_inst_dmem_n18251, MEM_stage_inst_dmem_n18250, MEM_stage_inst_dmem_n18249, MEM_stage_inst_dmem_n18248, MEM_stage_inst_dmem_n18247, MEM_stage_inst_dmem_n18246, MEM_stage_inst_dmem_n18245, MEM_stage_inst_dmem_n18244, MEM_stage_inst_dmem_n18243, MEM_stage_inst_dmem_n18242, MEM_stage_inst_dmem_n18241, MEM_stage_inst_dmem_n18240, MEM_stage_inst_dmem_n18239, MEM_stage_inst_dmem_n18238, MEM_stage_inst_dmem_n18237, MEM_stage_inst_dmem_n18236, MEM_stage_inst_dmem_n18235, MEM_stage_inst_dmem_n18234, MEM_stage_inst_dmem_n18233, MEM_stage_inst_dmem_n18232, MEM_stage_inst_dmem_n18231, MEM_stage_inst_dmem_n18230, MEM_stage_inst_dmem_n18229, MEM_stage_inst_dmem_n18228, MEM_stage_inst_dmem_n18227, MEM_stage_inst_dmem_n18226, MEM_stage_inst_dmem_n18225, MEM_stage_inst_dmem_n18224, MEM_stage_inst_dmem_n18223, MEM_stage_inst_dmem_n18222, MEM_stage_inst_dmem_n18221, MEM_stage_inst_dmem_n18220, MEM_stage_inst_dmem_n18219, MEM_stage_inst_dmem_n18218, MEM_stage_inst_dmem_n18217, MEM_stage_inst_dmem_n18216, MEM_stage_inst_dmem_n18215, MEM_stage_inst_dmem_n18214, MEM_stage_inst_dmem_n18213, MEM_stage_inst_dmem_n18212, MEM_stage_inst_dmem_n18211, MEM_stage_inst_dmem_n18210, MEM_stage_inst_dmem_n18209, MEM_stage_inst_dmem_n18208, MEM_stage_inst_dmem_n18207, MEM_stage_inst_dmem_n18206, MEM_stage_inst_dmem_n18205, MEM_stage_inst_dmem_n18204, MEM_stage_inst_dmem_n18203, MEM_stage_inst_dmem_n18202, MEM_stage_inst_dmem_n18201, MEM_stage_inst_dmem_n18200, MEM_stage_inst_dmem_n18199, MEM_stage_inst_dmem_n18198, MEM_stage_inst_dmem_n18197, MEM_stage_inst_dmem_n18196, MEM_stage_inst_dmem_n18195, MEM_stage_inst_dmem_n18194, MEM_stage_inst_dmem_n18193, MEM_stage_inst_dmem_n18192, MEM_stage_inst_dmem_n18191, MEM_stage_inst_dmem_n18190, MEM_stage_inst_dmem_n18189, MEM_stage_inst_dmem_n18188, MEM_stage_inst_dmem_n18187, MEM_stage_inst_dmem_n18186, MEM_stage_inst_dmem_n18185, MEM_stage_inst_dmem_n18184, MEM_stage_inst_dmem_n18183, MEM_stage_inst_dmem_n18182, MEM_stage_inst_dmem_n18181, MEM_stage_inst_dmem_n18180, MEM_stage_inst_dmem_n18179, MEM_stage_inst_dmem_n18178, MEM_stage_inst_dmem_n18177, MEM_stage_inst_dmem_n18176, MEM_stage_inst_dmem_n18175, MEM_stage_inst_dmem_n18174, MEM_stage_inst_dmem_n18173, MEM_stage_inst_dmem_n18172, MEM_stage_inst_dmem_n18171, MEM_stage_inst_dmem_n18170, MEM_stage_inst_dmem_n18169, MEM_stage_inst_dmem_n18168, MEM_stage_inst_dmem_n18167, MEM_stage_inst_dmem_n18166, MEM_stage_inst_dmem_n18165, MEM_stage_inst_dmem_n18164, MEM_stage_inst_dmem_n18163, MEM_stage_inst_dmem_n18162, MEM_stage_inst_dmem_n18161, MEM_stage_inst_dmem_n18160, MEM_stage_inst_dmem_n18159, MEM_stage_inst_dmem_n18158, MEM_stage_inst_dmem_n18157, MEM_stage_inst_dmem_n18156, MEM_stage_inst_dmem_n18155, MEM_stage_inst_dmem_n18154, MEM_stage_inst_dmem_n18153, MEM_stage_inst_dmem_n18152, MEM_stage_inst_dmem_n18151, MEM_stage_inst_dmem_n18150, MEM_stage_inst_dmem_n18149, MEM_stage_inst_dmem_n18148, MEM_stage_inst_dmem_n18147, MEM_stage_inst_dmem_n18146, MEM_stage_inst_dmem_n18145, MEM_stage_inst_dmem_n18144, MEM_stage_inst_dmem_n18143, MEM_stage_inst_dmem_n18142, MEM_stage_inst_dmem_n18141, MEM_stage_inst_dmem_n18140, MEM_stage_inst_dmem_n18139, MEM_stage_inst_dmem_n18138, MEM_stage_inst_dmem_n18137, MEM_stage_inst_dmem_n18136, MEM_stage_inst_dmem_n18135, MEM_stage_inst_dmem_n18134, MEM_stage_inst_dmem_n18133, MEM_stage_inst_dmem_n18132, MEM_stage_inst_dmem_n18131, MEM_stage_inst_dmem_n18130, MEM_stage_inst_dmem_n18129, MEM_stage_inst_dmem_n18128, MEM_stage_inst_dmem_n18127, MEM_stage_inst_dmem_n18126, MEM_stage_inst_dmem_n18125, MEM_stage_inst_dmem_n18124, MEM_stage_inst_dmem_n18123, MEM_stage_inst_dmem_n18122, MEM_stage_inst_dmem_n18121, MEM_stage_inst_dmem_n18120, MEM_stage_inst_dmem_n18119, MEM_stage_inst_dmem_n18118, MEM_stage_inst_dmem_n18117, MEM_stage_inst_dmem_n18116, MEM_stage_inst_dmem_n18115, MEM_stage_inst_dmem_n18114, MEM_stage_inst_dmem_n18113, MEM_stage_inst_dmem_n18112, MEM_stage_inst_dmem_n18111, MEM_stage_inst_dmem_n18110, MEM_stage_inst_dmem_n18109, MEM_stage_inst_dmem_n18108, MEM_stage_inst_dmem_n18107, MEM_stage_inst_dmem_n18106, MEM_stage_inst_dmem_n18105, MEM_stage_inst_dmem_n18104, MEM_stage_inst_dmem_n18103, MEM_stage_inst_dmem_n18102, MEM_stage_inst_dmem_n18101, MEM_stage_inst_dmem_n18100, MEM_stage_inst_dmem_n18099, MEM_stage_inst_dmem_n18098, MEM_stage_inst_dmem_n18097, MEM_stage_inst_dmem_n18096, MEM_stage_inst_dmem_n18095, MEM_stage_inst_dmem_n18094, MEM_stage_inst_dmem_n18093, MEM_stage_inst_dmem_n18092, MEM_stage_inst_dmem_n18091, MEM_stage_inst_dmem_n18090, MEM_stage_inst_dmem_n18089, MEM_stage_inst_dmem_n18088, MEM_stage_inst_dmem_n18087, MEM_stage_inst_dmem_n18086, MEM_stage_inst_dmem_n18085, MEM_stage_inst_dmem_n18084, MEM_stage_inst_dmem_n18083, MEM_stage_inst_dmem_n18082, MEM_stage_inst_dmem_n18081, MEM_stage_inst_dmem_n18080, MEM_stage_inst_dmem_n18079, MEM_stage_inst_dmem_n18078, MEM_stage_inst_dmem_n18077, MEM_stage_inst_dmem_n18076, MEM_stage_inst_dmem_n18075, MEM_stage_inst_dmem_n18074, MEM_stage_inst_dmem_n18073, MEM_stage_inst_dmem_n18072, MEM_stage_inst_dmem_n18071, MEM_stage_inst_dmem_n18070, MEM_stage_inst_dmem_n18069, MEM_stage_inst_dmem_n18068, MEM_stage_inst_dmem_n18067, MEM_stage_inst_dmem_n18066, MEM_stage_inst_dmem_n18065, MEM_stage_inst_dmem_n18064, MEM_stage_inst_dmem_n18063, MEM_stage_inst_dmem_n18062, MEM_stage_inst_dmem_n18061, MEM_stage_inst_dmem_n18060, MEM_stage_inst_dmem_n18059, MEM_stage_inst_dmem_n18058, MEM_stage_inst_dmem_n18057, MEM_stage_inst_dmem_n18056, MEM_stage_inst_dmem_n18055, MEM_stage_inst_dmem_n18054, MEM_stage_inst_dmem_n18053, MEM_stage_inst_dmem_n18052, MEM_stage_inst_dmem_n18051, MEM_stage_inst_dmem_n18050, MEM_stage_inst_dmem_n18049, MEM_stage_inst_dmem_n18048, MEM_stage_inst_dmem_n18047, MEM_stage_inst_dmem_n18046, MEM_stage_inst_dmem_n18045, MEM_stage_inst_dmem_n18044, MEM_stage_inst_dmem_n18043, MEM_stage_inst_dmem_n18042, MEM_stage_inst_dmem_n18041, MEM_stage_inst_dmem_n18040, MEM_stage_inst_dmem_n18039, MEM_stage_inst_dmem_n18038, MEM_stage_inst_dmem_n18037, MEM_stage_inst_dmem_n18036, MEM_stage_inst_dmem_n18035, MEM_stage_inst_dmem_n18034, MEM_stage_inst_dmem_n18033, MEM_stage_inst_dmem_n18032, MEM_stage_inst_dmem_n18031, MEM_stage_inst_dmem_n18030, MEM_stage_inst_dmem_n18029, MEM_stage_inst_dmem_n18028, MEM_stage_inst_dmem_n18027, MEM_stage_inst_dmem_n18026, MEM_stage_inst_dmem_n18025, MEM_stage_inst_dmem_n18024, MEM_stage_inst_dmem_n18023, MEM_stage_inst_dmem_n18022, MEM_stage_inst_dmem_n18021, MEM_stage_inst_dmem_n18020, MEM_stage_inst_dmem_n18019, MEM_stage_inst_dmem_n18018, MEM_stage_inst_dmem_n18017, MEM_stage_inst_dmem_n18016, MEM_stage_inst_dmem_n18015, MEM_stage_inst_dmem_n18014, MEM_stage_inst_dmem_n18013, MEM_stage_inst_dmem_n18012, MEM_stage_inst_dmem_n18011, MEM_stage_inst_dmem_n18009, MEM_stage_inst_dmem_n18008, MEM_stage_inst_dmem_n18007, MEM_stage_inst_dmem_n18006, MEM_stage_inst_dmem_n18005, MEM_stage_inst_dmem_n18004, MEM_stage_inst_dmem_n18003, MEM_stage_inst_dmem_n18002, MEM_stage_inst_dmem_n18001, MEM_stage_inst_dmem_n18000, MEM_stage_inst_dmem_n17999, MEM_stage_inst_dmem_n17998, MEM_stage_inst_dmem_n17997, MEM_stage_inst_dmem_n17996, MEM_stage_inst_dmem_n17995, MEM_stage_inst_dmem_n17994, MEM_stage_inst_dmem_n17993, MEM_stage_inst_dmem_n17992, MEM_stage_inst_dmem_n17991, MEM_stage_inst_dmem_n17990, MEM_stage_inst_dmem_n17989, MEM_stage_inst_dmem_n17988, MEM_stage_inst_dmem_n17987, MEM_stage_inst_dmem_n17986, MEM_stage_inst_dmem_n17985, MEM_stage_inst_dmem_n17984, MEM_stage_inst_dmem_n17983, MEM_stage_inst_dmem_n17982, MEM_stage_inst_dmem_n17981, MEM_stage_inst_dmem_n17980, MEM_stage_inst_dmem_n17979, MEM_stage_inst_dmem_n17978, MEM_stage_inst_dmem_n17977, MEM_stage_inst_dmem_n17976, MEM_stage_inst_dmem_n17975, MEM_stage_inst_dmem_n17974, MEM_stage_inst_dmem_n17973, MEM_stage_inst_dmem_n17972, MEM_stage_inst_dmem_n17971, MEM_stage_inst_dmem_n17970, MEM_stage_inst_dmem_n17969, MEM_stage_inst_dmem_n17968, MEM_stage_inst_dmem_n17967, MEM_stage_inst_dmem_n17966, MEM_stage_inst_dmem_n17965, MEM_stage_inst_dmem_n17964, MEM_stage_inst_dmem_n17963, MEM_stage_inst_dmem_n17962, MEM_stage_inst_dmem_n17961, MEM_stage_inst_dmem_n17960, MEM_stage_inst_dmem_n17959, MEM_stage_inst_dmem_n17958, MEM_stage_inst_dmem_n17957, MEM_stage_inst_dmem_n17956, MEM_stage_inst_dmem_n17955, MEM_stage_inst_dmem_n17954, MEM_stage_inst_dmem_n17953, MEM_stage_inst_dmem_n17952, MEM_stage_inst_dmem_n17951, MEM_stage_inst_dmem_n17950, MEM_stage_inst_dmem_n17949, MEM_stage_inst_dmem_n17948, MEM_stage_inst_dmem_n17947, MEM_stage_inst_dmem_n17946, MEM_stage_inst_dmem_n17945, MEM_stage_inst_dmem_n17944, MEM_stage_inst_dmem_n17943, MEM_stage_inst_dmem_n17942, MEM_stage_inst_dmem_n17941, MEM_stage_inst_dmem_n17940, MEM_stage_inst_dmem_n17939, MEM_stage_inst_dmem_n17938, MEM_stage_inst_dmem_n17937, MEM_stage_inst_dmem_n17936, MEM_stage_inst_dmem_n17935, MEM_stage_inst_dmem_n17934, MEM_stage_inst_dmem_n17933, MEM_stage_inst_dmem_n17932, MEM_stage_inst_dmem_n17931, MEM_stage_inst_dmem_n17930, MEM_stage_inst_dmem_n17929, MEM_stage_inst_dmem_n17928, MEM_stage_inst_dmem_n17927, MEM_stage_inst_dmem_n17926, MEM_stage_inst_dmem_n17925, MEM_stage_inst_dmem_n17924, MEM_stage_inst_dmem_n17923, MEM_stage_inst_dmem_n17922, MEM_stage_inst_dmem_n17921, MEM_stage_inst_dmem_n17920, MEM_stage_inst_dmem_n17919, MEM_stage_inst_dmem_n17918, MEM_stage_inst_dmem_n17917, MEM_stage_inst_dmem_n17916, MEM_stage_inst_dmem_n17915, MEM_stage_inst_dmem_n17914, MEM_stage_inst_dmem_n17913, MEM_stage_inst_dmem_n17912, MEM_stage_inst_dmem_n17911, MEM_stage_inst_dmem_n17910, MEM_stage_inst_dmem_n17909, MEM_stage_inst_dmem_n17908, MEM_stage_inst_dmem_n17907, MEM_stage_inst_dmem_n17906, MEM_stage_inst_dmem_n17905, MEM_stage_inst_dmem_n17904, MEM_stage_inst_dmem_n17903, MEM_stage_inst_dmem_n17902, MEM_stage_inst_dmem_n17901, MEM_stage_inst_dmem_n17900, MEM_stage_inst_dmem_n17899, MEM_stage_inst_dmem_n17898, MEM_stage_inst_dmem_n17897, MEM_stage_inst_dmem_n17896, MEM_stage_inst_dmem_n17895, MEM_stage_inst_dmem_n17894, MEM_stage_inst_dmem_n17893, MEM_stage_inst_dmem_n17892, MEM_stage_inst_dmem_n17891, MEM_stage_inst_dmem_n17890, MEM_stage_inst_dmem_n17889, MEM_stage_inst_dmem_n17888, MEM_stage_inst_dmem_n17887, MEM_stage_inst_dmem_n17886, MEM_stage_inst_dmem_n17885, MEM_stage_inst_dmem_n17884, MEM_stage_inst_dmem_n17883, MEM_stage_inst_dmem_n17882, MEM_stage_inst_dmem_n17881, MEM_stage_inst_dmem_n17880, MEM_stage_inst_dmem_n17879, MEM_stage_inst_dmem_n17878, MEM_stage_inst_dmem_n17877, MEM_stage_inst_dmem_n17876, MEM_stage_inst_dmem_n17875, MEM_stage_inst_dmem_n17874, MEM_stage_inst_dmem_n17873, MEM_stage_inst_dmem_n17872, MEM_stage_inst_dmem_n17871, MEM_stage_inst_dmem_n17870, MEM_stage_inst_dmem_n17869, MEM_stage_inst_dmem_n17868, MEM_stage_inst_dmem_n17867, MEM_stage_inst_dmem_n17866, MEM_stage_inst_dmem_n17865, MEM_stage_inst_dmem_n17864, MEM_stage_inst_dmem_n17863, MEM_stage_inst_dmem_n17862, MEM_stage_inst_dmem_n17861, MEM_stage_inst_dmem_n17860, MEM_stage_inst_dmem_n17859, MEM_stage_inst_dmem_n17858, MEM_stage_inst_dmem_n17857, MEM_stage_inst_dmem_n17856, MEM_stage_inst_dmem_n17855, MEM_stage_inst_dmem_n17854, MEM_stage_inst_dmem_n17853, MEM_stage_inst_dmem_n17852, MEM_stage_inst_dmem_n17851, MEM_stage_inst_dmem_n17850, MEM_stage_inst_dmem_n17849, MEM_stage_inst_dmem_n17848, MEM_stage_inst_dmem_n17847, MEM_stage_inst_dmem_n17846, MEM_stage_inst_dmem_n17845, MEM_stage_inst_dmem_n17844, MEM_stage_inst_dmem_n17843, MEM_stage_inst_dmem_n17842, MEM_stage_inst_dmem_n17841, MEM_stage_inst_dmem_n17840, MEM_stage_inst_dmem_n17839, MEM_stage_inst_dmem_n17838, MEM_stage_inst_dmem_n17837, MEM_stage_inst_dmem_n17836, MEM_stage_inst_dmem_n17835, MEM_stage_inst_dmem_n17834, MEM_stage_inst_dmem_n17833, MEM_stage_inst_dmem_n17832, MEM_stage_inst_dmem_n17831, MEM_stage_inst_dmem_n17830, MEM_stage_inst_dmem_n17829, MEM_stage_inst_dmem_n17828, MEM_stage_inst_dmem_n17827, MEM_stage_inst_dmem_n17826, MEM_stage_inst_dmem_n17825, MEM_stage_inst_dmem_n17824, MEM_stage_inst_dmem_n17823, MEM_stage_inst_dmem_n17822, MEM_stage_inst_dmem_n17821, MEM_stage_inst_dmem_n17820, MEM_stage_inst_dmem_n17819, MEM_stage_inst_dmem_n17818, MEM_stage_inst_dmem_n17817, MEM_stage_inst_dmem_n17816, MEM_stage_inst_dmem_n17815, MEM_stage_inst_dmem_n17814, MEM_stage_inst_dmem_n17813, MEM_stage_inst_dmem_n17812, MEM_stage_inst_dmem_n17811, MEM_stage_inst_dmem_n17810, MEM_stage_inst_dmem_n17809, MEM_stage_inst_dmem_n17808, MEM_stage_inst_dmem_n17807, MEM_stage_inst_dmem_n17806, MEM_stage_inst_dmem_n17805, MEM_stage_inst_dmem_n17804, MEM_stage_inst_dmem_n17803, MEM_stage_inst_dmem_n17802, MEM_stage_inst_dmem_n17801, MEM_stage_inst_dmem_n17800, MEM_stage_inst_dmem_n17799, MEM_stage_inst_dmem_n17798, MEM_stage_inst_dmem_n17797, MEM_stage_inst_dmem_n17796, MEM_stage_inst_dmem_n17795, MEM_stage_inst_dmem_n17794, MEM_stage_inst_dmem_n17793, MEM_stage_inst_dmem_n17792, MEM_stage_inst_dmem_n17791, MEM_stage_inst_dmem_n17790, MEM_stage_inst_dmem_n17789, MEM_stage_inst_dmem_n17788, MEM_stage_inst_dmem_n17787, MEM_stage_inst_dmem_n17786, MEM_stage_inst_dmem_n17785, MEM_stage_inst_dmem_n17784, MEM_stage_inst_dmem_n17783, MEM_stage_inst_dmem_n17782, MEM_stage_inst_dmem_n17781, MEM_stage_inst_dmem_n17780, MEM_stage_inst_dmem_n17779, MEM_stage_inst_dmem_n17778, MEM_stage_inst_dmem_n17777, MEM_stage_inst_dmem_n17776, MEM_stage_inst_dmem_n17775, MEM_stage_inst_dmem_n17774, MEM_stage_inst_dmem_n17773, MEM_stage_inst_dmem_n17772, MEM_stage_inst_dmem_n17771, MEM_stage_inst_dmem_n17770, MEM_stage_inst_dmem_n17769, MEM_stage_inst_dmem_n17768, MEM_stage_inst_dmem_n17767, MEM_stage_inst_dmem_n17766, MEM_stage_inst_dmem_n17765, MEM_stage_inst_dmem_n17764, MEM_stage_inst_dmem_n17763, MEM_stage_inst_dmem_n17762, MEM_stage_inst_dmem_n17761, MEM_stage_inst_dmem_n17760, MEM_stage_inst_dmem_n17759, MEM_stage_inst_dmem_n17758, MEM_stage_inst_dmem_n17757, MEM_stage_inst_dmem_n17756, MEM_stage_inst_dmem_n17755, MEM_stage_inst_dmem_n17754, MEM_stage_inst_dmem_n17753, MEM_stage_inst_dmem_n17752, MEM_stage_inst_dmem_n17751, MEM_stage_inst_dmem_n17750, MEM_stage_inst_dmem_n17749, MEM_stage_inst_dmem_n17748, MEM_stage_inst_dmem_n17747, MEM_stage_inst_dmem_n17746, MEM_stage_inst_dmem_n17745, MEM_stage_inst_dmem_n17744, MEM_stage_inst_dmem_n17743, MEM_stage_inst_dmem_n17742, MEM_stage_inst_dmem_n17741, MEM_stage_inst_dmem_n17740, MEM_stage_inst_dmem_n17739, MEM_stage_inst_dmem_n17738, MEM_stage_inst_dmem_n17737, MEM_stage_inst_dmem_n17736, MEM_stage_inst_dmem_n17735, MEM_stage_inst_dmem_n17734, MEM_stage_inst_dmem_n17733, MEM_stage_inst_dmem_n17732, MEM_stage_inst_dmem_n17731, MEM_stage_inst_dmem_n17730, MEM_stage_inst_dmem_n17729, MEM_stage_inst_dmem_n17728, MEM_stage_inst_dmem_n17727, MEM_stage_inst_dmem_n17726, MEM_stage_inst_dmem_n17725, MEM_stage_inst_dmem_n17724, MEM_stage_inst_dmem_n17723, MEM_stage_inst_dmem_n17722, MEM_stage_inst_dmem_n17721, MEM_stage_inst_dmem_n17720, MEM_stage_inst_dmem_n17719, MEM_stage_inst_dmem_n17718, MEM_stage_inst_dmem_n17717, MEM_stage_inst_dmem_n17716, MEM_stage_inst_dmem_n17715, MEM_stage_inst_dmem_n17714, MEM_stage_inst_dmem_n17713, MEM_stage_inst_dmem_n17712, MEM_stage_inst_dmem_n17711, MEM_stage_inst_dmem_n17710, MEM_stage_inst_dmem_n17709, MEM_stage_inst_dmem_n17708, MEM_stage_inst_dmem_n17707, MEM_stage_inst_dmem_n17706, MEM_stage_inst_dmem_n17705, MEM_stage_inst_dmem_n17704, MEM_stage_inst_dmem_n17703, MEM_stage_inst_dmem_n17702, MEM_stage_inst_dmem_n17701, MEM_stage_inst_dmem_n17700, MEM_stage_inst_dmem_n17699, MEM_stage_inst_dmem_n17698, MEM_stage_inst_dmem_n17697, MEM_stage_inst_dmem_n17696, MEM_stage_inst_dmem_n17695, MEM_stage_inst_dmem_n17694, MEM_stage_inst_dmem_n17693, MEM_stage_inst_dmem_n17692, MEM_stage_inst_dmem_n17691, MEM_stage_inst_dmem_n17690, MEM_stage_inst_dmem_n17689, MEM_stage_inst_dmem_n17688, MEM_stage_inst_dmem_n17687, MEM_stage_inst_dmem_n17686, MEM_stage_inst_dmem_n17685, MEM_stage_inst_dmem_n17684, MEM_stage_inst_dmem_n17683, MEM_stage_inst_dmem_n17682, MEM_stage_inst_dmem_n17681, MEM_stage_inst_dmem_n17680, MEM_stage_inst_dmem_n17679, MEM_stage_inst_dmem_n17678, MEM_stage_inst_dmem_n17677, MEM_stage_inst_dmem_n17676, MEM_stage_inst_dmem_n17675, MEM_stage_inst_dmem_n17674, MEM_stage_inst_dmem_n17673, MEM_stage_inst_dmem_n17672, MEM_stage_inst_dmem_n17671, MEM_stage_inst_dmem_n17670, MEM_stage_inst_dmem_n17669, MEM_stage_inst_dmem_n17668, MEM_stage_inst_dmem_n17667, MEM_stage_inst_dmem_n17666, MEM_stage_inst_dmem_n17665, MEM_stage_inst_dmem_n17664, MEM_stage_inst_dmem_n17663, MEM_stage_inst_dmem_n17662, MEM_stage_inst_dmem_n17661, MEM_stage_inst_dmem_n17660, MEM_stage_inst_dmem_n17659, MEM_stage_inst_dmem_n17658, MEM_stage_inst_dmem_n17657, MEM_stage_inst_dmem_n17656, MEM_stage_inst_dmem_n17655, MEM_stage_inst_dmem_n17654, MEM_stage_inst_dmem_n17653, MEM_stage_inst_dmem_n17652, MEM_stage_inst_dmem_n17651, MEM_stage_inst_dmem_n17650, MEM_stage_inst_dmem_n17649, MEM_stage_inst_dmem_n17648, MEM_stage_inst_dmem_n17647, MEM_stage_inst_dmem_n17646, MEM_stage_inst_dmem_n17645, MEM_stage_inst_dmem_n17644, MEM_stage_inst_dmem_n17643, MEM_stage_inst_dmem_n17642, MEM_stage_inst_dmem_n17641, MEM_stage_inst_dmem_n17640, MEM_stage_inst_dmem_n17639, MEM_stage_inst_dmem_n17638, MEM_stage_inst_dmem_n17637, MEM_stage_inst_dmem_n17636, MEM_stage_inst_dmem_n17635, MEM_stage_inst_dmem_n17634, MEM_stage_inst_dmem_n17633, MEM_stage_inst_dmem_n17632, MEM_stage_inst_dmem_n17631, MEM_stage_inst_dmem_n17630, MEM_stage_inst_dmem_n17629, MEM_stage_inst_dmem_n17628, MEM_stage_inst_dmem_n17627, MEM_stage_inst_dmem_n17626, MEM_stage_inst_dmem_n17625, MEM_stage_inst_dmem_n17624, MEM_stage_inst_dmem_n17623, MEM_stage_inst_dmem_n17622, MEM_stage_inst_dmem_n17621, MEM_stage_inst_dmem_n17620, MEM_stage_inst_dmem_n17619, MEM_stage_inst_dmem_n17618, MEM_stage_inst_dmem_n17617, MEM_stage_inst_dmem_n17616, MEM_stage_inst_dmem_n17615, MEM_stage_inst_dmem_n17614, MEM_stage_inst_dmem_n17613, MEM_stage_inst_dmem_n17612, MEM_stage_inst_dmem_n17611, MEM_stage_inst_dmem_n17610, MEM_stage_inst_dmem_n17609, MEM_stage_inst_dmem_n17608, MEM_stage_inst_dmem_n17607, MEM_stage_inst_dmem_n17606, MEM_stage_inst_dmem_n17605, MEM_stage_inst_dmem_n17604, MEM_stage_inst_dmem_n17603, MEM_stage_inst_dmem_n17602, MEM_stage_inst_dmem_n17601, MEM_stage_inst_dmem_n17600, MEM_stage_inst_dmem_n17599, MEM_stage_inst_dmem_n17598, MEM_stage_inst_dmem_n17597, MEM_stage_inst_dmem_n17596, MEM_stage_inst_dmem_n17595, MEM_stage_inst_dmem_n17594, MEM_stage_inst_dmem_n17593, MEM_stage_inst_dmem_n17592, MEM_stage_inst_dmem_n17591, MEM_stage_inst_dmem_n17590, MEM_stage_inst_dmem_n17589, MEM_stage_inst_dmem_n17588, MEM_stage_inst_dmem_n17587, MEM_stage_inst_dmem_n17586, MEM_stage_inst_dmem_n17585, MEM_stage_inst_dmem_n17584, MEM_stage_inst_dmem_n17583, MEM_stage_inst_dmem_n17582, MEM_stage_inst_dmem_n17581, MEM_stage_inst_dmem_n17580, MEM_stage_inst_dmem_n17579, MEM_stage_inst_dmem_n17578, MEM_stage_inst_dmem_n17577, MEM_stage_inst_dmem_n17576, MEM_stage_inst_dmem_n17575, MEM_stage_inst_dmem_n17574, MEM_stage_inst_dmem_n17573, MEM_stage_inst_dmem_n17572, MEM_stage_inst_dmem_n17571, MEM_stage_inst_dmem_n17570, MEM_stage_inst_dmem_n17569, MEM_stage_inst_dmem_n17568, MEM_stage_inst_dmem_n17567, MEM_stage_inst_dmem_n17566, MEM_stage_inst_dmem_n17565, MEM_stage_inst_dmem_n17564, MEM_stage_inst_dmem_n17563, MEM_stage_inst_dmem_n17562, MEM_stage_inst_dmem_n17561, MEM_stage_inst_dmem_n17560, MEM_stage_inst_dmem_n17559, MEM_stage_inst_dmem_n17558, MEM_stage_inst_dmem_n17557, MEM_stage_inst_dmem_n17556, MEM_stage_inst_dmem_n17555, MEM_stage_inst_dmem_n17554, MEM_stage_inst_dmem_n17553, MEM_stage_inst_dmem_n17552, MEM_stage_inst_dmem_n17551, MEM_stage_inst_dmem_n17550, MEM_stage_inst_dmem_n17549, MEM_stage_inst_dmem_n17548, MEM_stage_inst_dmem_n17547, MEM_stage_inst_dmem_n17546, MEM_stage_inst_dmem_n17545, MEM_stage_inst_dmem_n17544, MEM_stage_inst_dmem_n17543, MEM_stage_inst_dmem_n17542, MEM_stage_inst_dmem_n17541, MEM_stage_inst_dmem_n17540, MEM_stage_inst_dmem_n17539, MEM_stage_inst_dmem_n17538, MEM_stage_inst_dmem_n17537, MEM_stage_inst_dmem_n17536, MEM_stage_inst_dmem_n17535, MEM_stage_inst_dmem_n17534, MEM_stage_inst_dmem_n17533, MEM_stage_inst_dmem_n17532, MEM_stage_inst_dmem_n17531, MEM_stage_inst_dmem_n17530, MEM_stage_inst_dmem_n17529, MEM_stage_inst_dmem_n17528, MEM_stage_inst_dmem_n17527, MEM_stage_inst_dmem_n17526, MEM_stage_inst_dmem_n17525, MEM_stage_inst_dmem_n17524, MEM_stage_inst_dmem_n17523, MEM_stage_inst_dmem_n17522, MEM_stage_inst_dmem_n17521, MEM_stage_inst_dmem_n17520, MEM_stage_inst_dmem_n17519, MEM_stage_inst_dmem_n17518, MEM_stage_inst_dmem_n17517, MEM_stage_inst_dmem_n17516, MEM_stage_inst_dmem_n17515, MEM_stage_inst_dmem_n17514, MEM_stage_inst_dmem_n17513, MEM_stage_inst_dmem_n17512, MEM_stage_inst_dmem_n17511, MEM_stage_inst_dmem_n17510, MEM_stage_inst_dmem_n17509, MEM_stage_inst_dmem_n17508, MEM_stage_inst_dmem_n17507, MEM_stage_inst_dmem_n17506, MEM_stage_inst_dmem_n17505, MEM_stage_inst_dmem_n17504, MEM_stage_inst_dmem_n17503, MEM_stage_inst_dmem_n17502, MEM_stage_inst_dmem_n17501, MEM_stage_inst_dmem_n17500, MEM_stage_inst_dmem_n17499, MEM_stage_inst_dmem_n17498, MEM_stage_inst_dmem_n17497, MEM_stage_inst_dmem_n17496, MEM_stage_inst_dmem_n17495, MEM_stage_inst_dmem_n17494, MEM_stage_inst_dmem_n17493, MEM_stage_inst_dmem_n17492, MEM_stage_inst_dmem_n17491, MEM_stage_inst_dmem_n17490, MEM_stage_inst_dmem_n17489, MEM_stage_inst_dmem_n17488, MEM_stage_inst_dmem_n17487, MEM_stage_inst_dmem_n17486, MEM_stage_inst_dmem_n17485, MEM_stage_inst_dmem_n17484, MEM_stage_inst_dmem_n17483, MEM_stage_inst_dmem_n17482, MEM_stage_inst_dmem_n17481, MEM_stage_inst_dmem_n17480, MEM_stage_inst_dmem_n17479, MEM_stage_inst_dmem_n17478, MEM_stage_inst_dmem_n17477, MEM_stage_inst_dmem_n17476, MEM_stage_inst_dmem_n17475, MEM_stage_inst_dmem_n17474, MEM_stage_inst_dmem_n17473, MEM_stage_inst_dmem_n17472, MEM_stage_inst_dmem_n17471, MEM_stage_inst_dmem_n17470, MEM_stage_inst_dmem_n17469, MEM_stage_inst_dmem_n17468, MEM_stage_inst_dmem_n17467, MEM_stage_inst_dmem_n17466, MEM_stage_inst_dmem_n17465, MEM_stage_inst_dmem_n17464, MEM_stage_inst_dmem_n17463, MEM_stage_inst_dmem_n17462, MEM_stage_inst_dmem_n17461, MEM_stage_inst_dmem_n17460, MEM_stage_inst_dmem_n17459, MEM_stage_inst_dmem_n17458, MEM_stage_inst_dmem_n17457, MEM_stage_inst_dmem_n17456, MEM_stage_inst_dmem_n17455, MEM_stage_inst_dmem_n17454, MEM_stage_inst_dmem_n17453, MEM_stage_inst_dmem_n17452, MEM_stage_inst_dmem_n17451, MEM_stage_inst_dmem_n17450, MEM_stage_inst_dmem_n17449, MEM_stage_inst_dmem_n17448, MEM_stage_inst_dmem_n17447, MEM_stage_inst_dmem_n17446, MEM_stage_inst_dmem_n17445, MEM_stage_inst_dmem_n17444, MEM_stage_inst_dmem_n17443, MEM_stage_inst_dmem_n17442, MEM_stage_inst_dmem_n17441, MEM_stage_inst_dmem_n17440, MEM_stage_inst_dmem_n17439, MEM_stage_inst_dmem_n17438, MEM_stage_inst_dmem_n17437, MEM_stage_inst_dmem_n17436, MEM_stage_inst_dmem_n17435, MEM_stage_inst_dmem_n17434, MEM_stage_inst_dmem_n17433, MEM_stage_inst_dmem_n17432, MEM_stage_inst_dmem_n17431, MEM_stage_inst_dmem_n17430, MEM_stage_inst_dmem_n17429, MEM_stage_inst_dmem_n17428, MEM_stage_inst_dmem_n17427, MEM_stage_inst_dmem_n17426, MEM_stage_inst_dmem_n17425, MEM_stage_inst_dmem_n17424, MEM_stage_inst_dmem_n17423, MEM_stage_inst_dmem_n17422, MEM_stage_inst_dmem_n17421, MEM_stage_inst_dmem_n17420, MEM_stage_inst_dmem_n17419, MEM_stage_inst_dmem_n17418, MEM_stage_inst_dmem_n17417, MEM_stage_inst_dmem_n17416, MEM_stage_inst_dmem_n17415, MEM_stage_inst_dmem_n17414, MEM_stage_inst_dmem_n17413, MEM_stage_inst_dmem_n17412, MEM_stage_inst_dmem_n17411, MEM_stage_inst_dmem_n17410, MEM_stage_inst_dmem_n17409, MEM_stage_inst_dmem_n17408, MEM_stage_inst_dmem_n17407, MEM_stage_inst_dmem_n17406, MEM_stage_inst_dmem_n17405, MEM_stage_inst_dmem_n17404, MEM_stage_inst_dmem_n17403, MEM_stage_inst_dmem_n17402, MEM_stage_inst_dmem_n17401, MEM_stage_inst_dmem_n17400, MEM_stage_inst_dmem_n17399, MEM_stage_inst_dmem_n17398, MEM_stage_inst_dmem_n17397, MEM_stage_inst_dmem_n17396, MEM_stage_inst_dmem_n17395, MEM_stage_inst_dmem_n17394, MEM_stage_inst_dmem_n17393, MEM_stage_inst_dmem_n17392, MEM_stage_inst_dmem_n17391, MEM_stage_inst_dmem_n17390, MEM_stage_inst_dmem_n17389, MEM_stage_inst_dmem_n17388, MEM_stage_inst_dmem_n17387, MEM_stage_inst_dmem_n17386, MEM_stage_inst_dmem_n17385, MEM_stage_inst_dmem_n17384, MEM_stage_inst_dmem_n17383, MEM_stage_inst_dmem_n17382, MEM_stage_inst_dmem_n17381, MEM_stage_inst_dmem_n17380, MEM_stage_inst_dmem_n17379, MEM_stage_inst_dmem_n17378, MEM_stage_inst_dmem_n17377, MEM_stage_inst_dmem_n17376, MEM_stage_inst_dmem_n17375, MEM_stage_inst_dmem_n17374, MEM_stage_inst_dmem_n17373, MEM_stage_inst_dmem_n17372, MEM_stage_inst_dmem_n17371, MEM_stage_inst_dmem_n17370, MEM_stage_inst_dmem_n17369, MEM_stage_inst_dmem_n17368, MEM_stage_inst_dmem_n17367, MEM_stage_inst_dmem_n17366, MEM_stage_inst_dmem_n17365, MEM_stage_inst_dmem_n17364, MEM_stage_inst_dmem_n17363, MEM_stage_inst_dmem_n17362, MEM_stage_inst_dmem_n17361, MEM_stage_inst_dmem_n17360, MEM_stage_inst_dmem_n17359, MEM_stage_inst_dmem_n17358, MEM_stage_inst_dmem_n17357, MEM_stage_inst_dmem_n17356, MEM_stage_inst_dmem_n17355, MEM_stage_inst_dmem_n17354, MEM_stage_inst_dmem_n17353, MEM_stage_inst_dmem_n17352, MEM_stage_inst_dmem_n17351, MEM_stage_inst_dmem_n17350, MEM_stage_inst_dmem_n17349, MEM_stage_inst_dmem_n17348, MEM_stage_inst_dmem_n17347, MEM_stage_inst_dmem_n17346, MEM_stage_inst_dmem_n17345, MEM_stage_inst_dmem_n17344, MEM_stage_inst_dmem_n17343, MEM_stage_inst_dmem_n17342, MEM_stage_inst_dmem_n17341, MEM_stage_inst_dmem_n17340, MEM_stage_inst_dmem_n17339, MEM_stage_inst_dmem_n17338, MEM_stage_inst_dmem_n17337, MEM_stage_inst_dmem_n17336, MEM_stage_inst_dmem_n17335, MEM_stage_inst_dmem_n17334, MEM_stage_inst_dmem_n17333, MEM_stage_inst_dmem_n17332, MEM_stage_inst_dmem_n17331, MEM_stage_inst_dmem_n17330, MEM_stage_inst_dmem_n17329, MEM_stage_inst_dmem_n17328, MEM_stage_inst_dmem_n17327, MEM_stage_inst_dmem_n17326, MEM_stage_inst_dmem_n17325, MEM_stage_inst_dmem_n17324, MEM_stage_inst_dmem_n17323, MEM_stage_inst_dmem_n17322, MEM_stage_inst_dmem_n17321, MEM_stage_inst_dmem_n17320, MEM_stage_inst_dmem_n17319, MEM_stage_inst_dmem_n17318, MEM_stage_inst_dmem_n17317, MEM_stage_inst_dmem_n17316, MEM_stage_inst_dmem_n17315, MEM_stage_inst_dmem_n17314, MEM_stage_inst_dmem_n17313, MEM_stage_inst_dmem_n17312, MEM_stage_inst_dmem_n17311, MEM_stage_inst_dmem_n17310, MEM_stage_inst_dmem_n17309, MEM_stage_inst_dmem_n17308, MEM_stage_inst_dmem_n17307, MEM_stage_inst_dmem_n17306, MEM_stage_inst_dmem_n17305, MEM_stage_inst_dmem_n17304, MEM_stage_inst_dmem_n17303, MEM_stage_inst_dmem_n17302, MEM_stage_inst_dmem_n17301, MEM_stage_inst_dmem_n17300, MEM_stage_inst_dmem_n17299, MEM_stage_inst_dmem_n17298, MEM_stage_inst_dmem_n17297, MEM_stage_inst_dmem_n17296, MEM_stage_inst_dmem_n17295, MEM_stage_inst_dmem_n17294, MEM_stage_inst_dmem_n17293, MEM_stage_inst_dmem_n17292, MEM_stage_inst_dmem_n17291, MEM_stage_inst_dmem_n17290, MEM_stage_inst_dmem_n17289, MEM_stage_inst_dmem_n17288, MEM_stage_inst_dmem_n17287, MEM_stage_inst_dmem_n17286, MEM_stage_inst_dmem_n17285, MEM_stage_inst_dmem_n17284, MEM_stage_inst_dmem_n17283, MEM_stage_inst_dmem_n17282, MEM_stage_inst_dmem_n17281, MEM_stage_inst_dmem_n17280, MEM_stage_inst_dmem_n17279, MEM_stage_inst_dmem_n17278, MEM_stage_inst_dmem_n17277, MEM_stage_inst_dmem_n17276, MEM_stage_inst_dmem_n17275, MEM_stage_inst_dmem_n17274, MEM_stage_inst_dmem_n17273, MEM_stage_inst_dmem_n17272, MEM_stage_inst_dmem_n17271, MEM_stage_inst_dmem_n17270, MEM_stage_inst_dmem_n17269, MEM_stage_inst_dmem_n17268, MEM_stage_inst_dmem_n17267, MEM_stage_inst_dmem_n17266, MEM_stage_inst_dmem_n17265, MEM_stage_inst_dmem_n17264, MEM_stage_inst_dmem_n17263, MEM_stage_inst_dmem_n17262, MEM_stage_inst_dmem_n17261, MEM_stage_inst_dmem_n17260, MEM_stage_inst_dmem_n17259, MEM_stage_inst_dmem_n17258, MEM_stage_inst_dmem_n17257, MEM_stage_inst_dmem_n17256, MEM_stage_inst_dmem_n17255, MEM_stage_inst_dmem_n17254, MEM_stage_inst_dmem_n17253, MEM_stage_inst_dmem_n17252, MEM_stage_inst_dmem_n17251, MEM_stage_inst_dmem_n17250, MEM_stage_inst_dmem_n17249, MEM_stage_inst_dmem_n17248, MEM_stage_inst_dmem_n17247, MEM_stage_inst_dmem_n17246, MEM_stage_inst_dmem_n17245, MEM_stage_inst_dmem_n17244, MEM_stage_inst_dmem_n17243, MEM_stage_inst_dmem_n17242, MEM_stage_inst_dmem_n17241, MEM_stage_inst_dmem_n17240, MEM_stage_inst_dmem_n17239, MEM_stage_inst_dmem_n17238, MEM_stage_inst_dmem_n17237, MEM_stage_inst_dmem_n17236, MEM_stage_inst_dmem_n17235, MEM_stage_inst_dmem_n17234, MEM_stage_inst_dmem_n17233, MEM_stage_inst_dmem_n17232, MEM_stage_inst_dmem_n17231, MEM_stage_inst_dmem_n17230, MEM_stage_inst_dmem_n17229, MEM_stage_inst_dmem_n17228, MEM_stage_inst_dmem_n17227, MEM_stage_inst_dmem_n17226, MEM_stage_inst_dmem_n17225, MEM_stage_inst_dmem_n17224, MEM_stage_inst_dmem_n17223, MEM_stage_inst_dmem_n17222, MEM_stage_inst_dmem_n17221, MEM_stage_inst_dmem_n17220, MEM_stage_inst_dmem_n17219, MEM_stage_inst_dmem_n17218, MEM_stage_inst_dmem_n17217, MEM_stage_inst_dmem_n17216, MEM_stage_inst_dmem_n17215, MEM_stage_inst_dmem_n17214, MEM_stage_inst_dmem_n17213, MEM_stage_inst_dmem_n17212, MEM_stage_inst_dmem_n17211, MEM_stage_inst_dmem_n17210, MEM_stage_inst_dmem_n17209, MEM_stage_inst_dmem_n17208, MEM_stage_inst_dmem_n17207, MEM_stage_inst_dmem_n17206, MEM_stage_inst_dmem_n17205, MEM_stage_inst_dmem_n17204, MEM_stage_inst_dmem_n17203, MEM_stage_inst_dmem_n17202, MEM_stage_inst_dmem_n17201, MEM_stage_inst_dmem_n17200, MEM_stage_inst_dmem_n17199, MEM_stage_inst_dmem_n17198, MEM_stage_inst_dmem_n17197, MEM_stage_inst_dmem_n17196, MEM_stage_inst_dmem_n17195, MEM_stage_inst_dmem_n17194, MEM_stage_inst_dmem_n17193, MEM_stage_inst_dmem_n17192, MEM_stage_inst_dmem_n17191, MEM_stage_inst_dmem_n17190, MEM_stage_inst_dmem_n17189, MEM_stage_inst_dmem_n17188, MEM_stage_inst_dmem_n17187, MEM_stage_inst_dmem_n17186, MEM_stage_inst_dmem_n17185, MEM_stage_inst_dmem_n17184, MEM_stage_inst_dmem_n17183, MEM_stage_inst_dmem_n17182, MEM_stage_inst_dmem_n17181, MEM_stage_inst_dmem_n17180, MEM_stage_inst_dmem_n17179, MEM_stage_inst_dmem_n17178, MEM_stage_inst_dmem_n17177, MEM_stage_inst_dmem_n17176, MEM_stage_inst_dmem_n17175, MEM_stage_inst_dmem_n17174, MEM_stage_inst_dmem_n17173, MEM_stage_inst_dmem_n17172, MEM_stage_inst_dmem_n17171, MEM_stage_inst_dmem_n17170, MEM_stage_inst_dmem_n17169, MEM_stage_inst_dmem_n17168, MEM_stage_inst_dmem_n17167, MEM_stage_inst_dmem_n17166, MEM_stage_inst_dmem_n17165, MEM_stage_inst_dmem_n17164, MEM_stage_inst_dmem_n17163, MEM_stage_inst_dmem_n17162, MEM_stage_inst_dmem_n17161, MEM_stage_inst_dmem_n17160, MEM_stage_inst_dmem_n17159, MEM_stage_inst_dmem_n17158, MEM_stage_inst_dmem_n17157, MEM_stage_inst_dmem_n17156, MEM_stage_inst_dmem_n17155, MEM_stage_inst_dmem_n17154, MEM_stage_inst_dmem_n17153, MEM_stage_inst_dmem_n17152, MEM_stage_inst_dmem_n17151, MEM_stage_inst_dmem_n17150, MEM_stage_inst_dmem_n17149, MEM_stage_inst_dmem_n17148, MEM_stage_inst_dmem_n17147, MEM_stage_inst_dmem_n17146, MEM_stage_inst_dmem_n17145, MEM_stage_inst_dmem_n17144, MEM_stage_inst_dmem_n17143, MEM_stage_inst_dmem_n17142, MEM_stage_inst_dmem_n17141, MEM_stage_inst_dmem_n17140, MEM_stage_inst_dmem_n17139, MEM_stage_inst_dmem_n17138, MEM_stage_inst_dmem_n17137, MEM_stage_inst_dmem_n17136, MEM_stage_inst_dmem_n17135, MEM_stage_inst_dmem_n17134, MEM_stage_inst_dmem_n17133, MEM_stage_inst_dmem_n17132, MEM_stage_inst_dmem_n17131, MEM_stage_inst_dmem_n17130, MEM_stage_inst_dmem_n17129, MEM_stage_inst_dmem_n17128, MEM_stage_inst_dmem_n17127, MEM_stage_inst_dmem_n17126, MEM_stage_inst_dmem_n17125, MEM_stage_inst_dmem_n17124, MEM_stage_inst_dmem_n17123, MEM_stage_inst_dmem_n17122, MEM_stage_inst_dmem_n17121, MEM_stage_inst_dmem_n17120, MEM_stage_inst_dmem_n17119, MEM_stage_inst_dmem_n17118, MEM_stage_inst_dmem_n17117, MEM_stage_inst_dmem_n17116, MEM_stage_inst_dmem_n17115, MEM_stage_inst_dmem_n17114, MEM_stage_inst_dmem_n17113, MEM_stage_inst_dmem_n17112, MEM_stage_inst_dmem_n17111, MEM_stage_inst_dmem_n17110, MEM_stage_inst_dmem_n17109, MEM_stage_inst_dmem_n17108, MEM_stage_inst_dmem_n17107, MEM_stage_inst_dmem_n17106, MEM_stage_inst_dmem_n17105, MEM_stage_inst_dmem_n17104, MEM_stage_inst_dmem_n17103, MEM_stage_inst_dmem_n17102, MEM_stage_inst_dmem_n17101, MEM_stage_inst_dmem_n17100, MEM_stage_inst_dmem_n17099, MEM_stage_inst_dmem_n17098, MEM_stage_inst_dmem_n17097, MEM_stage_inst_dmem_n17096, MEM_stage_inst_dmem_n17095, MEM_stage_inst_dmem_n17094, MEM_stage_inst_dmem_n17093, MEM_stage_inst_dmem_n17092, MEM_stage_inst_dmem_n17091, MEM_stage_inst_dmem_n17090, MEM_stage_inst_dmem_n17089, MEM_stage_inst_dmem_n17088, MEM_stage_inst_dmem_n17087, MEM_stage_inst_dmem_n17086, MEM_stage_inst_dmem_n17085, MEM_stage_inst_dmem_n17084, MEM_stage_inst_dmem_n17083, MEM_stage_inst_dmem_n17082, MEM_stage_inst_dmem_n17081, MEM_stage_inst_dmem_n17080, MEM_stage_inst_dmem_n17079, MEM_stage_inst_dmem_n17078, MEM_stage_inst_dmem_n17077, MEM_stage_inst_dmem_n17076, MEM_stage_inst_dmem_n17075, MEM_stage_inst_dmem_n17074, MEM_stage_inst_dmem_n17073, MEM_stage_inst_dmem_n17072, MEM_stage_inst_dmem_n17071, MEM_stage_inst_dmem_n17070, MEM_stage_inst_dmem_n17069, MEM_stage_inst_dmem_n17068, MEM_stage_inst_dmem_n17067, MEM_stage_inst_dmem_n17066, MEM_stage_inst_dmem_n17065, MEM_stage_inst_dmem_n17064, MEM_stage_inst_dmem_n17063, MEM_stage_inst_dmem_n17062, MEM_stage_inst_dmem_n17061, MEM_stage_inst_dmem_n17060, MEM_stage_inst_dmem_n17059, MEM_stage_inst_dmem_n17058, MEM_stage_inst_dmem_n17057, MEM_stage_inst_dmem_n17056, MEM_stage_inst_dmem_n17055, MEM_stage_inst_dmem_n17054, MEM_stage_inst_dmem_n17053, MEM_stage_inst_dmem_n17052, MEM_stage_inst_dmem_n17051, MEM_stage_inst_dmem_n17050, MEM_stage_inst_dmem_n17049, MEM_stage_inst_dmem_n17048, MEM_stage_inst_dmem_n17047, MEM_stage_inst_dmem_n17046, MEM_stage_inst_dmem_n17045, MEM_stage_inst_dmem_n17044, MEM_stage_inst_dmem_n17043, MEM_stage_inst_dmem_n17042, MEM_stage_inst_dmem_n17041, MEM_stage_inst_dmem_n17040, MEM_stage_inst_dmem_n17039, MEM_stage_inst_dmem_n17038, MEM_stage_inst_dmem_n17037, MEM_stage_inst_dmem_n17036, MEM_stage_inst_dmem_n17035, MEM_stage_inst_dmem_n17034, MEM_stage_inst_dmem_n17033, MEM_stage_inst_dmem_n17032, MEM_stage_inst_dmem_n17031, MEM_stage_inst_dmem_n17030, MEM_stage_inst_dmem_n17029, MEM_stage_inst_dmem_n17028, MEM_stage_inst_dmem_n17027, MEM_stage_inst_dmem_n17026, MEM_stage_inst_dmem_n17025, MEM_stage_inst_dmem_n17024, MEM_stage_inst_dmem_n17023, MEM_stage_inst_dmem_n17022, MEM_stage_inst_dmem_n17021, MEM_stage_inst_dmem_n17020, MEM_stage_inst_dmem_n17019, MEM_stage_inst_dmem_n17018, MEM_stage_inst_dmem_n17017, MEM_stage_inst_dmem_n17016, MEM_stage_inst_dmem_n17015, MEM_stage_inst_dmem_n17014, MEM_stage_inst_dmem_n17013, MEM_stage_inst_dmem_n17012, MEM_stage_inst_dmem_n17011, MEM_stage_inst_dmem_n17010, MEM_stage_inst_dmem_n17009, MEM_stage_inst_dmem_n17008, MEM_stage_inst_dmem_n17007, MEM_stage_inst_dmem_n17006, MEM_stage_inst_dmem_n17005, MEM_stage_inst_dmem_n17004, MEM_stage_inst_dmem_n17003, MEM_stage_inst_dmem_n17002, MEM_stage_inst_dmem_n17001, MEM_stage_inst_dmem_n17000, MEM_stage_inst_dmem_n16999, MEM_stage_inst_dmem_n16998, MEM_stage_inst_dmem_n16997, MEM_stage_inst_dmem_n16996, MEM_stage_inst_dmem_n16995, MEM_stage_inst_dmem_n16994, MEM_stage_inst_dmem_n16993, MEM_stage_inst_dmem_n16992, MEM_stage_inst_dmem_n16991, MEM_stage_inst_dmem_n16990, MEM_stage_inst_dmem_n16989, MEM_stage_inst_dmem_n16988, MEM_stage_inst_dmem_n16987, MEM_stage_inst_dmem_n16986, MEM_stage_inst_dmem_n16985, MEM_stage_inst_dmem_n16984, MEM_stage_inst_dmem_n16983, MEM_stage_inst_dmem_n16982, MEM_stage_inst_dmem_n16981, MEM_stage_inst_dmem_n16980, MEM_stage_inst_dmem_n16979, MEM_stage_inst_dmem_n16978, MEM_stage_inst_dmem_n16977, MEM_stage_inst_dmem_n16976, MEM_stage_inst_dmem_n16975, MEM_stage_inst_dmem_n16974, MEM_stage_inst_dmem_n16973, MEM_stage_inst_dmem_n16972, MEM_stage_inst_dmem_n16971, MEM_stage_inst_dmem_n16970, MEM_stage_inst_dmem_n16969, MEM_stage_inst_dmem_n16968, MEM_stage_inst_dmem_n16967, MEM_stage_inst_dmem_n16966, MEM_stage_inst_dmem_n16965, MEM_stage_inst_dmem_n16964, MEM_stage_inst_dmem_n16963, MEM_stage_inst_dmem_n16962, MEM_stage_inst_dmem_n16961, MEM_stage_inst_dmem_n16960, MEM_stage_inst_dmem_n16959, MEM_stage_inst_dmem_n16958, MEM_stage_inst_dmem_n16957, MEM_stage_inst_dmem_n16956, MEM_stage_inst_dmem_n16955, MEM_stage_inst_dmem_n16954, MEM_stage_inst_dmem_n16953, MEM_stage_inst_dmem_n16952, MEM_stage_inst_dmem_n16951, MEM_stage_inst_dmem_n16950, MEM_stage_inst_dmem_n16949, MEM_stage_inst_dmem_n16948, MEM_stage_inst_dmem_n16947, MEM_stage_inst_dmem_n16946, MEM_stage_inst_dmem_n16945, MEM_stage_inst_dmem_n16944, MEM_stage_inst_dmem_n16943, MEM_stage_inst_dmem_n16942, MEM_stage_inst_dmem_n16941, MEM_stage_inst_dmem_n16940, MEM_stage_inst_dmem_n16939, MEM_stage_inst_dmem_n16938, MEM_stage_inst_dmem_n16937, MEM_stage_inst_dmem_n16936, MEM_stage_inst_dmem_n16935, MEM_stage_inst_dmem_n16934, MEM_stage_inst_dmem_n16933, MEM_stage_inst_dmem_n16932, MEM_stage_inst_dmem_n16931, MEM_stage_inst_dmem_n16930, MEM_stage_inst_dmem_n16929, MEM_stage_inst_dmem_n16928, MEM_stage_inst_dmem_n16927, MEM_stage_inst_dmem_n16926, MEM_stage_inst_dmem_n16925, MEM_stage_inst_dmem_n16924, MEM_stage_inst_dmem_n16923, MEM_stage_inst_dmem_n16922, MEM_stage_inst_dmem_n16921, MEM_stage_inst_dmem_n16920, MEM_stage_inst_dmem_n16919, MEM_stage_inst_dmem_n16918, MEM_stage_inst_dmem_n16917, MEM_stage_inst_dmem_n16916, MEM_stage_inst_dmem_n16915, MEM_stage_inst_dmem_n16914, MEM_stage_inst_dmem_n16913, MEM_stage_inst_dmem_n16912, MEM_stage_inst_dmem_n16911, MEM_stage_inst_dmem_n16910, MEM_stage_inst_dmem_n16909, MEM_stage_inst_dmem_n16908, MEM_stage_inst_dmem_n16907, MEM_stage_inst_dmem_n16906, MEM_stage_inst_dmem_n16905, MEM_stage_inst_dmem_n16904, MEM_stage_inst_dmem_n16903, MEM_stage_inst_dmem_n16902, MEM_stage_inst_dmem_n16901, MEM_stage_inst_dmem_n16900, MEM_stage_inst_dmem_n16899, MEM_stage_inst_dmem_n16898, MEM_stage_inst_dmem_n16897, MEM_stage_inst_dmem_n16896, MEM_stage_inst_dmem_n16895, MEM_stage_inst_dmem_n16894, MEM_stage_inst_dmem_n16893, MEM_stage_inst_dmem_n16892, MEM_stage_inst_dmem_n16891, MEM_stage_inst_dmem_n16890, MEM_stage_inst_dmem_n16889, MEM_stage_inst_dmem_n16888, MEM_stage_inst_dmem_n16887, MEM_stage_inst_dmem_n16886, MEM_stage_inst_dmem_n16885, MEM_stage_inst_dmem_n16884, MEM_stage_inst_dmem_n16883, MEM_stage_inst_dmem_n16882, MEM_stage_inst_dmem_n16881, MEM_stage_inst_dmem_n16880, MEM_stage_inst_dmem_n16879, MEM_stage_inst_dmem_n16878, MEM_stage_inst_dmem_n16877, MEM_stage_inst_dmem_n16876, MEM_stage_inst_dmem_n16875, MEM_stage_inst_dmem_n16874, MEM_stage_inst_dmem_n16873, MEM_stage_inst_dmem_n16872, MEM_stage_inst_dmem_n16871, MEM_stage_inst_dmem_n16870, MEM_stage_inst_dmem_n16869, MEM_stage_inst_dmem_n16868, MEM_stage_inst_dmem_n16867, MEM_stage_inst_dmem_n16866, MEM_stage_inst_dmem_n16865, MEM_stage_inst_dmem_n16864, MEM_stage_inst_dmem_n16863, MEM_stage_inst_dmem_n16862, MEM_stage_inst_dmem_n16861, MEM_stage_inst_dmem_n16860, MEM_stage_inst_dmem_n16859, MEM_stage_inst_dmem_n16858, MEM_stage_inst_dmem_n16857, MEM_stage_inst_dmem_n16856, MEM_stage_inst_dmem_n16855, MEM_stage_inst_dmem_n16854, MEM_stage_inst_dmem_n16853, MEM_stage_inst_dmem_n16852, MEM_stage_inst_dmem_n16851, MEM_stage_inst_dmem_n16850, MEM_stage_inst_dmem_n16849, MEM_stage_inst_dmem_n16848, MEM_stage_inst_dmem_n16847, MEM_stage_inst_dmem_n16846, MEM_stage_inst_dmem_n16845, MEM_stage_inst_dmem_n16844, MEM_stage_inst_dmem_n16843, MEM_stage_inst_dmem_n16842, MEM_stage_inst_dmem_n16841, MEM_stage_inst_dmem_n16840, MEM_stage_inst_dmem_n16839, MEM_stage_inst_dmem_n16838, MEM_stage_inst_dmem_n16837, MEM_stage_inst_dmem_n16836, MEM_stage_inst_dmem_n16835, MEM_stage_inst_dmem_n16834, MEM_stage_inst_dmem_n16833, MEM_stage_inst_dmem_n16832, MEM_stage_inst_dmem_n16831, MEM_stage_inst_dmem_n16830, MEM_stage_inst_dmem_n16829, MEM_stage_inst_dmem_n16828, MEM_stage_inst_dmem_n16827, MEM_stage_inst_dmem_n16826, MEM_stage_inst_dmem_n16825, MEM_stage_inst_dmem_n16824, MEM_stage_inst_dmem_n16823, MEM_stage_inst_dmem_n16822, MEM_stage_inst_dmem_n16821, MEM_stage_inst_dmem_n16820, MEM_stage_inst_dmem_n16819, MEM_stage_inst_dmem_n16818, MEM_stage_inst_dmem_n16817, MEM_stage_inst_dmem_n16816, MEM_stage_inst_dmem_n16815, MEM_stage_inst_dmem_n16814, MEM_stage_inst_dmem_n16813, MEM_stage_inst_dmem_n16812, MEM_stage_inst_dmem_n16811, MEM_stage_inst_dmem_n16810, MEM_stage_inst_dmem_n16809, MEM_stage_inst_dmem_n16808, MEM_stage_inst_dmem_n16807, MEM_stage_inst_dmem_n16806, MEM_stage_inst_dmem_n16805, MEM_stage_inst_dmem_n16804, MEM_stage_inst_dmem_n16803, MEM_stage_inst_dmem_n16802, MEM_stage_inst_dmem_n16801, MEM_stage_inst_dmem_n16800, MEM_stage_inst_dmem_n16799, MEM_stage_inst_dmem_n16798, MEM_stage_inst_dmem_n16797, MEM_stage_inst_dmem_n16796, MEM_stage_inst_dmem_n16795, MEM_stage_inst_dmem_n16794, MEM_stage_inst_dmem_n16793, MEM_stage_inst_dmem_n16791, MEM_stage_inst_dmem_n16790, MEM_stage_inst_dmem_n16789, MEM_stage_inst_dmem_n16788, MEM_stage_inst_dmem_n16787, MEM_stage_inst_dmem_n16786, MEM_stage_inst_dmem_n16785, MEM_stage_inst_dmem_n16784, MEM_stage_inst_dmem_n16783, MEM_stage_inst_dmem_n16782, MEM_stage_inst_dmem_n16781, MEM_stage_inst_dmem_n16780, MEM_stage_inst_dmem_n16779, MEM_stage_inst_dmem_n16778, MEM_stage_inst_dmem_n16777, MEM_stage_inst_dmem_n16776, MEM_stage_inst_dmem_n16775, MEM_stage_inst_dmem_n16774, MEM_stage_inst_dmem_n16773, MEM_stage_inst_dmem_n16772, MEM_stage_inst_dmem_n16771, MEM_stage_inst_dmem_n16770, MEM_stage_inst_dmem_n16769, MEM_stage_inst_dmem_n16768, MEM_stage_inst_dmem_n16767, MEM_stage_inst_dmem_n16766, MEM_stage_inst_dmem_n16765, MEM_stage_inst_dmem_n16764, MEM_stage_inst_dmem_n16763, MEM_stage_inst_dmem_n16762, MEM_stage_inst_dmem_n16761, MEM_stage_inst_dmem_n16760, MEM_stage_inst_dmem_n16759, MEM_stage_inst_dmem_n16758, MEM_stage_inst_dmem_n16757, MEM_stage_inst_dmem_n16756, MEM_stage_inst_dmem_n16755, MEM_stage_inst_dmem_n16754, MEM_stage_inst_dmem_n16753, MEM_stage_inst_dmem_n16752, MEM_stage_inst_dmem_n16751, MEM_stage_inst_dmem_n16750, MEM_stage_inst_dmem_n16749, MEM_stage_inst_dmem_n16748, MEM_stage_inst_dmem_n16747, MEM_stage_inst_dmem_n16746, MEM_stage_inst_dmem_n16745, MEM_stage_inst_dmem_n16744, MEM_stage_inst_dmem_n16743, MEM_stage_inst_dmem_n16742, MEM_stage_inst_dmem_n16741, MEM_stage_inst_dmem_n16740, MEM_stage_inst_dmem_n16739, MEM_stage_inst_dmem_n16738, MEM_stage_inst_dmem_n16737, MEM_stage_inst_dmem_n16736, MEM_stage_inst_dmem_n16735, MEM_stage_inst_dmem_n16734, MEM_stage_inst_dmem_n16733, MEM_stage_inst_dmem_n16732, MEM_stage_inst_dmem_n16731, MEM_stage_inst_dmem_n16730, MEM_stage_inst_dmem_n16729, MEM_stage_inst_dmem_n16728, MEM_stage_inst_dmem_n16727, MEM_stage_inst_dmem_n16726, MEM_stage_inst_dmem_n16725, MEM_stage_inst_dmem_n16724, MEM_stage_inst_dmem_n16723, MEM_stage_inst_dmem_n16722, MEM_stage_inst_dmem_n16721, MEM_stage_inst_dmem_n16720, MEM_stage_inst_dmem_n16719, MEM_stage_inst_dmem_n16718, MEM_stage_inst_dmem_n16717, MEM_stage_inst_dmem_n16716, MEM_stage_inst_dmem_n16715, MEM_stage_inst_dmem_n16714, MEM_stage_inst_dmem_n16713, MEM_stage_inst_dmem_n16712, MEM_stage_inst_dmem_n16711, MEM_stage_inst_dmem_n16710, MEM_stage_inst_dmem_n16709, MEM_stage_inst_dmem_n16708, MEM_stage_inst_dmem_n16707, MEM_stage_inst_dmem_n16706, MEM_stage_inst_dmem_n16705, MEM_stage_inst_dmem_n16704, MEM_stage_inst_dmem_n16703, MEM_stage_inst_dmem_n16702, MEM_stage_inst_dmem_n16701, MEM_stage_inst_dmem_n16700, MEM_stage_inst_dmem_n16699, MEM_stage_inst_dmem_n16698, MEM_stage_inst_dmem_n16697, MEM_stage_inst_dmem_n16696, MEM_stage_inst_dmem_n16695, MEM_stage_inst_dmem_n16694, MEM_stage_inst_dmem_n16693, MEM_stage_inst_dmem_n16692, MEM_stage_inst_dmem_n16691, MEM_stage_inst_dmem_n16690, MEM_stage_inst_dmem_n16689, MEM_stage_inst_dmem_n16688, MEM_stage_inst_dmem_n16687, MEM_stage_inst_dmem_n16686, MEM_stage_inst_dmem_n16685, MEM_stage_inst_dmem_n16684, MEM_stage_inst_dmem_n16683, MEM_stage_inst_dmem_n16682, MEM_stage_inst_dmem_n16681, MEM_stage_inst_dmem_n16680, MEM_stage_inst_dmem_n16679, MEM_stage_inst_dmem_n16678, MEM_stage_inst_dmem_n16677, MEM_stage_inst_dmem_n16676, MEM_stage_inst_dmem_n16675, MEM_stage_inst_dmem_n16674, MEM_stage_inst_dmem_n16673, MEM_stage_inst_dmem_n16672, MEM_stage_inst_dmem_n16671, MEM_stage_inst_dmem_n16670, MEM_stage_inst_dmem_n16669, MEM_stage_inst_dmem_n16668, MEM_stage_inst_dmem_n16667, MEM_stage_inst_dmem_n16666, MEM_stage_inst_dmem_n16665, MEM_stage_inst_dmem_n16664, MEM_stage_inst_dmem_n16663, MEM_stage_inst_dmem_n16662, MEM_stage_inst_dmem_n16661, MEM_stage_inst_dmem_n16660, MEM_stage_inst_dmem_n16659, MEM_stage_inst_dmem_n16658, MEM_stage_inst_dmem_n16657, MEM_stage_inst_dmem_n16656, MEM_stage_inst_dmem_n16655, MEM_stage_inst_dmem_n16654, MEM_stage_inst_dmem_n16653, MEM_stage_inst_dmem_n16652, MEM_stage_inst_dmem_n16651, MEM_stage_inst_dmem_n16650, MEM_stage_inst_dmem_n16649, MEM_stage_inst_dmem_n16648, MEM_stage_inst_dmem_n16647, MEM_stage_inst_dmem_n16646, MEM_stage_inst_dmem_n16645, MEM_stage_inst_dmem_n16644, MEM_stage_inst_dmem_n16643, MEM_stage_inst_dmem_n16642, MEM_stage_inst_dmem_n16641, MEM_stage_inst_dmem_n16640, MEM_stage_inst_dmem_n16639, MEM_stage_inst_dmem_n16638, MEM_stage_inst_dmem_n16637, MEM_stage_inst_dmem_n16636, MEM_stage_inst_dmem_n16635, MEM_stage_inst_dmem_n16634, MEM_stage_inst_dmem_n16633, MEM_stage_inst_dmem_n16632, MEM_stage_inst_dmem_n16631, MEM_stage_inst_dmem_n16630, MEM_stage_inst_dmem_n16629, MEM_stage_inst_dmem_n16628, MEM_stage_inst_dmem_n16627, MEM_stage_inst_dmem_n16626, MEM_stage_inst_dmem_n16625, MEM_stage_inst_dmem_n16624, MEM_stage_inst_dmem_n16623, MEM_stage_inst_dmem_n16622, MEM_stage_inst_dmem_n16621, MEM_stage_inst_dmem_n16620, MEM_stage_inst_dmem_n16619, MEM_stage_inst_dmem_n16618, MEM_stage_inst_dmem_n16617, MEM_stage_inst_dmem_n16616, MEM_stage_inst_dmem_n16615, MEM_stage_inst_dmem_n16614, MEM_stage_inst_dmem_n16613, MEM_stage_inst_dmem_n16612, MEM_stage_inst_dmem_n16611, MEM_stage_inst_dmem_n16610, MEM_stage_inst_dmem_n16609, MEM_stage_inst_dmem_n16608, MEM_stage_inst_dmem_n16607, MEM_stage_inst_dmem_n16606, MEM_stage_inst_dmem_n16605, MEM_stage_inst_dmem_n16604, MEM_stage_inst_dmem_n16603, MEM_stage_inst_dmem_n16602, MEM_stage_inst_dmem_n16601, MEM_stage_inst_dmem_n16600, MEM_stage_inst_dmem_n16599, MEM_stage_inst_dmem_n16598, MEM_stage_inst_dmem_n16597, MEM_stage_inst_dmem_n16596, MEM_stage_inst_dmem_n16595, MEM_stage_inst_dmem_n16594, MEM_stage_inst_dmem_n16593, MEM_stage_inst_dmem_n16592, MEM_stage_inst_dmem_n16591, MEM_stage_inst_dmem_n16590, MEM_stage_inst_dmem_n16589, MEM_stage_inst_dmem_n16588, MEM_stage_inst_dmem_n16587, MEM_stage_inst_dmem_n16586, MEM_stage_inst_dmem_n16585, MEM_stage_inst_dmem_n16584, MEM_stage_inst_dmem_n16583, MEM_stage_inst_dmem_n16582, MEM_stage_inst_dmem_n16581, MEM_stage_inst_dmem_n16580, MEM_stage_inst_dmem_n16579, MEM_stage_inst_dmem_n16578, MEM_stage_inst_dmem_n16577, MEM_stage_inst_dmem_n16576, MEM_stage_inst_dmem_n16575, MEM_stage_inst_dmem_n16574, MEM_stage_inst_dmem_n16573, MEM_stage_inst_dmem_n16572, MEM_stage_inst_dmem_n16571, MEM_stage_inst_dmem_n16570, MEM_stage_inst_dmem_n16569, MEM_stage_inst_dmem_n16568, MEM_stage_inst_dmem_n16567, MEM_stage_inst_dmem_n16566, MEM_stage_inst_dmem_n16565, MEM_stage_inst_dmem_n16564, MEM_stage_inst_dmem_n16563, MEM_stage_inst_dmem_n16562, MEM_stage_inst_dmem_n16561, MEM_stage_inst_dmem_n16560, MEM_stage_inst_dmem_n16559, MEM_stage_inst_dmem_n16558, MEM_stage_inst_dmem_n16557, MEM_stage_inst_dmem_n16556, MEM_stage_inst_dmem_n16555, MEM_stage_inst_dmem_n16554, MEM_stage_inst_dmem_n16553, MEM_stage_inst_dmem_n16552, MEM_stage_inst_dmem_n16551, MEM_stage_inst_dmem_n16550, MEM_stage_inst_dmem_n16549, MEM_stage_inst_dmem_n16548, MEM_stage_inst_dmem_n16547, MEM_stage_inst_dmem_n16546, MEM_stage_inst_dmem_n16545, MEM_stage_inst_dmem_n16544, MEM_stage_inst_dmem_n16543, MEM_stage_inst_dmem_n16542, MEM_stage_inst_dmem_n16541, MEM_stage_inst_dmem_n16540, MEM_stage_inst_dmem_n16539, MEM_stage_inst_dmem_n16538, MEM_stage_inst_dmem_n16537, MEM_stage_inst_dmem_n16536, MEM_stage_inst_dmem_n16535, MEM_stage_inst_dmem_n16534, MEM_stage_inst_dmem_n16533, MEM_stage_inst_dmem_n16532, MEM_stage_inst_dmem_n16531, MEM_stage_inst_dmem_n16530, MEM_stage_inst_dmem_n16529, MEM_stage_inst_dmem_n16528, MEM_stage_inst_dmem_n16527, MEM_stage_inst_dmem_n16526, MEM_stage_inst_dmem_n16525, MEM_stage_inst_dmem_n16524, MEM_stage_inst_dmem_n16523, MEM_stage_inst_dmem_n16522, MEM_stage_inst_dmem_n16521, MEM_stage_inst_dmem_n16520, MEM_stage_inst_dmem_n16519, MEM_stage_inst_dmem_n16518, MEM_stage_inst_dmem_n16517, MEM_stage_inst_dmem_n16516, MEM_stage_inst_dmem_n16515, MEM_stage_inst_dmem_n16514, MEM_stage_inst_dmem_n16513, MEM_stage_inst_dmem_n16512, MEM_stage_inst_dmem_n16511, MEM_stage_inst_dmem_n16510, MEM_stage_inst_dmem_n16509, MEM_stage_inst_dmem_n16508, MEM_stage_inst_dmem_n16507, MEM_stage_inst_dmem_n16506, MEM_stage_inst_dmem_n16505, MEM_stage_inst_dmem_n16504, MEM_stage_inst_dmem_n16503, MEM_stage_inst_dmem_n16502, MEM_stage_inst_dmem_n16501, MEM_stage_inst_dmem_n16500, MEM_stage_inst_dmem_n16499, MEM_stage_inst_dmem_n16498, MEM_stage_inst_dmem_n16497, MEM_stage_inst_dmem_n16496, MEM_stage_inst_dmem_n16495, MEM_stage_inst_dmem_n16494, MEM_stage_inst_dmem_n16493, MEM_stage_inst_dmem_n16492, MEM_stage_inst_dmem_n16491, MEM_stage_inst_dmem_n16490, MEM_stage_inst_dmem_n16489, MEM_stage_inst_dmem_n16488, MEM_stage_inst_dmem_n16487, MEM_stage_inst_dmem_n16486, MEM_stage_inst_dmem_n16485, MEM_stage_inst_dmem_n16484, MEM_stage_inst_dmem_n16483, MEM_stage_inst_dmem_n16482, MEM_stage_inst_dmem_n16481, MEM_stage_inst_dmem_n16480, MEM_stage_inst_dmem_n16479, MEM_stage_inst_dmem_n16478, MEM_stage_inst_dmem_n16477, MEM_stage_inst_dmem_n16476, MEM_stage_inst_dmem_n16475, MEM_stage_inst_dmem_n16474, MEM_stage_inst_dmem_n16473, MEM_stage_inst_dmem_n16472, MEM_stage_inst_dmem_n16471, MEM_stage_inst_dmem_n16470, MEM_stage_inst_dmem_n16469, MEM_stage_inst_dmem_n16468, MEM_stage_inst_dmem_n16467, MEM_stage_inst_dmem_n16466, MEM_stage_inst_dmem_n16465, MEM_stage_inst_dmem_n16464, MEM_stage_inst_dmem_n16463, MEM_stage_inst_dmem_n16462, MEM_stage_inst_dmem_n16461, MEM_stage_inst_dmem_n16460, MEM_stage_inst_dmem_n16459, MEM_stage_inst_dmem_n16458, MEM_stage_inst_dmem_n16457, MEM_stage_inst_dmem_n16456, MEM_stage_inst_dmem_n16455, MEM_stage_inst_dmem_n16454, MEM_stage_inst_dmem_n16453, MEM_stage_inst_dmem_n16452, MEM_stage_inst_dmem_n16451, MEM_stage_inst_dmem_n16450, MEM_stage_inst_dmem_n16449, MEM_stage_inst_dmem_n16448, MEM_stage_inst_dmem_n16447, MEM_stage_inst_dmem_n16446, MEM_stage_inst_dmem_n16445, MEM_stage_inst_dmem_n16444, MEM_stage_inst_dmem_n16443, MEM_stage_inst_dmem_n16442, MEM_stage_inst_dmem_n16441, MEM_stage_inst_dmem_n16440, MEM_stage_inst_dmem_n16439, MEM_stage_inst_dmem_n16438, MEM_stage_inst_dmem_n16437, MEM_stage_inst_dmem_n16436, MEM_stage_inst_dmem_n16435, MEM_stage_inst_dmem_n16434, MEM_stage_inst_dmem_n16433, MEM_stage_inst_dmem_n16432, MEM_stage_inst_dmem_n16431, MEM_stage_inst_dmem_n16430, MEM_stage_inst_dmem_n16429, MEM_stage_inst_dmem_n16428, MEM_stage_inst_dmem_n16427, MEM_stage_inst_dmem_n16426, MEM_stage_inst_dmem_n16425, MEM_stage_inst_dmem_n16424, MEM_stage_inst_dmem_n16423, MEM_stage_inst_dmem_n16422, MEM_stage_inst_dmem_n16421, MEM_stage_inst_dmem_n16420, MEM_stage_inst_dmem_n16419, MEM_stage_inst_dmem_n16418, MEM_stage_inst_dmem_n16417, MEM_stage_inst_dmem_n16416, MEM_stage_inst_dmem_n16415, MEM_stage_inst_dmem_n16414, MEM_stage_inst_dmem_n16413, MEM_stage_inst_dmem_n16412, MEM_stage_inst_dmem_n16411, MEM_stage_inst_dmem_n16410, MEM_stage_inst_dmem_n16409, MEM_stage_inst_dmem_n16408, MEM_stage_inst_dmem_n16407, MEM_stage_inst_dmem_n16406, MEM_stage_inst_dmem_n16405, MEM_stage_inst_dmem_n16404, MEM_stage_inst_dmem_n16403, MEM_stage_inst_dmem_n16402, MEM_stage_inst_dmem_n16401, MEM_stage_inst_dmem_n16400, MEM_stage_inst_dmem_n16399, MEM_stage_inst_dmem_n16398, MEM_stage_inst_dmem_n16397, MEM_stage_inst_dmem_n16396, MEM_stage_inst_dmem_n16395, MEM_stage_inst_dmem_n16394, MEM_stage_inst_dmem_n16393, MEM_stage_inst_dmem_n16392, MEM_stage_inst_dmem_n16391, MEM_stage_inst_dmem_n16390, MEM_stage_inst_dmem_n16389, MEM_stage_inst_dmem_n16388, MEM_stage_inst_dmem_n16387, MEM_stage_inst_dmem_n16386, MEM_stage_inst_dmem_n16385, MEM_stage_inst_dmem_n16384, MEM_stage_inst_dmem_n16383, MEM_stage_inst_dmem_n16382, MEM_stage_inst_dmem_n16381, MEM_stage_inst_dmem_n16380, MEM_stage_inst_dmem_n16379, MEM_stage_inst_dmem_n16378, MEM_stage_inst_dmem_n16377, MEM_stage_inst_dmem_n16376, MEM_stage_inst_dmem_n16375, MEM_stage_inst_dmem_n16374, MEM_stage_inst_dmem_n16373, MEM_stage_inst_dmem_n16372, MEM_stage_inst_dmem_n16371, MEM_stage_inst_dmem_n16370, MEM_stage_inst_dmem_n16369, MEM_stage_inst_dmem_n16368, MEM_stage_inst_dmem_n16367, MEM_stage_inst_dmem_n16366, MEM_stage_inst_dmem_n16365, MEM_stage_inst_dmem_n16364, MEM_stage_inst_dmem_n16363, MEM_stage_inst_dmem_n16362, MEM_stage_inst_dmem_n16361, MEM_stage_inst_dmem_n16360, MEM_stage_inst_dmem_n16359, MEM_stage_inst_dmem_n16358, MEM_stage_inst_dmem_n16357, MEM_stage_inst_dmem_n16356, MEM_stage_inst_dmem_n16355, MEM_stage_inst_dmem_n16354, MEM_stage_inst_dmem_n16353, MEM_stage_inst_dmem_n16352, MEM_stage_inst_dmem_n16351, MEM_stage_inst_dmem_n16350, MEM_stage_inst_dmem_n16349, MEM_stage_inst_dmem_n16348, MEM_stage_inst_dmem_n16347, MEM_stage_inst_dmem_n16346, MEM_stage_inst_dmem_n16345, MEM_stage_inst_dmem_n16344, MEM_stage_inst_dmem_n16343, MEM_stage_inst_dmem_n16342, MEM_stage_inst_dmem_n16341, MEM_stage_inst_dmem_n16340, MEM_stage_inst_dmem_n16339, MEM_stage_inst_dmem_n16338, MEM_stage_inst_dmem_n16337, MEM_stage_inst_dmem_n16336, MEM_stage_inst_dmem_n16335, MEM_stage_inst_dmem_n16334, MEM_stage_inst_dmem_n16333, MEM_stage_inst_dmem_n16332, MEM_stage_inst_dmem_n16331, MEM_stage_inst_dmem_n16330, MEM_stage_inst_dmem_n16329, MEM_stage_inst_dmem_n16328, MEM_stage_inst_dmem_n16327, MEM_stage_inst_dmem_n16326, MEM_stage_inst_dmem_n16325, MEM_stage_inst_dmem_n16324, MEM_stage_inst_dmem_n16323, MEM_stage_inst_dmem_n16322, MEM_stage_inst_dmem_n16321, MEM_stage_inst_dmem_n16320, MEM_stage_inst_dmem_n16319, MEM_stage_inst_dmem_n16318, MEM_stage_inst_dmem_n16317, MEM_stage_inst_dmem_n16316, MEM_stage_inst_dmem_n16315, MEM_stage_inst_dmem_n16314, MEM_stage_inst_dmem_n16313, MEM_stage_inst_dmem_n16312, MEM_stage_inst_dmem_n16311, MEM_stage_inst_dmem_n16310, MEM_stage_inst_dmem_n16309, MEM_stage_inst_dmem_n16308, MEM_stage_inst_dmem_n16307, MEM_stage_inst_dmem_n16306, MEM_stage_inst_dmem_n16305, MEM_stage_inst_dmem_n16304, MEM_stage_inst_dmem_n16303, MEM_stage_inst_dmem_n16302, MEM_stage_inst_dmem_n16301, MEM_stage_inst_dmem_n16300, MEM_stage_inst_dmem_n16299, MEM_stage_inst_dmem_n16298, MEM_stage_inst_dmem_n16297, MEM_stage_inst_dmem_n16296, MEM_stage_inst_dmem_n16295, MEM_stage_inst_dmem_n16294, MEM_stage_inst_dmem_n16293, MEM_stage_inst_dmem_n16292, MEM_stage_inst_dmem_n16291, MEM_stage_inst_dmem_n16290, MEM_stage_inst_dmem_n16289, MEM_stage_inst_dmem_n16288, MEM_stage_inst_dmem_n16287, MEM_stage_inst_dmem_n16286, MEM_stage_inst_dmem_n16285, MEM_stage_inst_dmem_n16284, MEM_stage_inst_dmem_n16283, MEM_stage_inst_dmem_n16282, MEM_stage_inst_dmem_n16281, MEM_stage_inst_dmem_n16280, MEM_stage_inst_dmem_n16279, MEM_stage_inst_dmem_n16278, MEM_stage_inst_dmem_n16277, MEM_stage_inst_dmem_n16276, MEM_stage_inst_dmem_n16275, MEM_stage_inst_dmem_n16274, MEM_stage_inst_dmem_n16273, MEM_stage_inst_dmem_n16272, MEM_stage_inst_dmem_n16271, MEM_stage_inst_dmem_n16270, MEM_stage_inst_dmem_n16269, MEM_stage_inst_dmem_n16268, MEM_stage_inst_dmem_n16267, MEM_stage_inst_dmem_n16266, MEM_stage_inst_dmem_n16265, MEM_stage_inst_dmem_n16264, MEM_stage_inst_dmem_n16263, MEM_stage_inst_dmem_n16262, MEM_stage_inst_dmem_n16261, MEM_stage_inst_dmem_n16260, MEM_stage_inst_dmem_n16259, MEM_stage_inst_dmem_n16258, MEM_stage_inst_dmem_n16257, MEM_stage_inst_dmem_n16256, MEM_stage_inst_dmem_n16255, MEM_stage_inst_dmem_n16254, MEM_stage_inst_dmem_n16253, MEM_stage_inst_dmem_n16252, MEM_stage_inst_dmem_n16251, MEM_stage_inst_dmem_n16250, MEM_stage_inst_dmem_n16249, MEM_stage_inst_dmem_n16248, MEM_stage_inst_dmem_n16247, MEM_stage_inst_dmem_n16246, MEM_stage_inst_dmem_n16245, MEM_stage_inst_dmem_n16244, MEM_stage_inst_dmem_n16243, MEM_stage_inst_dmem_n16242, MEM_stage_inst_dmem_n16241, MEM_stage_inst_dmem_n16240, MEM_stage_inst_dmem_n16239, MEM_stage_inst_dmem_n16238, MEM_stage_inst_dmem_n16237, MEM_stage_inst_dmem_n16236, MEM_stage_inst_dmem_n16235, MEM_stage_inst_dmem_n16234, MEM_stage_inst_dmem_n16233, MEM_stage_inst_dmem_n16232, MEM_stage_inst_dmem_n16231, MEM_stage_inst_dmem_n16230, MEM_stage_inst_dmem_n16229, MEM_stage_inst_dmem_n16228, MEM_stage_inst_dmem_n16227, MEM_stage_inst_dmem_n16226, MEM_stage_inst_dmem_n16225, MEM_stage_inst_dmem_n16224, MEM_stage_inst_dmem_n16223, MEM_stage_inst_dmem_n16222, MEM_stage_inst_dmem_n16221, MEM_stage_inst_dmem_n16220, MEM_stage_inst_dmem_n16219, MEM_stage_inst_dmem_n16218, MEM_stage_inst_dmem_n16217, MEM_stage_inst_dmem_n16216, MEM_stage_inst_dmem_n16215, MEM_stage_inst_dmem_n16214, MEM_stage_inst_dmem_n16213, MEM_stage_inst_dmem_n16212, MEM_stage_inst_dmem_n16211, MEM_stage_inst_dmem_n16210, MEM_stage_inst_dmem_n16209, MEM_stage_inst_dmem_n16208, MEM_stage_inst_dmem_n16207, MEM_stage_inst_dmem_n16206, MEM_stage_inst_dmem_n16205, MEM_stage_inst_dmem_n16204, MEM_stage_inst_dmem_n16203, MEM_stage_inst_dmem_n16202, MEM_stage_inst_dmem_n16201, MEM_stage_inst_dmem_n16200, MEM_stage_inst_dmem_n16199, MEM_stage_inst_dmem_n16198, MEM_stage_inst_dmem_n16197, MEM_stage_inst_dmem_n16196, MEM_stage_inst_dmem_n16195, MEM_stage_inst_dmem_n16194, MEM_stage_inst_dmem_n16193, MEM_stage_inst_dmem_n16192, MEM_stage_inst_dmem_n16191, MEM_stage_inst_dmem_n16190, MEM_stage_inst_dmem_n16189, MEM_stage_inst_dmem_n16188, MEM_stage_inst_dmem_n16187, MEM_stage_inst_dmem_n16186, MEM_stage_inst_dmem_n16185, MEM_stage_inst_dmem_n16184, MEM_stage_inst_dmem_n16183, MEM_stage_inst_dmem_n16182, MEM_stage_inst_dmem_n16181, MEM_stage_inst_dmem_n16180, MEM_stage_inst_dmem_n16179, MEM_stage_inst_dmem_n16178, MEM_stage_inst_dmem_n16177, MEM_stage_inst_dmem_n16176, MEM_stage_inst_dmem_n16175, MEM_stage_inst_dmem_n16174, MEM_stage_inst_dmem_n16173, MEM_stage_inst_dmem_n16172, MEM_stage_inst_dmem_n16171, MEM_stage_inst_dmem_n16170, MEM_stage_inst_dmem_n16169, MEM_stage_inst_dmem_n16168, MEM_stage_inst_dmem_n16167, MEM_stage_inst_dmem_n16166, MEM_stage_inst_dmem_n16165, MEM_stage_inst_dmem_n16164, MEM_stage_inst_dmem_n16163, MEM_stage_inst_dmem_n16162, MEM_stage_inst_dmem_n16161, MEM_stage_inst_dmem_n16160, MEM_stage_inst_dmem_n16159, MEM_stage_inst_dmem_n16158, MEM_stage_inst_dmem_n16157, MEM_stage_inst_dmem_n16156, MEM_stage_inst_dmem_n16155, MEM_stage_inst_dmem_n16154, MEM_stage_inst_dmem_n16153, MEM_stage_inst_dmem_n16152, MEM_stage_inst_dmem_n16151, MEM_stage_inst_dmem_n16150, MEM_stage_inst_dmem_n16149, MEM_stage_inst_dmem_n16148, MEM_stage_inst_dmem_n16147, MEM_stage_inst_dmem_n16146, MEM_stage_inst_dmem_n16145, MEM_stage_inst_dmem_n16144, MEM_stage_inst_dmem_n16143, MEM_stage_inst_dmem_n16142, MEM_stage_inst_dmem_n16141, MEM_stage_inst_dmem_n16140, MEM_stage_inst_dmem_n16139, MEM_stage_inst_dmem_n16138, MEM_stage_inst_dmem_n16137, MEM_stage_inst_dmem_n16136, MEM_stage_inst_dmem_n16135, MEM_stage_inst_dmem_n16134, MEM_stage_inst_dmem_n16133, MEM_stage_inst_dmem_n16132, MEM_stage_inst_dmem_n16131, MEM_stage_inst_dmem_n16130, MEM_stage_inst_dmem_n16129, MEM_stage_inst_dmem_n16128, MEM_stage_inst_dmem_n16127, MEM_stage_inst_dmem_n16126, MEM_stage_inst_dmem_n16125, MEM_stage_inst_dmem_n16124, MEM_stage_inst_dmem_n16123, MEM_stage_inst_dmem_n16122, MEM_stage_inst_dmem_n16121, MEM_stage_inst_dmem_n16120, MEM_stage_inst_dmem_n16119, MEM_stage_inst_dmem_n16118, MEM_stage_inst_dmem_n16117, MEM_stage_inst_dmem_n16116, MEM_stage_inst_dmem_n16115, MEM_stage_inst_dmem_n16114, MEM_stage_inst_dmem_n16113, MEM_stage_inst_dmem_n16112, MEM_stage_inst_dmem_n16111, MEM_stage_inst_dmem_n16110, MEM_stage_inst_dmem_n16109, MEM_stage_inst_dmem_n16108, MEM_stage_inst_dmem_n16107, MEM_stage_inst_dmem_n16106, MEM_stage_inst_dmem_n16105, MEM_stage_inst_dmem_n16104, MEM_stage_inst_dmem_n16103, MEM_stage_inst_dmem_n16102, MEM_stage_inst_dmem_n16101, MEM_stage_inst_dmem_n16100, MEM_stage_inst_dmem_n16099, MEM_stage_inst_dmem_n16098, MEM_stage_inst_dmem_n16097, MEM_stage_inst_dmem_n16096, MEM_stage_inst_dmem_n16095, MEM_stage_inst_dmem_n16094, MEM_stage_inst_dmem_n16093, MEM_stage_inst_dmem_n16092, MEM_stage_inst_dmem_n16091, MEM_stage_inst_dmem_n16090, MEM_stage_inst_dmem_n16089, MEM_stage_inst_dmem_n16088, MEM_stage_inst_dmem_n16087, MEM_stage_inst_dmem_n16086, MEM_stage_inst_dmem_n16085, MEM_stage_inst_dmem_n16084, MEM_stage_inst_dmem_n16083, MEM_stage_inst_dmem_n16082, MEM_stage_inst_dmem_n16081, MEM_stage_inst_dmem_n16080, MEM_stage_inst_dmem_n16079, MEM_stage_inst_dmem_n16078, MEM_stage_inst_dmem_n16077, MEM_stage_inst_dmem_n16076, MEM_stage_inst_dmem_n16075, MEM_stage_inst_dmem_n16074, MEM_stage_inst_dmem_n16073, MEM_stage_inst_dmem_n16072, MEM_stage_inst_dmem_n16071, MEM_stage_inst_dmem_n16070, MEM_stage_inst_dmem_n16069, MEM_stage_inst_dmem_n16068, MEM_stage_inst_dmem_n16067, MEM_stage_inst_dmem_n16066, MEM_stage_inst_dmem_n16065, MEM_stage_inst_dmem_n16064, MEM_stage_inst_dmem_n16063, MEM_stage_inst_dmem_n16062, MEM_stage_inst_dmem_n16061, MEM_stage_inst_dmem_n16060, MEM_stage_inst_dmem_n16059, MEM_stage_inst_dmem_n16058, MEM_stage_inst_dmem_n16057, MEM_stage_inst_dmem_n16056, MEM_stage_inst_dmem_n16055, MEM_stage_inst_dmem_n16054, MEM_stage_inst_dmem_n16053, MEM_stage_inst_dmem_n16052, MEM_stage_inst_dmem_n16051, MEM_stage_inst_dmem_n16050, MEM_stage_inst_dmem_n16049, MEM_stage_inst_dmem_n16048, MEM_stage_inst_dmem_n16047, MEM_stage_inst_dmem_n16046, MEM_stage_inst_dmem_n16045, MEM_stage_inst_dmem_n16044, MEM_stage_inst_dmem_n16043, MEM_stage_inst_dmem_n16042, MEM_stage_inst_dmem_n16041, MEM_stage_inst_dmem_n16040, MEM_stage_inst_dmem_n16039, MEM_stage_inst_dmem_n16038, MEM_stage_inst_dmem_n16037, MEM_stage_inst_dmem_n16036, MEM_stage_inst_dmem_n16035, MEM_stage_inst_dmem_n16034, MEM_stage_inst_dmem_n16033, MEM_stage_inst_dmem_n16032, MEM_stage_inst_dmem_n16031, MEM_stage_inst_dmem_n16030, MEM_stage_inst_dmem_n16029, MEM_stage_inst_dmem_n16028, MEM_stage_inst_dmem_n16027, MEM_stage_inst_dmem_n16026, MEM_stage_inst_dmem_n16025, MEM_stage_inst_dmem_n16024, MEM_stage_inst_dmem_n16023, MEM_stage_inst_dmem_n16022, MEM_stage_inst_dmem_n16021, MEM_stage_inst_dmem_n16020, MEM_stage_inst_dmem_n16019, MEM_stage_inst_dmem_n16018, MEM_stage_inst_dmem_n16017, MEM_stage_inst_dmem_n16016, MEM_stage_inst_dmem_n16015, MEM_stage_inst_dmem_n16014, MEM_stage_inst_dmem_n16013, MEM_stage_inst_dmem_n16012, MEM_stage_inst_dmem_n16011, MEM_stage_inst_dmem_n16010, MEM_stage_inst_dmem_n16009, MEM_stage_inst_dmem_n16008, MEM_stage_inst_dmem_n16007, MEM_stage_inst_dmem_n16006, MEM_stage_inst_dmem_n16005, MEM_stage_inst_dmem_n16004, MEM_stage_inst_dmem_n16003, MEM_stage_inst_dmem_n16002, MEM_stage_inst_dmem_n16001, MEM_stage_inst_dmem_n16000, MEM_stage_inst_dmem_n15999, MEM_stage_inst_dmem_n15998, MEM_stage_inst_dmem_n15997, MEM_stage_inst_dmem_n15996, MEM_stage_inst_dmem_n15995, MEM_stage_inst_dmem_n15994, MEM_stage_inst_dmem_n15993, MEM_stage_inst_dmem_n15992, MEM_stage_inst_dmem_n15991, MEM_stage_inst_dmem_n15990, MEM_stage_inst_dmem_n15989, MEM_stage_inst_dmem_n15988, MEM_stage_inst_dmem_n15987, MEM_stage_inst_dmem_n15986, MEM_stage_inst_dmem_n15985, MEM_stage_inst_dmem_n15984, MEM_stage_inst_dmem_n15983, MEM_stage_inst_dmem_n15982, MEM_stage_inst_dmem_n15981, MEM_stage_inst_dmem_n15980, MEM_stage_inst_dmem_n15979, MEM_stage_inst_dmem_n15978, MEM_stage_inst_dmem_n15977, MEM_stage_inst_dmem_n15976, MEM_stage_inst_dmem_n15975, MEM_stage_inst_dmem_n15974, MEM_stage_inst_dmem_n15973, MEM_stage_inst_dmem_n15972, MEM_stage_inst_dmem_n15971, MEM_stage_inst_dmem_n15970, MEM_stage_inst_dmem_n15969, MEM_stage_inst_dmem_n15968, MEM_stage_inst_dmem_n15967, MEM_stage_inst_dmem_n15966, MEM_stage_inst_dmem_n15965, MEM_stage_inst_dmem_n15964, MEM_stage_inst_dmem_n15963, MEM_stage_inst_dmem_n15962, MEM_stage_inst_dmem_n15961, MEM_stage_inst_dmem_n15960, MEM_stage_inst_dmem_n15959, MEM_stage_inst_dmem_n15958, MEM_stage_inst_dmem_n15957, MEM_stage_inst_dmem_n15956, MEM_stage_inst_dmem_n15955, MEM_stage_inst_dmem_n15954, MEM_stage_inst_dmem_n15953, MEM_stage_inst_dmem_n15952, MEM_stage_inst_dmem_n15951, MEM_stage_inst_dmem_n15950, MEM_stage_inst_dmem_n15949, MEM_stage_inst_dmem_n15948, MEM_stage_inst_dmem_n15947, MEM_stage_inst_dmem_n15946, MEM_stage_inst_dmem_n15945, MEM_stage_inst_dmem_n15944, MEM_stage_inst_dmem_n15943, MEM_stage_inst_dmem_n15942, MEM_stage_inst_dmem_n15941, MEM_stage_inst_dmem_n15940, MEM_stage_inst_dmem_n15939, MEM_stage_inst_dmem_n15938, MEM_stage_inst_dmem_n15937, MEM_stage_inst_dmem_n15936, MEM_stage_inst_dmem_n15935, MEM_stage_inst_dmem_n15934, MEM_stage_inst_dmem_n15933, MEM_stage_inst_dmem_n15932, MEM_stage_inst_dmem_n15931, MEM_stage_inst_dmem_n15930, MEM_stage_inst_dmem_n15929, MEM_stage_inst_dmem_n15928, MEM_stage_inst_dmem_n15927, MEM_stage_inst_dmem_n15926, MEM_stage_inst_dmem_n15925, MEM_stage_inst_dmem_n15924, MEM_stage_inst_dmem_n15923, MEM_stage_inst_dmem_n15922, MEM_stage_inst_dmem_n15921, MEM_stage_inst_dmem_n15920, MEM_stage_inst_dmem_n15919, MEM_stage_inst_dmem_n15918, MEM_stage_inst_dmem_n15917, MEM_stage_inst_dmem_n15916, MEM_stage_inst_dmem_n15915, MEM_stage_inst_dmem_n15914, MEM_stage_inst_dmem_n15913, MEM_stage_inst_dmem_n15912, MEM_stage_inst_dmem_n15911, MEM_stage_inst_dmem_n15910, MEM_stage_inst_dmem_n15909, MEM_stage_inst_dmem_n15908, MEM_stage_inst_dmem_n15907, MEM_stage_inst_dmem_n15906, MEM_stage_inst_dmem_n15905, MEM_stage_inst_dmem_n15904, MEM_stage_inst_dmem_n15903, MEM_stage_inst_dmem_n15902, MEM_stage_inst_dmem_n15901, MEM_stage_inst_dmem_n15900, MEM_stage_inst_dmem_n15899, MEM_stage_inst_dmem_n15898, MEM_stage_inst_dmem_n15897, MEM_stage_inst_dmem_n15896, MEM_stage_inst_dmem_n15895, MEM_stage_inst_dmem_n15894, MEM_stage_inst_dmem_n15893, MEM_stage_inst_dmem_n15892, MEM_stage_inst_dmem_n15891, MEM_stage_inst_dmem_n15890, MEM_stage_inst_dmem_n15889, MEM_stage_inst_dmem_n15888, MEM_stage_inst_dmem_n15887, MEM_stage_inst_dmem_n15886, MEM_stage_inst_dmem_n15885, MEM_stage_inst_dmem_n15884, MEM_stage_inst_dmem_n15883, MEM_stage_inst_dmem_n15882, MEM_stage_inst_dmem_n15881, MEM_stage_inst_dmem_n15880, MEM_stage_inst_dmem_n15879, MEM_stage_inst_dmem_n15878, MEM_stage_inst_dmem_n15877, MEM_stage_inst_dmem_n15876, MEM_stage_inst_dmem_n15875, MEM_stage_inst_dmem_n15874, MEM_stage_inst_dmem_n15873, MEM_stage_inst_dmem_n15872, MEM_stage_inst_dmem_n15871, MEM_stage_inst_dmem_n15870, MEM_stage_inst_dmem_n15869, MEM_stage_inst_dmem_n15868, MEM_stage_inst_dmem_n15867, MEM_stage_inst_dmem_n15866, MEM_stage_inst_dmem_n15865, MEM_stage_inst_dmem_n15864, MEM_stage_inst_dmem_n15863, MEM_stage_inst_dmem_n15862, MEM_stage_inst_dmem_n15861, MEM_stage_inst_dmem_n15860, MEM_stage_inst_dmem_n15859, MEM_stage_inst_dmem_n15858, MEM_stage_inst_dmem_n15857, MEM_stage_inst_dmem_n15856, MEM_stage_inst_dmem_n15855, MEM_stage_inst_dmem_n15854, MEM_stage_inst_dmem_n15853, MEM_stage_inst_dmem_n15852, MEM_stage_inst_dmem_n15851, MEM_stage_inst_dmem_n15850, MEM_stage_inst_dmem_n15849, MEM_stage_inst_dmem_n15848, MEM_stage_inst_dmem_n15847, MEM_stage_inst_dmem_n15846, MEM_stage_inst_dmem_n15845, MEM_stage_inst_dmem_n15844, MEM_stage_inst_dmem_n15843, MEM_stage_inst_dmem_n15842, MEM_stage_inst_dmem_n15841, MEM_stage_inst_dmem_n15840, MEM_stage_inst_dmem_n15839, MEM_stage_inst_dmem_n15838, MEM_stage_inst_dmem_n15837, MEM_stage_inst_dmem_n15836, MEM_stage_inst_dmem_n15835, MEM_stage_inst_dmem_n15834, MEM_stage_inst_dmem_n15833, MEM_stage_inst_dmem_n15832, MEM_stage_inst_dmem_n15831, MEM_stage_inst_dmem_n15830, MEM_stage_inst_dmem_n15829, MEM_stage_inst_dmem_n15828, MEM_stage_inst_dmem_n15827, MEM_stage_inst_dmem_n15826, MEM_stage_inst_dmem_n15825, MEM_stage_inst_dmem_n15824, MEM_stage_inst_dmem_n15823, MEM_stage_inst_dmem_n15822, MEM_stage_inst_dmem_n15821, MEM_stage_inst_dmem_n15820, MEM_stage_inst_dmem_n15819, MEM_stage_inst_dmem_n15818, MEM_stage_inst_dmem_n15817, MEM_stage_inst_dmem_n15816, MEM_stage_inst_dmem_n15815, MEM_stage_inst_dmem_n15814, MEM_stage_inst_dmem_n15813, MEM_stage_inst_dmem_n15812, MEM_stage_inst_dmem_n15811, MEM_stage_inst_dmem_n15810, MEM_stage_inst_dmem_n15809, MEM_stage_inst_dmem_n15808, MEM_stage_inst_dmem_n15807, MEM_stage_inst_dmem_n15806, MEM_stage_inst_dmem_n15805, MEM_stage_inst_dmem_n15804, MEM_stage_inst_dmem_n15803, MEM_stage_inst_dmem_n15802, MEM_stage_inst_dmem_n15801, MEM_stage_inst_dmem_n15800, MEM_stage_inst_dmem_n15799, MEM_stage_inst_dmem_n15798, MEM_stage_inst_dmem_n15797, MEM_stage_inst_dmem_n15796, MEM_stage_inst_dmem_n15795, MEM_stage_inst_dmem_n15794, MEM_stage_inst_dmem_n15793, MEM_stage_inst_dmem_n15792, MEM_stage_inst_dmem_n15791, MEM_stage_inst_dmem_n15790, MEM_stage_inst_dmem_n15789, MEM_stage_inst_dmem_n15788, MEM_stage_inst_dmem_n15787, MEM_stage_inst_dmem_n15786, MEM_stage_inst_dmem_n15785, MEM_stage_inst_dmem_n15784, MEM_stage_inst_dmem_n15783, MEM_stage_inst_dmem_n15782, MEM_stage_inst_dmem_n15781, MEM_stage_inst_dmem_n15780, MEM_stage_inst_dmem_n15779, MEM_stage_inst_dmem_n15778, MEM_stage_inst_dmem_n15777, MEM_stage_inst_dmem_n15776, MEM_stage_inst_dmem_n15775, MEM_stage_inst_dmem_n15774, MEM_stage_inst_dmem_n15773, MEM_stage_inst_dmem_n15772, MEM_stage_inst_dmem_n15771, MEM_stage_inst_dmem_n15770, MEM_stage_inst_dmem_n15769, MEM_stage_inst_dmem_n15768, MEM_stage_inst_dmem_n15767, MEM_stage_inst_dmem_n15766, MEM_stage_inst_dmem_n15765, MEM_stage_inst_dmem_n15764, MEM_stage_inst_dmem_n15763, MEM_stage_inst_dmem_n15762, MEM_stage_inst_dmem_n15761, MEM_stage_inst_dmem_n15760, MEM_stage_inst_dmem_n15759, MEM_stage_inst_dmem_n15758, MEM_stage_inst_dmem_n15757, MEM_stage_inst_dmem_n15756, MEM_stage_inst_dmem_n15755, MEM_stage_inst_dmem_n15754, MEM_stage_inst_dmem_n15753, MEM_stage_inst_dmem_n15752, MEM_stage_inst_dmem_n15751, MEM_stage_inst_dmem_n15750, MEM_stage_inst_dmem_n15749, MEM_stage_inst_dmem_n15748, MEM_stage_inst_dmem_n15747, MEM_stage_inst_dmem_n15746, MEM_stage_inst_dmem_n15745, MEM_stage_inst_dmem_n15744, MEM_stage_inst_dmem_n15743, MEM_stage_inst_dmem_n15742, MEM_stage_inst_dmem_n15741, MEM_stage_inst_dmem_n15740, MEM_stage_inst_dmem_n15739, MEM_stage_inst_dmem_n15738, MEM_stage_inst_dmem_n15737, MEM_stage_inst_dmem_n15736, MEM_stage_inst_dmem_n15735, MEM_stage_inst_dmem_n15734, MEM_stage_inst_dmem_n15733, MEM_stage_inst_dmem_n15732, MEM_stage_inst_dmem_n15731, MEM_stage_inst_dmem_n15730, MEM_stage_inst_dmem_n15729, MEM_stage_inst_dmem_n15728, MEM_stage_inst_dmem_n15727, MEM_stage_inst_dmem_n15726, MEM_stage_inst_dmem_n15725, MEM_stage_inst_dmem_n15724, MEM_stage_inst_dmem_n15723, MEM_stage_inst_dmem_n15722, MEM_stage_inst_dmem_n15721, MEM_stage_inst_dmem_n15720, MEM_stage_inst_dmem_n15719, MEM_stage_inst_dmem_n15718, MEM_stage_inst_dmem_n15717, MEM_stage_inst_dmem_n15716, MEM_stage_inst_dmem_n15715, MEM_stage_inst_dmem_n15714, MEM_stage_inst_dmem_n15713, MEM_stage_inst_dmem_n15712, MEM_stage_inst_dmem_n15711, MEM_stage_inst_dmem_n15710, MEM_stage_inst_dmem_n15709, MEM_stage_inst_dmem_n15708, MEM_stage_inst_dmem_n15707, MEM_stage_inst_dmem_n15706, MEM_stage_inst_dmem_n15705, MEM_stage_inst_dmem_n15704, MEM_stage_inst_dmem_n15703, MEM_stage_inst_dmem_n15702, MEM_stage_inst_dmem_n15701, MEM_stage_inst_dmem_n15700, MEM_stage_inst_dmem_n15699, MEM_stage_inst_dmem_n15698, MEM_stage_inst_dmem_n15697, MEM_stage_inst_dmem_n15696, MEM_stage_inst_dmem_n15695, MEM_stage_inst_dmem_n15694, MEM_stage_inst_dmem_n15693, MEM_stage_inst_dmem_n15692, MEM_stage_inst_dmem_n15691, MEM_stage_inst_dmem_n15690, MEM_stage_inst_dmem_n15689, MEM_stage_inst_dmem_n15688, MEM_stage_inst_dmem_n15687, MEM_stage_inst_dmem_n15686, MEM_stage_inst_dmem_n15685, MEM_stage_inst_dmem_n15684, MEM_stage_inst_dmem_n15683, MEM_stage_inst_dmem_n15682, MEM_stage_inst_dmem_n15681, MEM_stage_inst_dmem_n15680, MEM_stage_inst_dmem_n15679, MEM_stage_inst_dmem_n15678, MEM_stage_inst_dmem_n15677, MEM_stage_inst_dmem_n15676, MEM_stage_inst_dmem_n15675, MEM_stage_inst_dmem_n15674, MEM_stage_inst_dmem_n15673, MEM_stage_inst_dmem_n15672, MEM_stage_inst_dmem_n15671, MEM_stage_inst_dmem_n15670, MEM_stage_inst_dmem_n15669, MEM_stage_inst_dmem_n15668, MEM_stage_inst_dmem_n15667, MEM_stage_inst_dmem_n15666, MEM_stage_inst_dmem_n15665, MEM_stage_inst_dmem_n15664, MEM_stage_inst_dmem_n15663, MEM_stage_inst_dmem_n15662, MEM_stage_inst_dmem_n15661, MEM_stage_inst_dmem_n15660, MEM_stage_inst_dmem_n15659, MEM_stage_inst_dmem_n15658, MEM_stage_inst_dmem_n15657, MEM_stage_inst_dmem_n15656, MEM_stage_inst_dmem_n15655, MEM_stage_inst_dmem_n15654, MEM_stage_inst_dmem_n15653, MEM_stage_inst_dmem_n15652, MEM_stage_inst_dmem_n15651, MEM_stage_inst_dmem_n15650, MEM_stage_inst_dmem_n15649, MEM_stage_inst_dmem_n15648, MEM_stage_inst_dmem_n15647, MEM_stage_inst_dmem_n15646, MEM_stage_inst_dmem_n15645, MEM_stage_inst_dmem_n15644, MEM_stage_inst_dmem_n15643, MEM_stage_inst_dmem_n15642, MEM_stage_inst_dmem_n15641, MEM_stage_inst_dmem_n15640, MEM_stage_inst_dmem_n15639, MEM_stage_inst_dmem_n15638, MEM_stage_inst_dmem_n15637, MEM_stage_inst_dmem_n15636, MEM_stage_inst_dmem_n15635, MEM_stage_inst_dmem_n15634, MEM_stage_inst_dmem_n15633, MEM_stage_inst_dmem_n15632, MEM_stage_inst_dmem_n15631, MEM_stage_inst_dmem_n15630, MEM_stage_inst_dmem_n15629, MEM_stage_inst_dmem_n15628, MEM_stage_inst_dmem_n15627, MEM_stage_inst_dmem_n15626, MEM_stage_inst_dmem_n15625, MEM_stage_inst_dmem_n15624, MEM_stage_inst_dmem_n15623, MEM_stage_inst_dmem_n15622, MEM_stage_inst_dmem_n15621, MEM_stage_inst_dmem_n15620, MEM_stage_inst_dmem_n15619, MEM_stage_inst_dmem_n15618, MEM_stage_inst_dmem_n15617, MEM_stage_inst_dmem_n15616, MEM_stage_inst_dmem_n15615, MEM_stage_inst_dmem_n15614, MEM_stage_inst_dmem_n15613, MEM_stage_inst_dmem_n15612, MEM_stage_inst_dmem_n15611, MEM_stage_inst_dmem_n15610, MEM_stage_inst_dmem_n15609, MEM_stage_inst_dmem_n15608, MEM_stage_inst_dmem_n15607, MEM_stage_inst_dmem_n15606, MEM_stage_inst_dmem_n15605, MEM_stage_inst_dmem_n15604, MEM_stage_inst_dmem_n15603, MEM_stage_inst_dmem_n15602, MEM_stage_inst_dmem_n15601, MEM_stage_inst_dmem_n15600, MEM_stage_inst_dmem_n15599, MEM_stage_inst_dmem_n15598, MEM_stage_inst_dmem_n15597, MEM_stage_inst_dmem_n15596, MEM_stage_inst_dmem_n15595, MEM_stage_inst_dmem_n15594, MEM_stage_inst_dmem_n15593, MEM_stage_inst_dmem_n15592, MEM_stage_inst_dmem_n15591, MEM_stage_inst_dmem_n15590, MEM_stage_inst_dmem_n15589, MEM_stage_inst_dmem_n15588, MEM_stage_inst_dmem_n15587, MEM_stage_inst_dmem_n15586, MEM_stage_inst_dmem_n15585, MEM_stage_inst_dmem_n15584, MEM_stage_inst_dmem_n15583, MEM_stage_inst_dmem_n15582, MEM_stage_inst_dmem_n15581, MEM_stage_inst_dmem_n15580, MEM_stage_inst_dmem_n15579, MEM_stage_inst_dmem_n15578, MEM_stage_inst_dmem_n15577, MEM_stage_inst_dmem_n15576, MEM_stage_inst_dmem_n15575, MEM_stage_inst_dmem_n15574, MEM_stage_inst_dmem_n15573, MEM_stage_inst_dmem_n15572, MEM_stage_inst_dmem_n15571, MEM_stage_inst_dmem_n15570, MEM_stage_inst_dmem_n15569, MEM_stage_inst_dmem_n15568, MEM_stage_inst_dmem_n15567, MEM_stage_inst_dmem_n15566, MEM_stage_inst_dmem_n15565, MEM_stage_inst_dmem_n15564, MEM_stage_inst_dmem_n15563, MEM_stage_inst_dmem_n15562, MEM_stage_inst_dmem_n15561, MEM_stage_inst_dmem_n15560, MEM_stage_inst_dmem_n15559, MEM_stage_inst_dmem_n15558, MEM_stage_inst_dmem_n15557, MEM_stage_inst_dmem_n15556, MEM_stage_inst_dmem_n15555, MEM_stage_inst_dmem_n15554, MEM_stage_inst_dmem_n15553, MEM_stage_inst_dmem_n15552, MEM_stage_inst_dmem_n15551, MEM_stage_inst_dmem_n15550, MEM_stage_inst_dmem_n15549, MEM_stage_inst_dmem_n15548, MEM_stage_inst_dmem_n15547, MEM_stage_inst_dmem_n15546, MEM_stage_inst_dmem_n15545, MEM_stage_inst_dmem_n15544, MEM_stage_inst_dmem_n15543, MEM_stage_inst_dmem_n15542, MEM_stage_inst_dmem_n15541, MEM_stage_inst_dmem_n15540, MEM_stage_inst_dmem_n15539, MEM_stage_inst_dmem_n15538, MEM_stage_inst_dmem_n15537, MEM_stage_inst_dmem_n15536, MEM_stage_inst_dmem_n15535, MEM_stage_inst_dmem_n15534, MEM_stage_inst_dmem_n15533, MEM_stage_inst_dmem_n15532, MEM_stage_inst_dmem_n15531, MEM_stage_inst_dmem_n15530, MEM_stage_inst_dmem_n15529, MEM_stage_inst_dmem_n15528, MEM_stage_inst_dmem_n15527, MEM_stage_inst_dmem_n15526, MEM_stage_inst_dmem_n15525, MEM_stage_inst_dmem_n15524, MEM_stage_inst_dmem_n15523, MEM_stage_inst_dmem_n15522, MEM_stage_inst_dmem_n15521, MEM_stage_inst_dmem_n15520, MEM_stage_inst_dmem_n15519, MEM_stage_inst_dmem_n15518, MEM_stage_inst_dmem_n15517, MEM_stage_inst_dmem_n15516, MEM_stage_inst_dmem_n15515, MEM_stage_inst_dmem_n15514, MEM_stage_inst_dmem_n15513, MEM_stage_inst_dmem_n15512, MEM_stage_inst_dmem_n15511, MEM_stage_inst_dmem_n15510, MEM_stage_inst_dmem_n15509, MEM_stage_inst_dmem_n15508, MEM_stage_inst_dmem_n15507, MEM_stage_inst_dmem_n15506, MEM_stage_inst_dmem_n15505, MEM_stage_inst_dmem_n15504, MEM_stage_inst_dmem_n15503, MEM_stage_inst_dmem_n15502, MEM_stage_inst_dmem_n15501, MEM_stage_inst_dmem_n15500, MEM_stage_inst_dmem_n15499, MEM_stage_inst_dmem_n15498, MEM_stage_inst_dmem_n15497, MEM_stage_inst_dmem_n15496, MEM_stage_inst_dmem_n15495, MEM_stage_inst_dmem_n15494, MEM_stage_inst_dmem_n15493, MEM_stage_inst_dmem_n15492, MEM_stage_inst_dmem_n15491, MEM_stage_inst_dmem_n15490, MEM_stage_inst_dmem_n15489, MEM_stage_inst_dmem_n15488, MEM_stage_inst_dmem_n15487, MEM_stage_inst_dmem_n15486, MEM_stage_inst_dmem_n15485, MEM_stage_inst_dmem_n15484, MEM_stage_inst_dmem_n15483, MEM_stage_inst_dmem_n15482, MEM_stage_inst_dmem_n15481, MEM_stage_inst_dmem_n15480, MEM_stage_inst_dmem_n15479, MEM_stage_inst_dmem_n15478, MEM_stage_inst_dmem_n15477, MEM_stage_inst_dmem_n15476, MEM_stage_inst_dmem_n15475, MEM_stage_inst_dmem_n15474, MEM_stage_inst_dmem_n15473, MEM_stage_inst_dmem_n15472, MEM_stage_inst_dmem_n15471, MEM_stage_inst_dmem_n15470, MEM_stage_inst_dmem_n15469, MEM_stage_inst_dmem_n15468, MEM_stage_inst_dmem_n15467, MEM_stage_inst_dmem_n15466, MEM_stage_inst_dmem_n15465, MEM_stage_inst_dmem_n15464, MEM_stage_inst_dmem_n15463, MEM_stage_inst_dmem_n15462, MEM_stage_inst_dmem_n15461, MEM_stage_inst_dmem_n15460, MEM_stage_inst_dmem_n15459, MEM_stage_inst_dmem_n15458, MEM_stage_inst_dmem_n15457, MEM_stage_inst_dmem_n15456, MEM_stage_inst_dmem_n15455, MEM_stage_inst_dmem_n15454, MEM_stage_inst_dmem_n15453, MEM_stage_inst_dmem_n15452, MEM_stage_inst_dmem_n15451, MEM_stage_inst_dmem_n15450, MEM_stage_inst_dmem_n15449, MEM_stage_inst_dmem_n15448, MEM_stage_inst_dmem_n15447, MEM_stage_inst_dmem_n15446, MEM_stage_inst_dmem_n15445, MEM_stage_inst_dmem_n15444, MEM_stage_inst_dmem_n15443, MEM_stage_inst_dmem_n15442, MEM_stage_inst_dmem_n15441, MEM_stage_inst_dmem_n15440, MEM_stage_inst_dmem_n15439, MEM_stage_inst_dmem_n15438, MEM_stage_inst_dmem_n15437, MEM_stage_inst_dmem_n15436, MEM_stage_inst_dmem_n15435, MEM_stage_inst_dmem_n15434, MEM_stage_inst_dmem_n15433, MEM_stage_inst_dmem_n15432, MEM_stage_inst_dmem_n15431, MEM_stage_inst_dmem_n15430, MEM_stage_inst_dmem_n15429, MEM_stage_inst_dmem_n15428, MEM_stage_inst_dmem_n15427, MEM_stage_inst_dmem_n15426, MEM_stage_inst_dmem_n15425, MEM_stage_inst_dmem_n15424, MEM_stage_inst_dmem_n15423, MEM_stage_inst_dmem_n15422, MEM_stage_inst_dmem_n15421, MEM_stage_inst_dmem_n15420, MEM_stage_inst_dmem_n15419, MEM_stage_inst_dmem_n15418, MEM_stage_inst_dmem_n15417, MEM_stage_inst_dmem_n15416, MEM_stage_inst_dmem_n15415, MEM_stage_inst_dmem_n15414, MEM_stage_inst_dmem_n15413, MEM_stage_inst_dmem_n15412, MEM_stage_inst_dmem_n15411, MEM_stage_inst_dmem_n15410, MEM_stage_inst_dmem_n15409, MEM_stage_inst_dmem_n15408, MEM_stage_inst_dmem_n15407, MEM_stage_inst_dmem_n15406, MEM_stage_inst_dmem_n15405, MEM_stage_inst_dmem_n15404, MEM_stage_inst_dmem_n15403, MEM_stage_inst_dmem_n15402, MEM_stage_inst_dmem_n15401, MEM_stage_inst_dmem_n15400, MEM_stage_inst_dmem_n15399, MEM_stage_inst_dmem_n15398, MEM_stage_inst_dmem_n15397, MEM_stage_inst_dmem_n15396, MEM_stage_inst_dmem_n15395, MEM_stage_inst_dmem_n15394, MEM_stage_inst_dmem_n15393, MEM_stage_inst_dmem_n15392, MEM_stage_inst_dmem_n15391, MEM_stage_inst_dmem_n15390, MEM_stage_inst_dmem_n15389, MEM_stage_inst_dmem_n15388, MEM_stage_inst_dmem_n15387, MEM_stage_inst_dmem_n15386, MEM_stage_inst_dmem_n15385, MEM_stage_inst_dmem_n15384, MEM_stage_inst_dmem_n15383, MEM_stage_inst_dmem_n15382, MEM_stage_inst_dmem_n15381, MEM_stage_inst_dmem_n15380, MEM_stage_inst_dmem_n15379, MEM_stage_inst_dmem_n15378, MEM_stage_inst_dmem_n15377, MEM_stage_inst_dmem_n15376, MEM_stage_inst_dmem_n15375, MEM_stage_inst_dmem_n15374, MEM_stage_inst_dmem_n15373, MEM_stage_inst_dmem_n15372, MEM_stage_inst_dmem_n15371, MEM_stage_inst_dmem_n15370, MEM_stage_inst_dmem_n15369, MEM_stage_inst_dmem_n15368, MEM_stage_inst_dmem_n15367, MEM_stage_inst_dmem_n15366, MEM_stage_inst_dmem_n15365, MEM_stage_inst_dmem_n15364, MEM_stage_inst_dmem_n15363, MEM_stage_inst_dmem_n15362, MEM_stage_inst_dmem_n15361, MEM_stage_inst_dmem_n15360, MEM_stage_inst_dmem_n15359, MEM_stage_inst_dmem_n15358, MEM_stage_inst_dmem_n15357, MEM_stage_inst_dmem_n15356, MEM_stage_inst_dmem_n15355, MEM_stage_inst_dmem_n15354, MEM_stage_inst_dmem_n15353, MEM_stage_inst_dmem_n15352, MEM_stage_inst_dmem_n15351, MEM_stage_inst_dmem_n15350, MEM_stage_inst_dmem_n15349, MEM_stage_inst_dmem_n15348, MEM_stage_inst_dmem_n15347, MEM_stage_inst_dmem_n15346, MEM_stage_inst_dmem_n15345, MEM_stage_inst_dmem_n15344, MEM_stage_inst_dmem_n15343, MEM_stage_inst_dmem_n15342, MEM_stage_inst_dmem_n15341, MEM_stage_inst_dmem_n15340, MEM_stage_inst_dmem_n15339, MEM_stage_inst_dmem_n15338, MEM_stage_inst_dmem_n15337, MEM_stage_inst_dmem_n15336, MEM_stage_inst_dmem_n15335, MEM_stage_inst_dmem_n15334, MEM_stage_inst_dmem_n15333, MEM_stage_inst_dmem_n15332, MEM_stage_inst_dmem_n15331, MEM_stage_inst_dmem_n15330, MEM_stage_inst_dmem_n15329, MEM_stage_inst_dmem_n15328, MEM_stage_inst_dmem_n15327, MEM_stage_inst_dmem_n15326, MEM_stage_inst_dmem_n15325, MEM_stage_inst_dmem_n15324, MEM_stage_inst_dmem_n15323, MEM_stage_inst_dmem_n15322, MEM_stage_inst_dmem_n15321, MEM_stage_inst_dmem_n15320, MEM_stage_inst_dmem_n15319, MEM_stage_inst_dmem_n15318, MEM_stage_inst_dmem_n15317, MEM_stage_inst_dmem_n15316, MEM_stage_inst_dmem_n15315, MEM_stage_inst_dmem_n15314, MEM_stage_inst_dmem_n15313, MEM_stage_inst_dmem_n15312, MEM_stage_inst_dmem_n15311, MEM_stage_inst_dmem_n15310, MEM_stage_inst_dmem_n15309, MEM_stage_inst_dmem_n15308, MEM_stage_inst_dmem_n15307, MEM_stage_inst_dmem_n15306, MEM_stage_inst_dmem_n15305, MEM_stage_inst_dmem_n15304, MEM_stage_inst_dmem_n15303, MEM_stage_inst_dmem_n15302, MEM_stage_inst_dmem_n15301, MEM_stage_inst_dmem_n15300, MEM_stage_inst_dmem_n15299, MEM_stage_inst_dmem_n15298, MEM_stage_inst_dmem_n15297, MEM_stage_inst_dmem_n15296, MEM_stage_inst_dmem_n15295, MEM_stage_inst_dmem_n15294, MEM_stage_inst_dmem_n15293, MEM_stage_inst_dmem_n15292, MEM_stage_inst_dmem_n15291, MEM_stage_inst_dmem_n15290, MEM_stage_inst_dmem_n15289, MEM_stage_inst_dmem_n15288, MEM_stage_inst_dmem_n15287, MEM_stage_inst_dmem_n15286, MEM_stage_inst_dmem_n15285, MEM_stage_inst_dmem_n15284, MEM_stage_inst_dmem_n15283, MEM_stage_inst_dmem_n15282, MEM_stage_inst_dmem_n15281, MEM_stage_inst_dmem_n15280, MEM_stage_inst_dmem_n15279, MEM_stage_inst_dmem_n15278, MEM_stage_inst_dmem_n15277, MEM_stage_inst_dmem_n15276, MEM_stage_inst_dmem_n15275, MEM_stage_inst_dmem_n15274, MEM_stage_inst_dmem_n15273, MEM_stage_inst_dmem_n15272, MEM_stage_inst_dmem_n15271, MEM_stage_inst_dmem_n15270, MEM_stage_inst_dmem_n15269, MEM_stage_inst_dmem_n15268, MEM_stage_inst_dmem_n15267, MEM_stage_inst_dmem_n15266, MEM_stage_inst_dmem_n15265, MEM_stage_inst_dmem_n15264, MEM_stage_inst_dmem_n15263, MEM_stage_inst_dmem_n15262, MEM_stage_inst_dmem_n15261, MEM_stage_inst_dmem_n15260, MEM_stage_inst_dmem_n15259, MEM_stage_inst_dmem_n15258, MEM_stage_inst_dmem_n15257, MEM_stage_inst_dmem_n15256, MEM_stage_inst_dmem_n15255, MEM_stage_inst_dmem_n15254, MEM_stage_inst_dmem_n15253, MEM_stage_inst_dmem_n15252, MEM_stage_inst_dmem_n15251, MEM_stage_inst_dmem_n15250, MEM_stage_inst_dmem_n15249, MEM_stage_inst_dmem_n15248, MEM_stage_inst_dmem_n15247, MEM_stage_inst_dmem_n15246, MEM_stage_inst_dmem_n15245, MEM_stage_inst_dmem_n15244, MEM_stage_inst_dmem_n15243, MEM_stage_inst_dmem_n15242, MEM_stage_inst_dmem_n15241, MEM_stage_inst_dmem_n15240, MEM_stage_inst_dmem_n15239, MEM_stage_inst_dmem_n15238, MEM_stage_inst_dmem_n15237, MEM_stage_inst_dmem_n15236, MEM_stage_inst_dmem_n15235, MEM_stage_inst_dmem_n15234, MEM_stage_inst_dmem_n15233, MEM_stage_inst_dmem_n15232, MEM_stage_inst_dmem_n15231, MEM_stage_inst_dmem_n15230, MEM_stage_inst_dmem_n15229, MEM_stage_inst_dmem_n15228, MEM_stage_inst_dmem_n15227, MEM_stage_inst_dmem_n15226, MEM_stage_inst_dmem_n15225, MEM_stage_inst_dmem_n15224, MEM_stage_inst_dmem_n15223, MEM_stage_inst_dmem_n15222, MEM_stage_inst_dmem_n15221, MEM_stage_inst_dmem_n15220, MEM_stage_inst_dmem_n15219, MEM_stage_inst_dmem_n15218, MEM_stage_inst_dmem_n15217, MEM_stage_inst_dmem_n15216, MEM_stage_inst_dmem_n15215, MEM_stage_inst_dmem_n15214, MEM_stage_inst_dmem_n15213, MEM_stage_inst_dmem_n15212, MEM_stage_inst_dmem_n15211, MEM_stage_inst_dmem_n15210, MEM_stage_inst_dmem_n15209, MEM_stage_inst_dmem_n15208, MEM_stage_inst_dmem_n15207, MEM_stage_inst_dmem_n15206, MEM_stage_inst_dmem_n15205, MEM_stage_inst_dmem_n15204, MEM_stage_inst_dmem_n15203, MEM_stage_inst_dmem_n15202, MEM_stage_inst_dmem_n15201, MEM_stage_inst_dmem_n15200, MEM_stage_inst_dmem_n15199, MEM_stage_inst_dmem_n15198, MEM_stage_inst_dmem_n15197, MEM_stage_inst_dmem_n15196, MEM_stage_inst_dmem_n15195, MEM_stage_inst_dmem_n15194, MEM_stage_inst_dmem_n15193, MEM_stage_inst_dmem_n15192, MEM_stage_inst_dmem_n15191, MEM_stage_inst_dmem_n15190, MEM_stage_inst_dmem_n15189, MEM_stage_inst_dmem_n15188, MEM_stage_inst_dmem_n15187, MEM_stage_inst_dmem_n15186, MEM_stage_inst_dmem_n15185, MEM_stage_inst_dmem_n15184, MEM_stage_inst_dmem_n15183, MEM_stage_inst_dmem_n15182, MEM_stage_inst_dmem_n15181, MEM_stage_inst_dmem_n15180, MEM_stage_inst_dmem_n15179, MEM_stage_inst_dmem_n15178, MEM_stage_inst_dmem_n15177, MEM_stage_inst_dmem_n15176, MEM_stage_inst_dmem_n15175, MEM_stage_inst_dmem_n15174, MEM_stage_inst_dmem_n15173, MEM_stage_inst_dmem_n15172, MEM_stage_inst_dmem_n15171, MEM_stage_inst_dmem_n15170, MEM_stage_inst_dmem_n15169, MEM_stage_inst_dmem_n15168, MEM_stage_inst_dmem_n15167, MEM_stage_inst_dmem_n15166, MEM_stage_inst_dmem_n15165, MEM_stage_inst_dmem_n15164, MEM_stage_inst_dmem_n15163, MEM_stage_inst_dmem_n15162, MEM_stage_inst_dmem_n15161, MEM_stage_inst_dmem_n15160, MEM_stage_inst_dmem_n15159, MEM_stage_inst_dmem_n15158, MEM_stage_inst_dmem_n15157, MEM_stage_inst_dmem_n15156, MEM_stage_inst_dmem_n15155, MEM_stage_inst_dmem_n15154, MEM_stage_inst_dmem_n15153, MEM_stage_inst_dmem_n15152, MEM_stage_inst_dmem_n15151, MEM_stage_inst_dmem_n15150, MEM_stage_inst_dmem_n15149, MEM_stage_inst_dmem_n15148, MEM_stage_inst_dmem_n15147, MEM_stage_inst_dmem_n15146, MEM_stage_inst_dmem_n15145, MEM_stage_inst_dmem_n15144, MEM_stage_inst_dmem_n15143, MEM_stage_inst_dmem_n15142, MEM_stage_inst_dmem_n15141, MEM_stage_inst_dmem_n15140, MEM_stage_inst_dmem_n15139, MEM_stage_inst_dmem_n15138, MEM_stage_inst_dmem_n15137, MEM_stage_inst_dmem_n15136, MEM_stage_inst_dmem_n15135, MEM_stage_inst_dmem_n15134, MEM_stage_inst_dmem_n15133, MEM_stage_inst_dmem_n15132, MEM_stage_inst_dmem_n15131, MEM_stage_inst_dmem_n15130, MEM_stage_inst_dmem_n15129, MEM_stage_inst_dmem_n15128, MEM_stage_inst_dmem_n15127, MEM_stage_inst_dmem_n15126, MEM_stage_inst_dmem_n15125, MEM_stage_inst_dmem_n15124, MEM_stage_inst_dmem_n15123, MEM_stage_inst_dmem_n15122, MEM_stage_inst_dmem_n15121, MEM_stage_inst_dmem_n15120, MEM_stage_inst_dmem_n15119, MEM_stage_inst_dmem_n15118, MEM_stage_inst_dmem_n15117, MEM_stage_inst_dmem_n15116, MEM_stage_inst_dmem_n15115, MEM_stage_inst_dmem_n15114, MEM_stage_inst_dmem_n15113, MEM_stage_inst_dmem_n15112, MEM_stage_inst_dmem_n15111, MEM_stage_inst_dmem_n15110, MEM_stage_inst_dmem_n15109, MEM_stage_inst_dmem_n15108, MEM_stage_inst_dmem_n15107, MEM_stage_inst_dmem_n15106, MEM_stage_inst_dmem_n15105, MEM_stage_inst_dmem_n15104, MEM_stage_inst_dmem_n15103, MEM_stage_inst_dmem_n15102, MEM_stage_inst_dmem_n15101, MEM_stage_inst_dmem_n15100, MEM_stage_inst_dmem_n15099, MEM_stage_inst_dmem_n15098, MEM_stage_inst_dmem_n15097, MEM_stage_inst_dmem_n15096, MEM_stage_inst_dmem_n15095, MEM_stage_inst_dmem_n15094, MEM_stage_inst_dmem_n15093, MEM_stage_inst_dmem_n15092, MEM_stage_inst_dmem_n15091, MEM_stage_inst_dmem_n15090, MEM_stage_inst_dmem_n15089, MEM_stage_inst_dmem_n15088, MEM_stage_inst_dmem_n15087, MEM_stage_inst_dmem_n15086, MEM_stage_inst_dmem_n15085, MEM_stage_inst_dmem_n15084, MEM_stage_inst_dmem_n15083, MEM_stage_inst_dmem_n15082, MEM_stage_inst_dmem_n15081, MEM_stage_inst_dmem_n15080, MEM_stage_inst_dmem_n15079, MEM_stage_inst_dmem_n15078, MEM_stage_inst_dmem_n15077, MEM_stage_inst_dmem_n15076, MEM_stage_inst_dmem_n15075, MEM_stage_inst_dmem_n15074, MEM_stage_inst_dmem_n15073, MEM_stage_inst_dmem_n15072, MEM_stage_inst_dmem_n15071, MEM_stage_inst_dmem_n15070, MEM_stage_inst_dmem_n15069, MEM_stage_inst_dmem_n15068, MEM_stage_inst_dmem_n15067, MEM_stage_inst_dmem_n15066, MEM_stage_inst_dmem_n15065, MEM_stage_inst_dmem_n15064, MEM_stage_inst_dmem_n15063, MEM_stage_inst_dmem_n15062, MEM_stage_inst_dmem_n15061, MEM_stage_inst_dmem_n15060, MEM_stage_inst_dmem_n15059, MEM_stage_inst_dmem_n15058, MEM_stage_inst_dmem_n15057, MEM_stage_inst_dmem_n15056, MEM_stage_inst_dmem_n15055, MEM_stage_inst_dmem_n15054, MEM_stage_inst_dmem_n15053, MEM_stage_inst_dmem_n15052, MEM_stage_inst_dmem_n15051, MEM_stage_inst_dmem_n15050, MEM_stage_inst_dmem_n15049, MEM_stage_inst_dmem_n15048, MEM_stage_inst_dmem_n15047, MEM_stage_inst_dmem_n15046, MEM_stage_inst_dmem_n15045, MEM_stage_inst_dmem_n15044, MEM_stage_inst_dmem_n15043, MEM_stage_inst_dmem_n15042, MEM_stage_inst_dmem_n15041, MEM_stage_inst_dmem_n15040, MEM_stage_inst_dmem_n15039, MEM_stage_inst_dmem_n15038, MEM_stage_inst_dmem_n15037, MEM_stage_inst_dmem_n15036, MEM_stage_inst_dmem_n15035, MEM_stage_inst_dmem_n15034, MEM_stage_inst_dmem_n15033, MEM_stage_inst_dmem_n15032, MEM_stage_inst_dmem_n15031, MEM_stage_inst_dmem_n15030, MEM_stage_inst_dmem_n15029, MEM_stage_inst_dmem_n15028, MEM_stage_inst_dmem_n15027, MEM_stage_inst_dmem_n15026, MEM_stage_inst_dmem_n15025, MEM_stage_inst_dmem_n15024, MEM_stage_inst_dmem_n15023, MEM_stage_inst_dmem_n15022, MEM_stage_inst_dmem_n15021, MEM_stage_inst_dmem_n15020, MEM_stage_inst_dmem_n15019, MEM_stage_inst_dmem_n15018, MEM_stage_inst_dmem_n15017, MEM_stage_inst_dmem_n15016, MEM_stage_inst_dmem_n15015, MEM_stage_inst_dmem_n15014, MEM_stage_inst_dmem_n15013, MEM_stage_inst_dmem_n15012, MEM_stage_inst_dmem_n15011, MEM_stage_inst_dmem_n15010, MEM_stage_inst_dmem_n15009, MEM_stage_inst_dmem_n15008, MEM_stage_inst_dmem_n15007, MEM_stage_inst_dmem_n15006, MEM_stage_inst_dmem_n15005, MEM_stage_inst_dmem_n15004, MEM_stage_inst_dmem_n15003, MEM_stage_inst_dmem_n15002, MEM_stage_inst_dmem_n15001, MEM_stage_inst_dmem_n15000, MEM_stage_inst_dmem_n14999, MEM_stage_inst_dmem_n14998, MEM_stage_inst_dmem_n14997, MEM_stage_inst_dmem_n14996, MEM_stage_inst_dmem_n14995, MEM_stage_inst_dmem_n14994, MEM_stage_inst_dmem_n14993, MEM_stage_inst_dmem_n14992, MEM_stage_inst_dmem_n14991, MEM_stage_inst_dmem_n14990, MEM_stage_inst_dmem_n14989, MEM_stage_inst_dmem_n14988, MEM_stage_inst_dmem_n14987, MEM_stage_inst_dmem_n14986, MEM_stage_inst_dmem_n14985, MEM_stage_inst_dmem_n14984, MEM_stage_inst_dmem_n14983, MEM_stage_inst_dmem_n14982, MEM_stage_inst_dmem_n14981, MEM_stage_inst_dmem_n14980, MEM_stage_inst_dmem_n14979, MEM_stage_inst_dmem_n14978, MEM_stage_inst_dmem_n14977, MEM_stage_inst_dmem_n14976, MEM_stage_inst_dmem_n14975, MEM_stage_inst_dmem_n14974, MEM_stage_inst_dmem_n14973, MEM_stage_inst_dmem_n14972, MEM_stage_inst_dmem_n14971, MEM_stage_inst_dmem_n14970, MEM_stage_inst_dmem_n14969, MEM_stage_inst_dmem_n14968, MEM_stage_inst_dmem_n14967, MEM_stage_inst_dmem_n14966, MEM_stage_inst_dmem_n14965, MEM_stage_inst_dmem_n14964, MEM_stage_inst_dmem_n14963, MEM_stage_inst_dmem_n14962, MEM_stage_inst_dmem_n14961, MEM_stage_inst_dmem_n14960, MEM_stage_inst_dmem_n14959, MEM_stage_inst_dmem_n14958, MEM_stage_inst_dmem_n14957, MEM_stage_inst_dmem_n14956, MEM_stage_inst_dmem_n14955, MEM_stage_inst_dmem_n14954, MEM_stage_inst_dmem_n14953, MEM_stage_inst_dmem_n14952, MEM_stage_inst_dmem_n14951, MEM_stage_inst_dmem_n14950, MEM_stage_inst_dmem_n14949, MEM_stage_inst_dmem_n14948, MEM_stage_inst_dmem_n14947, MEM_stage_inst_dmem_n14946, MEM_stage_inst_dmem_n14945, MEM_stage_inst_dmem_n14944, MEM_stage_inst_dmem_n14943, MEM_stage_inst_dmem_n14942, MEM_stage_inst_dmem_n14941, MEM_stage_inst_dmem_n14940, MEM_stage_inst_dmem_n14939, MEM_stage_inst_dmem_n14938, MEM_stage_inst_dmem_n14937, MEM_stage_inst_dmem_n14936, MEM_stage_inst_dmem_n14935, MEM_stage_inst_dmem_n14934, MEM_stage_inst_dmem_n14933, MEM_stage_inst_dmem_n14932, MEM_stage_inst_dmem_n14931, MEM_stage_inst_dmem_n14930, MEM_stage_inst_dmem_n14929, MEM_stage_inst_dmem_n14928, MEM_stage_inst_dmem_n14927, MEM_stage_inst_dmem_n14926, MEM_stage_inst_dmem_n14925, MEM_stage_inst_dmem_n14924, MEM_stage_inst_dmem_n14923, MEM_stage_inst_dmem_n14922, MEM_stage_inst_dmem_n14921, MEM_stage_inst_dmem_n14920, MEM_stage_inst_dmem_n14919, MEM_stage_inst_dmem_n14918, MEM_stage_inst_dmem_n14917, MEM_stage_inst_dmem_n14916, MEM_stage_inst_dmem_n14915, MEM_stage_inst_dmem_n14914, MEM_stage_inst_dmem_n14913, MEM_stage_inst_dmem_n14912, MEM_stage_inst_dmem_n14911, MEM_stage_inst_dmem_n14910, MEM_stage_inst_dmem_n14909, MEM_stage_inst_dmem_n14908, MEM_stage_inst_dmem_n14907, MEM_stage_inst_dmem_n14906, MEM_stage_inst_dmem_n14905, MEM_stage_inst_dmem_n14904, MEM_stage_inst_dmem_n14903, MEM_stage_inst_dmem_n14902, MEM_stage_inst_dmem_n14901, MEM_stage_inst_dmem_n14900, MEM_stage_inst_dmem_n14899, MEM_stage_inst_dmem_n14898, MEM_stage_inst_dmem_n14897, MEM_stage_inst_dmem_n14896, MEM_stage_inst_dmem_n14895, MEM_stage_inst_dmem_n14894, MEM_stage_inst_dmem_n14893, MEM_stage_inst_dmem_n14892, MEM_stage_inst_dmem_n14891, MEM_stage_inst_dmem_n14890, MEM_stage_inst_dmem_n14889, MEM_stage_inst_dmem_n14888, MEM_stage_inst_dmem_n14887, MEM_stage_inst_dmem_n14886, MEM_stage_inst_dmem_n14885, MEM_stage_inst_dmem_n14884, MEM_stage_inst_dmem_n14883, MEM_stage_inst_dmem_n14882, MEM_stage_inst_dmem_n14881, MEM_stage_inst_dmem_n14880, MEM_stage_inst_dmem_n14879, MEM_stage_inst_dmem_n14878, MEM_stage_inst_dmem_n14877, MEM_stage_inst_dmem_n14876, MEM_stage_inst_dmem_n14875, MEM_stage_inst_dmem_n14874, MEM_stage_inst_dmem_n14873, MEM_stage_inst_dmem_n14872, MEM_stage_inst_dmem_n14871, MEM_stage_inst_dmem_n14870, MEM_stage_inst_dmem_n14869, MEM_stage_inst_dmem_n14868, MEM_stage_inst_dmem_n14867, MEM_stage_inst_dmem_n14866, MEM_stage_inst_dmem_n14865, MEM_stage_inst_dmem_n14864, MEM_stage_inst_dmem_n14863, MEM_stage_inst_dmem_n14862, MEM_stage_inst_dmem_n14861, MEM_stage_inst_dmem_n14860, MEM_stage_inst_dmem_n14859, MEM_stage_inst_dmem_n14858, MEM_stage_inst_dmem_n14857, MEM_stage_inst_dmem_n14856, MEM_stage_inst_dmem_n14855, MEM_stage_inst_dmem_n14854, MEM_stage_inst_dmem_n14853, MEM_stage_inst_dmem_n14852, MEM_stage_inst_dmem_n14851, MEM_stage_inst_dmem_n14850, MEM_stage_inst_dmem_n14849, MEM_stage_inst_dmem_n14848, MEM_stage_inst_dmem_n14847, MEM_stage_inst_dmem_n14846, MEM_stage_inst_dmem_n14845, MEM_stage_inst_dmem_n14844, MEM_stage_inst_dmem_n14843, MEM_stage_inst_dmem_n14842, MEM_stage_inst_dmem_n14841, MEM_stage_inst_dmem_n14840, MEM_stage_inst_dmem_n14839, MEM_stage_inst_dmem_n14838, MEM_stage_inst_dmem_n14837, MEM_stage_inst_dmem_n14836, MEM_stage_inst_dmem_n14835, MEM_stage_inst_dmem_n14834, MEM_stage_inst_dmem_n14833, MEM_stage_inst_dmem_n14832, MEM_stage_inst_dmem_n14831, MEM_stage_inst_dmem_n14830, MEM_stage_inst_dmem_n14829, MEM_stage_inst_dmem_n14828, MEM_stage_inst_dmem_n14827, MEM_stage_inst_dmem_n14826, MEM_stage_inst_dmem_n14825, MEM_stage_inst_dmem_n14824, MEM_stage_inst_dmem_n14823, MEM_stage_inst_dmem_n14822, MEM_stage_inst_dmem_n14821, MEM_stage_inst_dmem_n14820, MEM_stage_inst_dmem_n14819, MEM_stage_inst_dmem_n14818, MEM_stage_inst_dmem_n14817, MEM_stage_inst_dmem_n14816, MEM_stage_inst_dmem_n14815, MEM_stage_inst_dmem_n14814, MEM_stage_inst_dmem_n14813, MEM_stage_inst_dmem_n14812, MEM_stage_inst_dmem_n14811, MEM_stage_inst_dmem_n14810, MEM_stage_inst_dmem_n14809, MEM_stage_inst_dmem_n14808, MEM_stage_inst_dmem_n14807, MEM_stage_inst_dmem_n14806, MEM_stage_inst_dmem_n14805, MEM_stage_inst_dmem_n14804, MEM_stage_inst_dmem_n14803, MEM_stage_inst_dmem_n14802, MEM_stage_inst_dmem_n14801, MEM_stage_inst_dmem_n14800, MEM_stage_inst_dmem_n14799, MEM_stage_inst_dmem_n14798, MEM_stage_inst_dmem_n14797, MEM_stage_inst_dmem_n14796, MEM_stage_inst_dmem_n14795, MEM_stage_inst_dmem_n14794, MEM_stage_inst_dmem_n14793, MEM_stage_inst_dmem_n14792, MEM_stage_inst_dmem_n14791, MEM_stage_inst_dmem_n14790, MEM_stage_inst_dmem_n14789, MEM_stage_inst_dmem_n14788, MEM_stage_inst_dmem_n14787, MEM_stage_inst_dmem_n14786, MEM_stage_inst_dmem_n14785, MEM_stage_inst_dmem_n14784, MEM_stage_inst_dmem_n14783, MEM_stage_inst_dmem_n14782, MEM_stage_inst_dmem_n14781, MEM_stage_inst_dmem_n14780, MEM_stage_inst_dmem_n14779, MEM_stage_inst_dmem_n14778, MEM_stage_inst_dmem_n14777, MEM_stage_inst_dmem_n14776, MEM_stage_inst_dmem_n14775, MEM_stage_inst_dmem_n14774, MEM_stage_inst_dmem_n14773, MEM_stage_inst_dmem_n14772, MEM_stage_inst_dmem_n14771, MEM_stage_inst_dmem_n14770, MEM_stage_inst_dmem_n14769, MEM_stage_inst_dmem_n14768, MEM_stage_inst_dmem_n14767, MEM_stage_inst_dmem_n14766, MEM_stage_inst_dmem_n14765, MEM_stage_inst_dmem_n14764, MEM_stage_inst_dmem_n14763, MEM_stage_inst_dmem_n14762, MEM_stage_inst_dmem_n14761, MEM_stage_inst_dmem_n14760, MEM_stage_inst_dmem_n14759, MEM_stage_inst_dmem_n14758, MEM_stage_inst_dmem_n14757, MEM_stage_inst_dmem_n14756, MEM_stage_inst_dmem_n14755, MEM_stage_inst_dmem_n14754, MEM_stage_inst_dmem_n14753, MEM_stage_inst_dmem_n14752, MEM_stage_inst_dmem_n14751, MEM_stage_inst_dmem_n14750, MEM_stage_inst_dmem_n14749, MEM_stage_inst_dmem_n14748, MEM_stage_inst_dmem_n14747, MEM_stage_inst_dmem_n14746, MEM_stage_inst_dmem_n14745, MEM_stage_inst_dmem_n14744, MEM_stage_inst_dmem_n14743, MEM_stage_inst_dmem_n14742, MEM_stage_inst_dmem_n14741, MEM_stage_inst_dmem_n14740, MEM_stage_inst_dmem_n14739, MEM_stage_inst_dmem_n14738, MEM_stage_inst_dmem_n14737, MEM_stage_inst_dmem_n14736, MEM_stage_inst_dmem_n14735, MEM_stage_inst_dmem_n14734, MEM_stage_inst_dmem_n14733, MEM_stage_inst_dmem_n14732, MEM_stage_inst_dmem_n14731, MEM_stage_inst_dmem_n14730, MEM_stage_inst_dmem_n14729, MEM_stage_inst_dmem_n14728, MEM_stage_inst_dmem_n14727, MEM_stage_inst_dmem_n14726, MEM_stage_inst_dmem_n14725, MEM_stage_inst_dmem_n14724, MEM_stage_inst_dmem_n14723, MEM_stage_inst_dmem_n14722, MEM_stage_inst_dmem_n14721, MEM_stage_inst_dmem_n14720, MEM_stage_inst_dmem_n14719, MEM_stage_inst_dmem_n14718, MEM_stage_inst_dmem_n14717, MEM_stage_inst_dmem_n14716, MEM_stage_inst_dmem_n14715, MEM_stage_inst_dmem_n14713, MEM_stage_inst_dmem_n14712, MEM_stage_inst_dmem_n14711, MEM_stage_inst_dmem_n14710, MEM_stage_inst_dmem_n14709, MEM_stage_inst_dmem_n14708, MEM_stage_inst_dmem_n14707, MEM_stage_inst_dmem_n14706, MEM_stage_inst_dmem_n14705, MEM_stage_inst_dmem_n14704, MEM_stage_inst_dmem_n14703, MEM_stage_inst_dmem_n14702, MEM_stage_inst_dmem_n14701, MEM_stage_inst_dmem_n14700, MEM_stage_inst_dmem_n14698, MEM_stage_inst_dmem_n14697, MEM_stage_inst_dmem_n14696, MEM_stage_inst_dmem_n14695, MEM_stage_inst_dmem_n14694, MEM_stage_inst_dmem_n14693, MEM_stage_inst_dmem_n14692, MEM_stage_inst_dmem_n14691, MEM_stage_inst_dmem_n14690, MEM_stage_inst_dmem_n14689, MEM_stage_inst_dmem_n14688, MEM_stage_inst_dmem_n14687, MEM_stage_inst_dmem_n14686, MEM_stage_inst_dmem_n14685, MEM_stage_inst_dmem_n14684, MEM_stage_inst_dmem_n14683, MEM_stage_inst_dmem_n14682, MEM_stage_inst_dmem_n14681, MEM_stage_inst_dmem_n14680, MEM_stage_inst_dmem_n14679, MEM_stage_inst_dmem_n14678, MEM_stage_inst_dmem_n14677, MEM_stage_inst_dmem_n14676, MEM_stage_inst_dmem_n14675, MEM_stage_inst_dmem_n14674, MEM_stage_inst_dmem_n14673, MEM_stage_inst_dmem_n14672, MEM_stage_inst_dmem_n14671, MEM_stage_inst_dmem_n14670, MEM_stage_inst_dmem_n14669, MEM_stage_inst_dmem_n14668, MEM_stage_inst_dmem_n14667, MEM_stage_inst_dmem_n14666, MEM_stage_inst_dmem_n14665, MEM_stage_inst_dmem_n14664, MEM_stage_inst_dmem_n14663, MEM_stage_inst_dmem_n14662, MEM_stage_inst_dmem_n14661, MEM_stage_inst_dmem_n14660, MEM_stage_inst_dmem_n14659, MEM_stage_inst_dmem_n14658, MEM_stage_inst_dmem_n14657, MEM_stage_inst_dmem_n14656, MEM_stage_inst_dmem_n14655, MEM_stage_inst_dmem_n14654, MEM_stage_inst_dmem_n14653, MEM_stage_inst_dmem_n14652, MEM_stage_inst_dmem_n14651, MEM_stage_inst_dmem_n14650, MEM_stage_inst_dmem_n14649, MEM_stage_inst_dmem_n14648, MEM_stage_inst_dmem_n14647, MEM_stage_inst_dmem_n14646, MEM_stage_inst_dmem_n14645, MEM_stage_inst_dmem_n14644, MEM_stage_inst_dmem_n14643, MEM_stage_inst_dmem_n14642, MEM_stage_inst_dmem_n14641, MEM_stage_inst_dmem_n14640, MEM_stage_inst_dmem_n14639, MEM_stage_inst_dmem_n14638, MEM_stage_inst_dmem_n14637, MEM_stage_inst_dmem_n14636, MEM_stage_inst_dmem_n14635, MEM_stage_inst_dmem_n14634, MEM_stage_inst_dmem_n14633, MEM_stage_inst_dmem_n14632, MEM_stage_inst_dmem_n14631, MEM_stage_inst_dmem_n14630, MEM_stage_inst_dmem_n14629, MEM_stage_inst_dmem_n14628, MEM_stage_inst_dmem_n14627, MEM_stage_inst_dmem_n14626, MEM_stage_inst_dmem_n14625, MEM_stage_inst_dmem_n14624, MEM_stage_inst_dmem_n14623, MEM_stage_inst_dmem_n14622, MEM_stage_inst_dmem_n14621, MEM_stage_inst_dmem_n14620, MEM_stage_inst_dmem_n14619, MEM_stage_inst_dmem_n14618, MEM_stage_inst_dmem_n14617, MEM_stage_inst_dmem_n14616, MEM_stage_inst_dmem_n14615, MEM_stage_inst_dmem_n14614, MEM_stage_inst_dmem_n14613, MEM_stage_inst_dmem_n14612, MEM_stage_inst_dmem_n14611, MEM_stage_inst_dmem_n14610, MEM_stage_inst_dmem_n14609, MEM_stage_inst_dmem_n14608, MEM_stage_inst_dmem_n14607, MEM_stage_inst_dmem_n14606, MEM_stage_inst_dmem_n14605, MEM_stage_inst_dmem_n14604, MEM_stage_inst_dmem_n14603, MEM_stage_inst_dmem_n14602, MEM_stage_inst_dmem_n14601, MEM_stage_inst_dmem_n14600, MEM_stage_inst_dmem_n14599, MEM_stage_inst_dmem_n14598, MEM_stage_inst_dmem_n14597, MEM_stage_inst_dmem_n14596, MEM_stage_inst_dmem_n14595, MEM_stage_inst_dmem_n14594, MEM_stage_inst_dmem_n14593, MEM_stage_inst_dmem_n14592, MEM_stage_inst_dmem_n14591, MEM_stage_inst_dmem_n14590, MEM_stage_inst_dmem_n14589, MEM_stage_inst_dmem_n14588, MEM_stage_inst_dmem_n14587, MEM_stage_inst_dmem_n14586, MEM_stage_inst_dmem_n14585, MEM_stage_inst_dmem_n14584, MEM_stage_inst_dmem_n14583, MEM_stage_inst_dmem_n14582, MEM_stage_inst_dmem_n14581, MEM_stage_inst_dmem_n14580, MEM_stage_inst_dmem_n14579, MEM_stage_inst_dmem_n14578, MEM_stage_inst_dmem_n14577, MEM_stage_inst_dmem_n14576, MEM_stage_inst_dmem_n14575, MEM_stage_inst_dmem_n14574, MEM_stage_inst_dmem_n14573, MEM_stage_inst_dmem_n14572, MEM_stage_inst_dmem_n14571, MEM_stage_inst_dmem_n14570, MEM_stage_inst_dmem_n14569, MEM_stage_inst_dmem_n14568, MEM_stage_inst_dmem_n14567, MEM_stage_inst_dmem_n14566, MEM_stage_inst_dmem_n14565, MEM_stage_inst_dmem_n14564, MEM_stage_inst_dmem_n14563, MEM_stage_inst_dmem_n14562, MEM_stage_inst_dmem_n14561, MEM_stage_inst_dmem_n14560, MEM_stage_inst_dmem_n14559, MEM_stage_inst_dmem_n14558, MEM_stage_inst_dmem_n14557, MEM_stage_inst_dmem_n14556, MEM_stage_inst_dmem_n14555, MEM_stage_inst_dmem_n14554, MEM_stage_inst_dmem_n14553, MEM_stage_inst_dmem_n14552, MEM_stage_inst_dmem_n14551, MEM_stage_inst_dmem_n14550, MEM_stage_inst_dmem_n14549, MEM_stage_inst_dmem_n14548, MEM_stage_inst_dmem_n14547, MEM_stage_inst_dmem_n14546, MEM_stage_inst_dmem_n14545, MEM_stage_inst_dmem_n14544, MEM_stage_inst_dmem_n14543, MEM_stage_inst_dmem_n14542, MEM_stage_inst_dmem_n14541, MEM_stage_inst_dmem_n14540, MEM_stage_inst_dmem_n14539, MEM_stage_inst_dmem_n14538, MEM_stage_inst_dmem_n14537, MEM_stage_inst_dmem_n14536, MEM_stage_inst_dmem_n14535, MEM_stage_inst_dmem_n14534, MEM_stage_inst_dmem_n14533, MEM_stage_inst_dmem_n14532, MEM_stage_inst_dmem_n14531, MEM_stage_inst_dmem_n14530, MEM_stage_inst_dmem_n14529, MEM_stage_inst_dmem_n14528, MEM_stage_inst_dmem_n14527, MEM_stage_inst_dmem_n14526, MEM_stage_inst_dmem_n14525, MEM_stage_inst_dmem_n14524, MEM_stage_inst_dmem_n14523, MEM_stage_inst_dmem_n14522, MEM_stage_inst_dmem_n14521, MEM_stage_inst_dmem_n14520, MEM_stage_inst_dmem_n14519, MEM_stage_inst_dmem_n14518, MEM_stage_inst_dmem_n14517, MEM_stage_inst_dmem_n14516, MEM_stage_inst_dmem_n14515, MEM_stage_inst_dmem_n14514, MEM_stage_inst_dmem_n14513, MEM_stage_inst_dmem_n14512, MEM_stage_inst_dmem_n14511, MEM_stage_inst_dmem_n14510, MEM_stage_inst_dmem_n14509, MEM_stage_inst_dmem_n14508, MEM_stage_inst_dmem_n14507, MEM_stage_inst_dmem_n14506, MEM_stage_inst_dmem_n14505, MEM_stage_inst_dmem_n14504, MEM_stage_inst_dmem_n14503, MEM_stage_inst_dmem_n14502, MEM_stage_inst_dmem_n14501, MEM_stage_inst_dmem_n14500, MEM_stage_inst_dmem_n14499, MEM_stage_inst_dmem_n14498, MEM_stage_inst_dmem_n14497, MEM_stage_inst_dmem_n14496, MEM_stage_inst_dmem_n14495, MEM_stage_inst_dmem_n14494, MEM_stage_inst_dmem_n14493, MEM_stage_inst_dmem_n14492, MEM_stage_inst_dmem_n14491, MEM_stage_inst_dmem_n14490, MEM_stage_inst_dmem_n14489, MEM_stage_inst_dmem_n14488, MEM_stage_inst_dmem_n14487, MEM_stage_inst_dmem_n14486, MEM_stage_inst_dmem_n14485, MEM_stage_inst_dmem_n14484, MEM_stage_inst_dmem_n14483, MEM_stage_inst_dmem_n14482, MEM_stage_inst_dmem_n14481, MEM_stage_inst_dmem_n14480, MEM_stage_inst_dmem_n14479, MEM_stage_inst_dmem_n14478, MEM_stage_inst_dmem_n14477, MEM_stage_inst_dmem_n14476, MEM_stage_inst_dmem_n14475, MEM_stage_inst_dmem_n14474, MEM_stage_inst_dmem_n14473, MEM_stage_inst_dmem_n14472, MEM_stage_inst_dmem_n14471, MEM_stage_inst_dmem_n14470, MEM_stage_inst_dmem_n14469, MEM_stage_inst_dmem_n14468, MEM_stage_inst_dmem_n14467, MEM_stage_inst_dmem_n14466, MEM_stage_inst_dmem_n14465, MEM_stage_inst_dmem_n14464, MEM_stage_inst_dmem_n14463, MEM_stage_inst_dmem_n14462, MEM_stage_inst_dmem_n14461, MEM_stage_inst_dmem_n14460, MEM_stage_inst_dmem_n14459, MEM_stage_inst_dmem_n14458, MEM_stage_inst_dmem_n14457, MEM_stage_inst_dmem_n14456, MEM_stage_inst_dmem_n14455, MEM_stage_inst_dmem_n14454, MEM_stage_inst_dmem_n14453, MEM_stage_inst_dmem_n14452, MEM_stage_inst_dmem_n14451, MEM_stage_inst_dmem_n14450, MEM_stage_inst_dmem_n14449, MEM_stage_inst_dmem_n14448, MEM_stage_inst_dmem_n14447, MEM_stage_inst_dmem_n14446, MEM_stage_inst_dmem_n14445, MEM_stage_inst_dmem_n14444, MEM_stage_inst_dmem_n14443, MEM_stage_inst_dmem_n14442, MEM_stage_inst_dmem_n14441, MEM_stage_inst_dmem_n14440, MEM_stage_inst_dmem_n14439, MEM_stage_inst_dmem_n14438, MEM_stage_inst_dmem_n14437, MEM_stage_inst_dmem_n14436, MEM_stage_inst_dmem_n14435, MEM_stage_inst_dmem_n14434, MEM_stage_inst_dmem_n14433, MEM_stage_inst_dmem_n14432, MEM_stage_inst_dmem_n14431, MEM_stage_inst_dmem_n14430, MEM_stage_inst_dmem_n14429, MEM_stage_inst_dmem_n14428, MEM_stage_inst_dmem_n14427, MEM_stage_inst_dmem_n14426, MEM_stage_inst_dmem_n14425, MEM_stage_inst_dmem_n14424, MEM_stage_inst_dmem_n14423, MEM_stage_inst_dmem_n14422, MEM_stage_inst_dmem_n14421, MEM_stage_inst_dmem_n14420, MEM_stage_inst_dmem_n14419, MEM_stage_inst_dmem_n14418, MEM_stage_inst_dmem_n14417, MEM_stage_inst_dmem_n14416, MEM_stage_inst_dmem_n14415, MEM_stage_inst_dmem_n14414, MEM_stage_inst_dmem_n14413, MEM_stage_inst_dmem_n14412, MEM_stage_inst_dmem_n14411, MEM_stage_inst_dmem_n14410, MEM_stage_inst_dmem_n14409, MEM_stage_inst_dmem_n14408, MEM_stage_inst_dmem_n14407, MEM_stage_inst_dmem_n14406, MEM_stage_inst_dmem_n14405, MEM_stage_inst_dmem_n14404, MEM_stage_inst_dmem_n14403, MEM_stage_inst_dmem_n14402, MEM_stage_inst_dmem_n14401, MEM_stage_inst_dmem_n14400, MEM_stage_inst_dmem_n14399, MEM_stage_inst_dmem_n14398, MEM_stage_inst_dmem_n14397, MEM_stage_inst_dmem_n14396, MEM_stage_inst_dmem_n14395, MEM_stage_inst_dmem_n14394, MEM_stage_inst_dmem_n14393, MEM_stage_inst_dmem_n14392, MEM_stage_inst_dmem_n14391, MEM_stage_inst_dmem_n14390, MEM_stage_inst_dmem_n14389, MEM_stage_inst_dmem_n14388, MEM_stage_inst_dmem_n14387, MEM_stage_inst_dmem_n14386, MEM_stage_inst_dmem_n14385, MEM_stage_inst_dmem_n14384, MEM_stage_inst_dmem_n14383, MEM_stage_inst_dmem_n14382, MEM_stage_inst_dmem_n14381, MEM_stage_inst_dmem_n14380, MEM_stage_inst_dmem_n14379, MEM_stage_inst_dmem_n14378, MEM_stage_inst_dmem_n14377, MEM_stage_inst_dmem_n14376, MEM_stage_inst_dmem_n14375, MEM_stage_inst_dmem_n14374, MEM_stage_inst_dmem_n14373, MEM_stage_inst_dmem_n14372, MEM_stage_inst_dmem_n14371, MEM_stage_inst_dmem_n14370, MEM_stage_inst_dmem_n14369, MEM_stage_inst_dmem_n14368, MEM_stage_inst_dmem_n14367, MEM_stage_inst_dmem_n14366, MEM_stage_inst_dmem_n14365, MEM_stage_inst_dmem_n14364, MEM_stage_inst_dmem_n14363, MEM_stage_inst_dmem_n14362, MEM_stage_inst_dmem_n14361, MEM_stage_inst_dmem_n14360, MEM_stage_inst_dmem_n14359, MEM_stage_inst_dmem_n14358, MEM_stage_inst_dmem_n14357, MEM_stage_inst_dmem_n14356, MEM_stage_inst_dmem_n14355, MEM_stage_inst_dmem_n14354, MEM_stage_inst_dmem_n14353, MEM_stage_inst_dmem_n14352, MEM_stage_inst_dmem_n14351, MEM_stage_inst_dmem_n14350, MEM_stage_inst_dmem_n14349, MEM_stage_inst_dmem_n14348, MEM_stage_inst_dmem_n14347, MEM_stage_inst_dmem_n14346, MEM_stage_inst_dmem_n14345, MEM_stage_inst_dmem_n14344, MEM_stage_inst_dmem_n14343, MEM_stage_inst_dmem_n14342, MEM_stage_inst_dmem_n14341, MEM_stage_inst_dmem_n14340, MEM_stage_inst_dmem_n14339, MEM_stage_inst_dmem_n14338, MEM_stage_inst_dmem_n14337, MEM_stage_inst_dmem_n14336, MEM_stage_inst_dmem_n14335, MEM_stage_inst_dmem_n14334, MEM_stage_inst_dmem_n14333, MEM_stage_inst_dmem_n14332, MEM_stage_inst_dmem_n14331, MEM_stage_inst_dmem_n14330, MEM_stage_inst_dmem_n14329, MEM_stage_inst_dmem_n14328, MEM_stage_inst_dmem_n14327, MEM_stage_inst_dmem_n14326, MEM_stage_inst_dmem_n14325, MEM_stage_inst_dmem_n14324, MEM_stage_inst_dmem_n14323, MEM_stage_inst_dmem_n14322, MEM_stage_inst_dmem_n14321, MEM_stage_inst_dmem_n14320, MEM_stage_inst_dmem_n14319, MEM_stage_inst_dmem_n14318, MEM_stage_inst_dmem_n14317, MEM_stage_inst_dmem_n14316, MEM_stage_inst_dmem_n14315, MEM_stage_inst_dmem_n14314, MEM_stage_inst_dmem_n14313, MEM_stage_inst_dmem_n14312, MEM_stage_inst_dmem_n14311, MEM_stage_inst_dmem_n14310, MEM_stage_inst_dmem_n14309, MEM_stage_inst_dmem_n14308, MEM_stage_inst_dmem_n14307, MEM_stage_inst_dmem_n14306, MEM_stage_inst_dmem_n14305, MEM_stage_inst_dmem_n14304, MEM_stage_inst_dmem_n14303, MEM_stage_inst_dmem_n14302, MEM_stage_inst_dmem_n14301, MEM_stage_inst_dmem_n14300, MEM_stage_inst_dmem_n14299, MEM_stage_inst_dmem_n14298, MEM_stage_inst_dmem_n14297, MEM_stage_inst_dmem_n14296, MEM_stage_inst_dmem_n14295, MEM_stage_inst_dmem_n14294, MEM_stage_inst_dmem_n14293, MEM_stage_inst_dmem_n14292, MEM_stage_inst_dmem_n14291, MEM_stage_inst_dmem_n14290, MEM_stage_inst_dmem_n14289, MEM_stage_inst_dmem_n14288, MEM_stage_inst_dmem_n14287, MEM_stage_inst_dmem_n14286, MEM_stage_inst_dmem_n14285, MEM_stage_inst_dmem_n14284, MEM_stage_inst_dmem_n14283, MEM_stage_inst_dmem_n14282, MEM_stage_inst_dmem_n14281, MEM_stage_inst_dmem_n14280, MEM_stage_inst_dmem_n14279, MEM_stage_inst_dmem_n14278, MEM_stage_inst_dmem_n14277, MEM_stage_inst_dmem_n14276, MEM_stage_inst_dmem_n14275, MEM_stage_inst_dmem_n14274, MEM_stage_inst_dmem_n14273, MEM_stage_inst_dmem_n14272, MEM_stage_inst_dmem_n14271, MEM_stage_inst_dmem_n14270, MEM_stage_inst_dmem_n14269, MEM_stage_inst_dmem_n14268, MEM_stage_inst_dmem_n14267, MEM_stage_inst_dmem_n14266, MEM_stage_inst_dmem_n14265, MEM_stage_inst_dmem_n14264, MEM_stage_inst_dmem_n14263, MEM_stage_inst_dmem_n14262, MEM_stage_inst_dmem_n14261, MEM_stage_inst_dmem_n14260, MEM_stage_inst_dmem_n14259, MEM_stage_inst_dmem_n14258, MEM_stage_inst_dmem_n14257, MEM_stage_inst_dmem_n14256, MEM_stage_inst_dmem_n14255, MEM_stage_inst_dmem_n14254, MEM_stage_inst_dmem_n14253, MEM_stage_inst_dmem_n14252, MEM_stage_inst_dmem_n14251, MEM_stage_inst_dmem_n14250, MEM_stage_inst_dmem_n14249, MEM_stage_inst_dmem_n14248, MEM_stage_inst_dmem_n14247, MEM_stage_inst_dmem_n14246, MEM_stage_inst_dmem_n14245, MEM_stage_inst_dmem_n14244, MEM_stage_inst_dmem_n14243, MEM_stage_inst_dmem_n14242, MEM_stage_inst_dmem_n14241, MEM_stage_inst_dmem_n14240, MEM_stage_inst_dmem_n14239, MEM_stage_inst_dmem_n14238, MEM_stage_inst_dmem_n14237, MEM_stage_inst_dmem_n14236, MEM_stage_inst_dmem_n14235, MEM_stage_inst_dmem_n14234, MEM_stage_inst_dmem_n14233, MEM_stage_inst_dmem_n14232, MEM_stage_inst_dmem_n14231, MEM_stage_inst_dmem_n14230, MEM_stage_inst_dmem_n14229, MEM_stage_inst_dmem_n14228, MEM_stage_inst_dmem_n14227, MEM_stage_inst_dmem_n14226, MEM_stage_inst_dmem_n14225, MEM_stage_inst_dmem_n14224, MEM_stage_inst_dmem_n14223, MEM_stage_inst_dmem_n14222, MEM_stage_inst_dmem_n14221, MEM_stage_inst_dmem_n14220, MEM_stage_inst_dmem_n14219, MEM_stage_inst_dmem_n14218, MEM_stage_inst_dmem_n14217, MEM_stage_inst_dmem_n14216, MEM_stage_inst_dmem_n14215, MEM_stage_inst_dmem_n14214, MEM_stage_inst_dmem_n14213, MEM_stage_inst_dmem_n14212, MEM_stage_inst_dmem_n14211, MEM_stage_inst_dmem_n14210, MEM_stage_inst_dmem_n14209, MEM_stage_inst_dmem_n14208, MEM_stage_inst_dmem_n14207, MEM_stage_inst_dmem_n14206, MEM_stage_inst_dmem_n14205, MEM_stage_inst_dmem_n14204, MEM_stage_inst_dmem_n14203, MEM_stage_inst_dmem_n14202, MEM_stage_inst_dmem_n14201, MEM_stage_inst_dmem_n14200, MEM_stage_inst_dmem_n14199, MEM_stage_inst_dmem_n14198, MEM_stage_inst_dmem_n14197, MEM_stage_inst_dmem_n14196, MEM_stage_inst_dmem_n14195, MEM_stage_inst_dmem_n14194, MEM_stage_inst_dmem_n14193, MEM_stage_inst_dmem_n14192, MEM_stage_inst_dmem_n14191, MEM_stage_inst_dmem_n14190, MEM_stage_inst_dmem_n14189, MEM_stage_inst_dmem_n14188, MEM_stage_inst_dmem_n14187, MEM_stage_inst_dmem_n14186, MEM_stage_inst_dmem_n14185, MEM_stage_inst_dmem_n14184, MEM_stage_inst_dmem_n14183, MEM_stage_inst_dmem_n14182, MEM_stage_inst_dmem_n14181, MEM_stage_inst_dmem_n14180, MEM_stage_inst_dmem_n14179, MEM_stage_inst_dmem_n14178, MEM_stage_inst_dmem_n14177, MEM_stage_inst_dmem_n14176, MEM_stage_inst_dmem_n14175, MEM_stage_inst_dmem_n14174, MEM_stage_inst_dmem_n14173, MEM_stage_inst_dmem_n14172, MEM_stage_inst_dmem_n14171, MEM_stage_inst_dmem_n14170, MEM_stage_inst_dmem_n14169, MEM_stage_inst_dmem_n14168, MEM_stage_inst_dmem_n14167, MEM_stage_inst_dmem_n14166, MEM_stage_inst_dmem_n14165, MEM_stage_inst_dmem_n14164, MEM_stage_inst_dmem_n14163, MEM_stage_inst_dmem_n14162, MEM_stage_inst_dmem_n14161, MEM_stage_inst_dmem_n14160, MEM_stage_inst_dmem_n14159, MEM_stage_inst_dmem_n14158, MEM_stage_inst_dmem_n14157, MEM_stage_inst_dmem_n14156, MEM_stage_inst_dmem_n14155, MEM_stage_inst_dmem_n14154, MEM_stage_inst_dmem_n14153, MEM_stage_inst_dmem_n14152, MEM_stage_inst_dmem_n14151, MEM_stage_inst_dmem_n14150, MEM_stage_inst_dmem_n14149, MEM_stage_inst_dmem_n14148, MEM_stage_inst_dmem_n14147, MEM_stage_inst_dmem_n14146, MEM_stage_inst_dmem_n14145, MEM_stage_inst_dmem_n14144, MEM_stage_inst_dmem_n14143, MEM_stage_inst_dmem_n14142, MEM_stage_inst_dmem_n14141, MEM_stage_inst_dmem_n14140, MEM_stage_inst_dmem_n14139, MEM_stage_inst_dmem_n14138, MEM_stage_inst_dmem_n14137, MEM_stage_inst_dmem_n14136, MEM_stage_inst_dmem_n14135, MEM_stage_inst_dmem_n14134, MEM_stage_inst_dmem_n14133, MEM_stage_inst_dmem_n14132, MEM_stage_inst_dmem_n14131, MEM_stage_inst_dmem_n14130, MEM_stage_inst_dmem_n14129, MEM_stage_inst_dmem_n14128, MEM_stage_inst_dmem_n14127, MEM_stage_inst_dmem_n14126, MEM_stage_inst_dmem_n14125, MEM_stage_inst_dmem_n14124, MEM_stage_inst_dmem_n14123, MEM_stage_inst_dmem_n14122, MEM_stage_inst_dmem_n14121, MEM_stage_inst_dmem_n14120, MEM_stage_inst_dmem_n14119, MEM_stage_inst_dmem_n14118, MEM_stage_inst_dmem_n14117, MEM_stage_inst_dmem_n14116, MEM_stage_inst_dmem_n14115, MEM_stage_inst_dmem_n14114, MEM_stage_inst_dmem_n14113, MEM_stage_inst_dmem_n14112, MEM_stage_inst_dmem_n14111, MEM_stage_inst_dmem_n14110, MEM_stage_inst_dmem_n14109, MEM_stage_inst_dmem_n14108, MEM_stage_inst_dmem_n14107, MEM_stage_inst_dmem_n14106, MEM_stage_inst_dmem_n14105, MEM_stage_inst_dmem_n14104, MEM_stage_inst_dmem_n14103, MEM_stage_inst_dmem_n14102, MEM_stage_inst_dmem_n14101, MEM_stage_inst_dmem_n14100, MEM_stage_inst_dmem_n14099, MEM_stage_inst_dmem_n14098, MEM_stage_inst_dmem_n14097, MEM_stage_inst_dmem_n14096, MEM_stage_inst_dmem_n14095, MEM_stage_inst_dmem_n14094, MEM_stage_inst_dmem_n14093, MEM_stage_inst_dmem_n14092, MEM_stage_inst_dmem_n14091, MEM_stage_inst_dmem_n14090, MEM_stage_inst_dmem_n14089, MEM_stage_inst_dmem_n14088, MEM_stage_inst_dmem_n14087, MEM_stage_inst_dmem_n14086, MEM_stage_inst_dmem_n14085, MEM_stage_inst_dmem_n14084, MEM_stage_inst_dmem_n14083, MEM_stage_inst_dmem_n14082, MEM_stage_inst_dmem_n14081, MEM_stage_inst_dmem_n14080, MEM_stage_inst_dmem_n14079, MEM_stage_inst_dmem_n14078, MEM_stage_inst_dmem_n14077, MEM_stage_inst_dmem_n14076, MEM_stage_inst_dmem_n14075, MEM_stage_inst_dmem_n14074, MEM_stage_inst_dmem_n14073, MEM_stage_inst_dmem_n14072, MEM_stage_inst_dmem_n14071, MEM_stage_inst_dmem_n14070, MEM_stage_inst_dmem_n14069, MEM_stage_inst_dmem_n14068, MEM_stage_inst_dmem_n14067, MEM_stage_inst_dmem_n14066, MEM_stage_inst_dmem_n14065, MEM_stage_inst_dmem_n14064, MEM_stage_inst_dmem_n14063, MEM_stage_inst_dmem_n14062, MEM_stage_inst_dmem_n14061, MEM_stage_inst_dmem_n14060, MEM_stage_inst_dmem_n14059, MEM_stage_inst_dmem_n14058, MEM_stage_inst_dmem_n14057, MEM_stage_inst_dmem_n14056, MEM_stage_inst_dmem_n14055, MEM_stage_inst_dmem_n14054, MEM_stage_inst_dmem_n14053, MEM_stage_inst_dmem_n14052, MEM_stage_inst_dmem_n14051, MEM_stage_inst_dmem_n14050, MEM_stage_inst_dmem_n14049, MEM_stage_inst_dmem_n14048, MEM_stage_inst_dmem_n14047, MEM_stage_inst_dmem_n14046, MEM_stage_inst_dmem_n14045, MEM_stage_inst_dmem_n14044, MEM_stage_inst_dmem_n14043, MEM_stage_inst_dmem_n14042, MEM_stage_inst_dmem_n14041, MEM_stage_inst_dmem_n14040, MEM_stage_inst_dmem_n14039, MEM_stage_inst_dmem_n14038, MEM_stage_inst_dmem_n14037, MEM_stage_inst_dmem_n14036, MEM_stage_inst_dmem_n14035, MEM_stage_inst_dmem_n14034, MEM_stage_inst_dmem_n14033, MEM_stage_inst_dmem_n14032, MEM_stage_inst_dmem_n14031, MEM_stage_inst_dmem_n14030, MEM_stage_inst_dmem_n14029, MEM_stage_inst_dmem_n14028, MEM_stage_inst_dmem_n14027, MEM_stage_inst_dmem_n14026, MEM_stage_inst_dmem_n14025, MEM_stage_inst_dmem_n14024, MEM_stage_inst_dmem_n14023, MEM_stage_inst_dmem_n14022, MEM_stage_inst_dmem_n14021, MEM_stage_inst_dmem_n14020, MEM_stage_inst_dmem_n14019, MEM_stage_inst_dmem_n14018, MEM_stage_inst_dmem_n14017, MEM_stage_inst_dmem_n14016, MEM_stage_inst_dmem_n14015, MEM_stage_inst_dmem_n14014, MEM_stage_inst_dmem_n14013, MEM_stage_inst_dmem_n14012, MEM_stage_inst_dmem_n14011, MEM_stage_inst_dmem_n14010, MEM_stage_inst_dmem_n14009, MEM_stage_inst_dmem_n14008, MEM_stage_inst_dmem_n14007, MEM_stage_inst_dmem_n14006, MEM_stage_inst_dmem_n14005, MEM_stage_inst_dmem_n14004, MEM_stage_inst_dmem_n14003, MEM_stage_inst_dmem_n14002, MEM_stage_inst_dmem_n14001, MEM_stage_inst_dmem_n14000, MEM_stage_inst_dmem_n13999, MEM_stage_inst_dmem_n13998, MEM_stage_inst_dmem_n13997, MEM_stage_inst_dmem_n13996, MEM_stage_inst_dmem_n13995, MEM_stage_inst_dmem_n13994, MEM_stage_inst_dmem_n13993, MEM_stage_inst_dmem_n13992, MEM_stage_inst_dmem_n13991, MEM_stage_inst_dmem_n13990, MEM_stage_inst_dmem_n13989, MEM_stage_inst_dmem_n13988, MEM_stage_inst_dmem_n13987, MEM_stage_inst_dmem_n13986, MEM_stage_inst_dmem_n13985, MEM_stage_inst_dmem_n13984, MEM_stage_inst_dmem_n13983, MEM_stage_inst_dmem_n13982, MEM_stage_inst_dmem_n13981, MEM_stage_inst_dmem_n13980, MEM_stage_inst_dmem_n13979, MEM_stage_inst_dmem_n13978, MEM_stage_inst_dmem_n13977, MEM_stage_inst_dmem_n13976, MEM_stage_inst_dmem_n13975, MEM_stage_inst_dmem_n13974, MEM_stage_inst_dmem_n13973, MEM_stage_inst_dmem_n13972, MEM_stage_inst_dmem_n13971, MEM_stage_inst_dmem_n13970, MEM_stage_inst_dmem_n13969, MEM_stage_inst_dmem_n13968, MEM_stage_inst_dmem_n13967, MEM_stage_inst_dmem_n13966, MEM_stage_inst_dmem_n13965, MEM_stage_inst_dmem_n13964, MEM_stage_inst_dmem_n13963, MEM_stage_inst_dmem_n13962, MEM_stage_inst_dmem_n13961, MEM_stage_inst_dmem_n13960, MEM_stage_inst_dmem_n13959, MEM_stage_inst_dmem_n13958, MEM_stage_inst_dmem_n13957, MEM_stage_inst_dmem_n13956, MEM_stage_inst_dmem_n13955, MEM_stage_inst_dmem_n13954, MEM_stage_inst_dmem_n13953, MEM_stage_inst_dmem_n13952, MEM_stage_inst_dmem_n13951, MEM_stage_inst_dmem_n13950, MEM_stage_inst_dmem_n13949, MEM_stage_inst_dmem_n13948, MEM_stage_inst_dmem_n13947, MEM_stage_inst_dmem_n13946, MEM_stage_inst_dmem_n13945, MEM_stage_inst_dmem_n13944, MEM_stage_inst_dmem_n13943, MEM_stage_inst_dmem_n13942, MEM_stage_inst_dmem_n13941, MEM_stage_inst_dmem_n13940, MEM_stage_inst_dmem_n13939, MEM_stage_inst_dmem_n13938, MEM_stage_inst_dmem_n13937, MEM_stage_inst_dmem_n13936, MEM_stage_inst_dmem_n13935, MEM_stage_inst_dmem_n13934, MEM_stage_inst_dmem_n13933, MEM_stage_inst_dmem_n13932, MEM_stage_inst_dmem_n13931, MEM_stage_inst_dmem_n13930, MEM_stage_inst_dmem_n13929, MEM_stage_inst_dmem_n13928, MEM_stage_inst_dmem_n13927, MEM_stage_inst_dmem_n13926, MEM_stage_inst_dmem_n13925, MEM_stage_inst_dmem_n13924, MEM_stage_inst_dmem_n13923, MEM_stage_inst_dmem_n13922, MEM_stage_inst_dmem_n13921, MEM_stage_inst_dmem_n13920, MEM_stage_inst_dmem_n13919, MEM_stage_inst_dmem_n13918, MEM_stage_inst_dmem_n13917, MEM_stage_inst_dmem_n13916, MEM_stage_inst_dmem_n13915, MEM_stage_inst_dmem_n13914, MEM_stage_inst_dmem_n13913, MEM_stage_inst_dmem_n13912, MEM_stage_inst_dmem_n13911, MEM_stage_inst_dmem_n13910, MEM_stage_inst_dmem_n13909, MEM_stage_inst_dmem_n13908, MEM_stage_inst_dmem_n13907, MEM_stage_inst_dmem_n13906, MEM_stage_inst_dmem_n13905, MEM_stage_inst_dmem_n13904, MEM_stage_inst_dmem_n13902, MEM_stage_inst_dmem_n13901, MEM_stage_inst_dmem_n13900, MEM_stage_inst_dmem_n13899, MEM_stage_inst_dmem_n13898, MEM_stage_inst_dmem_n13897, MEM_stage_inst_dmem_n13896, MEM_stage_inst_dmem_n13895, MEM_stage_inst_dmem_n13894, MEM_stage_inst_dmem_n13893, MEM_stage_inst_dmem_n13892, MEM_stage_inst_dmem_n13891, MEM_stage_inst_dmem_n13890, MEM_stage_inst_dmem_n13889, MEM_stage_inst_dmem_n13888, MEM_stage_inst_dmem_n13887, MEM_stage_inst_dmem_n13886, MEM_stage_inst_dmem_n13885, MEM_stage_inst_dmem_n13884, MEM_stage_inst_dmem_n13883, MEM_stage_inst_dmem_n13882, MEM_stage_inst_dmem_n13881, MEM_stage_inst_dmem_n13880, MEM_stage_inst_dmem_n13879, MEM_stage_inst_dmem_n13878, MEM_stage_inst_dmem_n13877, MEM_stage_inst_dmem_n13876, MEM_stage_inst_dmem_n13875, MEM_stage_inst_dmem_n13874, MEM_stage_inst_dmem_n13873, MEM_stage_inst_dmem_n13872, MEM_stage_inst_dmem_n13871, MEM_stage_inst_dmem_n13870, MEM_stage_inst_dmem_n13869, MEM_stage_inst_dmem_n13868, MEM_stage_inst_dmem_n13867, MEM_stage_inst_dmem_n13866, MEM_stage_inst_dmem_n13865, MEM_stage_inst_dmem_n13864, MEM_stage_inst_dmem_n13863, MEM_stage_inst_dmem_n13862, MEM_stage_inst_dmem_n13861, MEM_stage_inst_dmem_n13860, MEM_stage_inst_dmem_n13859, MEM_stage_inst_dmem_n13858, MEM_stage_inst_dmem_n13857, MEM_stage_inst_dmem_n13856, MEM_stage_inst_dmem_n13855, MEM_stage_inst_dmem_n13854, MEM_stage_inst_dmem_n13853, MEM_stage_inst_dmem_n13852, MEM_stage_inst_dmem_n13851, MEM_stage_inst_dmem_n13850, MEM_stage_inst_dmem_n13849, MEM_stage_inst_dmem_n13848, MEM_stage_inst_dmem_n13847, MEM_stage_inst_dmem_n13846, MEM_stage_inst_dmem_n13845, MEM_stage_inst_dmem_n13844, MEM_stage_inst_dmem_n13843, MEM_stage_inst_dmem_n13842, MEM_stage_inst_dmem_n13841, MEM_stage_inst_dmem_n13840, MEM_stage_inst_dmem_n13839, MEM_stage_inst_dmem_n13838, MEM_stage_inst_dmem_n13837, MEM_stage_inst_dmem_n13836, MEM_stage_inst_dmem_n13835, MEM_stage_inst_dmem_n13834, MEM_stage_inst_dmem_n13833, MEM_stage_inst_dmem_n13832, MEM_stage_inst_dmem_n13831, MEM_stage_inst_dmem_n13830, MEM_stage_inst_dmem_n13829, MEM_stage_inst_dmem_n13828, MEM_stage_inst_dmem_n13827, MEM_stage_inst_dmem_n13826, MEM_stage_inst_dmem_n13825, MEM_stage_inst_dmem_n13824, MEM_stage_inst_dmem_n13823, MEM_stage_inst_dmem_n13822, MEM_stage_inst_dmem_n13821, MEM_stage_inst_dmem_n13820, MEM_stage_inst_dmem_n13819, MEM_stage_inst_dmem_n13818, MEM_stage_inst_dmem_n13817, MEM_stage_inst_dmem_n13816, MEM_stage_inst_dmem_n13815, MEM_stage_inst_dmem_n13814, MEM_stage_inst_dmem_n13813, MEM_stage_inst_dmem_n13812, MEM_stage_inst_dmem_n13811, MEM_stage_inst_dmem_n13810, MEM_stage_inst_dmem_n13809, MEM_stage_inst_dmem_n13808, MEM_stage_inst_dmem_n13807, MEM_stage_inst_dmem_n13806, MEM_stage_inst_dmem_n13805, MEM_stage_inst_dmem_n13804, MEM_stage_inst_dmem_n13803, MEM_stage_inst_dmem_n13802, MEM_stage_inst_dmem_n13801, MEM_stage_inst_dmem_n13800, MEM_stage_inst_dmem_n13799, MEM_stage_inst_dmem_n13798, MEM_stage_inst_dmem_n13797, MEM_stage_inst_dmem_n13796, MEM_stage_inst_dmem_n13795, MEM_stage_inst_dmem_n13794, MEM_stage_inst_dmem_n13793, MEM_stage_inst_dmem_n13792, MEM_stage_inst_dmem_n13791, MEM_stage_inst_dmem_n13790, MEM_stage_inst_dmem_n13789, MEM_stage_inst_dmem_n13788, MEM_stage_inst_dmem_n13787, MEM_stage_inst_dmem_n13786, MEM_stage_inst_dmem_n13785, MEM_stage_inst_dmem_n13784, MEM_stage_inst_dmem_n13783, MEM_stage_inst_dmem_n13782, MEM_stage_inst_dmem_n13781, MEM_stage_inst_dmem_n13780, MEM_stage_inst_dmem_n13779, MEM_stage_inst_dmem_n13778, MEM_stage_inst_dmem_n13777, MEM_stage_inst_dmem_n13776, MEM_stage_inst_dmem_n13775, MEM_stage_inst_dmem_n13774, MEM_stage_inst_dmem_n13773, MEM_stage_inst_dmem_n13772, MEM_stage_inst_dmem_n13771, MEM_stage_inst_dmem_n13770, MEM_stage_inst_dmem_n13769, MEM_stage_inst_dmem_n13768, MEM_stage_inst_dmem_n13767, MEM_stage_inst_dmem_n13766, MEM_stage_inst_dmem_n13765, MEM_stage_inst_dmem_n13764, MEM_stage_inst_dmem_n13763, MEM_stage_inst_dmem_n13762, MEM_stage_inst_dmem_n13761, MEM_stage_inst_dmem_n13760, MEM_stage_inst_dmem_n13759, MEM_stage_inst_dmem_n13758, MEM_stage_inst_dmem_n13757, MEM_stage_inst_dmem_n13756, MEM_stage_inst_dmem_n13755, MEM_stage_inst_dmem_n13754, MEM_stage_inst_dmem_n13753, MEM_stage_inst_dmem_n13752, MEM_stage_inst_dmem_n13751, MEM_stage_inst_dmem_n13750, MEM_stage_inst_dmem_n13749, MEM_stage_inst_dmem_n13748, MEM_stage_inst_dmem_n13747, MEM_stage_inst_dmem_n13746, MEM_stage_inst_dmem_n13745, MEM_stage_inst_dmem_n13744, MEM_stage_inst_dmem_n13743, MEM_stage_inst_dmem_n13742, MEM_stage_inst_dmem_n13741, MEM_stage_inst_dmem_n13740, MEM_stage_inst_dmem_n13739, MEM_stage_inst_dmem_n13738, MEM_stage_inst_dmem_n13737, MEM_stage_inst_dmem_n13736, MEM_stage_inst_dmem_n13735, MEM_stage_inst_dmem_n13734, MEM_stage_inst_dmem_n13733, MEM_stage_inst_dmem_n13732, MEM_stage_inst_dmem_n13731, MEM_stage_inst_dmem_n13730, MEM_stage_inst_dmem_n13729, MEM_stage_inst_dmem_n13728, MEM_stage_inst_dmem_n13727, MEM_stage_inst_dmem_n13726, MEM_stage_inst_dmem_n13725, MEM_stage_inst_dmem_n13724, MEM_stage_inst_dmem_n13723, MEM_stage_inst_dmem_n13722, MEM_stage_inst_dmem_n13721, MEM_stage_inst_dmem_n13720, MEM_stage_inst_dmem_n13719, MEM_stage_inst_dmem_n13718, MEM_stage_inst_dmem_n13717, MEM_stage_inst_dmem_n13716, MEM_stage_inst_dmem_n13715, MEM_stage_inst_dmem_n13714, MEM_stage_inst_dmem_n13713, MEM_stage_inst_dmem_n13712, MEM_stage_inst_dmem_n13711, MEM_stage_inst_dmem_n13710, MEM_stage_inst_dmem_n13709, MEM_stage_inst_dmem_n13708, MEM_stage_inst_dmem_n13707, MEM_stage_inst_dmem_n13706, MEM_stage_inst_dmem_n13705, MEM_stage_inst_dmem_n13704, MEM_stage_inst_dmem_n13703, MEM_stage_inst_dmem_n13702, MEM_stage_inst_dmem_n13701, MEM_stage_inst_dmem_n13700, MEM_stage_inst_dmem_n13699, MEM_stage_inst_dmem_n13698, MEM_stage_inst_dmem_n13697, MEM_stage_inst_dmem_n13696, MEM_stage_inst_dmem_n13695, MEM_stage_inst_dmem_n13694, MEM_stage_inst_dmem_n13693, MEM_stage_inst_dmem_n13692, MEM_stage_inst_dmem_n13691, MEM_stage_inst_dmem_n13690, MEM_stage_inst_dmem_n13689, MEM_stage_inst_dmem_n13688, MEM_stage_inst_dmem_n13687, MEM_stage_inst_dmem_n13686, MEM_stage_inst_dmem_n13685, MEM_stage_inst_dmem_n13684, MEM_stage_inst_dmem_n13683, MEM_stage_inst_dmem_n13682, MEM_stage_inst_dmem_n13681, MEM_stage_inst_dmem_n13680, MEM_stage_inst_dmem_n13679, MEM_stage_inst_dmem_n13678, MEM_stage_inst_dmem_n13677, MEM_stage_inst_dmem_n13676, MEM_stage_inst_dmem_n13675, MEM_stage_inst_dmem_n13674, MEM_stage_inst_dmem_n13673, MEM_stage_inst_dmem_n13672, MEM_stage_inst_dmem_n13671, MEM_stage_inst_dmem_n13670, MEM_stage_inst_dmem_n13669, MEM_stage_inst_dmem_n13668, MEM_stage_inst_dmem_n13667, MEM_stage_inst_dmem_n13666, MEM_stage_inst_dmem_n13665, MEM_stage_inst_dmem_n13664, MEM_stage_inst_dmem_n13663, MEM_stage_inst_dmem_n13662, MEM_stage_inst_dmem_n13661, MEM_stage_inst_dmem_n13660, MEM_stage_inst_dmem_n13659, MEM_stage_inst_dmem_n13658, MEM_stage_inst_dmem_n13657, MEM_stage_inst_dmem_n13656, MEM_stage_inst_dmem_n13655, MEM_stage_inst_dmem_n13654, MEM_stage_inst_dmem_n13653, MEM_stage_inst_dmem_n13652, MEM_stage_inst_dmem_n13651, MEM_stage_inst_dmem_n13650, MEM_stage_inst_dmem_n13649, MEM_stage_inst_dmem_n13648, MEM_stage_inst_dmem_n13647, MEM_stage_inst_dmem_n13646, MEM_stage_inst_dmem_n13645, MEM_stage_inst_dmem_n13644, MEM_stage_inst_dmem_n13643, MEM_stage_inst_dmem_n13642, MEM_stage_inst_dmem_n13641, MEM_stage_inst_dmem_n13640, MEM_stage_inst_dmem_n13639, MEM_stage_inst_dmem_n13638, MEM_stage_inst_dmem_n13637, MEM_stage_inst_dmem_n13636, MEM_stage_inst_dmem_n13635, MEM_stage_inst_dmem_n13634, MEM_stage_inst_dmem_n13633, MEM_stage_inst_dmem_n13632, MEM_stage_inst_dmem_n13631, MEM_stage_inst_dmem_n13630, MEM_stage_inst_dmem_n13629, MEM_stage_inst_dmem_n13628, MEM_stage_inst_dmem_n13627, MEM_stage_inst_dmem_n13626, MEM_stage_inst_dmem_n13625, MEM_stage_inst_dmem_n13624, MEM_stage_inst_dmem_n13623, MEM_stage_inst_dmem_n13622, MEM_stage_inst_dmem_n13621, MEM_stage_inst_dmem_n13620, MEM_stage_inst_dmem_n13619, MEM_stage_inst_dmem_n13618, MEM_stage_inst_dmem_n13617, MEM_stage_inst_dmem_n13616, MEM_stage_inst_dmem_n13615, MEM_stage_inst_dmem_n13614, MEM_stage_inst_dmem_n13613, MEM_stage_inst_dmem_n13612, MEM_stage_inst_dmem_n13611, MEM_stage_inst_dmem_n13610, MEM_stage_inst_dmem_n13609, MEM_stage_inst_dmem_n13608, MEM_stage_inst_dmem_n13607, MEM_stage_inst_dmem_n13606, MEM_stage_inst_dmem_n13605, MEM_stage_inst_dmem_n13604, MEM_stage_inst_dmem_n13603, MEM_stage_inst_dmem_n13602, MEM_stage_inst_dmem_n13601, MEM_stage_inst_dmem_n13600, MEM_stage_inst_dmem_n13599, MEM_stage_inst_dmem_n13598, MEM_stage_inst_dmem_n13597, MEM_stage_inst_dmem_n13596, MEM_stage_inst_dmem_n13595, MEM_stage_inst_dmem_n13594, MEM_stage_inst_dmem_n13593, MEM_stage_inst_dmem_n13592, MEM_stage_inst_dmem_n13591, MEM_stage_inst_dmem_n13590, MEM_stage_inst_dmem_n13589, MEM_stage_inst_dmem_n13588, MEM_stage_inst_dmem_n13587, MEM_stage_inst_dmem_n13586, MEM_stage_inst_dmem_n13585, MEM_stage_inst_dmem_n13584, MEM_stage_inst_dmem_n13583, MEM_stage_inst_dmem_n13582, MEM_stage_inst_dmem_n13581, MEM_stage_inst_dmem_n13580, MEM_stage_inst_dmem_n13579, MEM_stage_inst_dmem_n13578, MEM_stage_inst_dmem_n13577, MEM_stage_inst_dmem_n13576, MEM_stage_inst_dmem_n13575, MEM_stage_inst_dmem_n13574, MEM_stage_inst_dmem_n13573, MEM_stage_inst_dmem_n13572, MEM_stage_inst_dmem_n13571, MEM_stage_inst_dmem_n13570, MEM_stage_inst_dmem_n13569, MEM_stage_inst_dmem_n13568, MEM_stage_inst_dmem_n13567, MEM_stage_inst_dmem_n13566, MEM_stage_inst_dmem_n13565, MEM_stage_inst_dmem_n13564, MEM_stage_inst_dmem_n13563, MEM_stage_inst_dmem_n13562, MEM_stage_inst_dmem_n13561, MEM_stage_inst_dmem_n13560, MEM_stage_inst_dmem_n13559, MEM_stage_inst_dmem_n13558, MEM_stage_inst_dmem_n13557, MEM_stage_inst_dmem_n13556, MEM_stage_inst_dmem_n13555, MEM_stage_inst_dmem_n13554, MEM_stage_inst_dmem_n13553, MEM_stage_inst_dmem_n13552, MEM_stage_inst_dmem_n13551, MEM_stage_inst_dmem_n13550, MEM_stage_inst_dmem_n13549, MEM_stage_inst_dmem_n13548, MEM_stage_inst_dmem_n13547, MEM_stage_inst_dmem_n13546, MEM_stage_inst_dmem_n13545, MEM_stage_inst_dmem_n13544, MEM_stage_inst_dmem_n13543, MEM_stage_inst_dmem_n13542, MEM_stage_inst_dmem_n13541, MEM_stage_inst_dmem_n13540, MEM_stage_inst_dmem_n13539, MEM_stage_inst_dmem_n13538, MEM_stage_inst_dmem_n13537, MEM_stage_inst_dmem_n13536, MEM_stage_inst_dmem_n13535, MEM_stage_inst_dmem_n13534, MEM_stage_inst_dmem_n13533, MEM_stage_inst_dmem_n13532, MEM_stage_inst_dmem_n13531, MEM_stage_inst_dmem_n13530, MEM_stage_inst_dmem_n13529, MEM_stage_inst_dmem_n13528, MEM_stage_inst_dmem_n13527, MEM_stage_inst_dmem_n13526, MEM_stage_inst_dmem_n13525, MEM_stage_inst_dmem_n13524, MEM_stage_inst_dmem_n13523, MEM_stage_inst_dmem_n13522, MEM_stage_inst_dmem_n13521, MEM_stage_inst_dmem_n13520, MEM_stage_inst_dmem_n13519, MEM_stage_inst_dmem_n13518, MEM_stage_inst_dmem_n13517, MEM_stage_inst_dmem_n13516, MEM_stage_inst_dmem_n13515, MEM_stage_inst_dmem_n13514, MEM_stage_inst_dmem_n13513, MEM_stage_inst_dmem_n13512, MEM_stage_inst_dmem_n13511, MEM_stage_inst_dmem_n13510, MEM_stage_inst_dmem_n13509, MEM_stage_inst_dmem_n13508, MEM_stage_inst_dmem_n13507, MEM_stage_inst_dmem_n13506, MEM_stage_inst_dmem_n13505, MEM_stage_inst_dmem_n13504, MEM_stage_inst_dmem_n13503, MEM_stage_inst_dmem_n13502, MEM_stage_inst_dmem_n13501, MEM_stage_inst_dmem_n13500, MEM_stage_inst_dmem_n13499, MEM_stage_inst_dmem_n13498, MEM_stage_inst_dmem_n13497, MEM_stage_inst_dmem_n13496, MEM_stage_inst_dmem_n13495, MEM_stage_inst_dmem_n13494, MEM_stage_inst_dmem_n13493, MEM_stage_inst_dmem_n13492, MEM_stage_inst_dmem_n13491, MEM_stage_inst_dmem_n13490, MEM_stage_inst_dmem_n13489, MEM_stage_inst_dmem_n13488, MEM_stage_inst_dmem_n13487, MEM_stage_inst_dmem_n13486, MEM_stage_inst_dmem_n13485, MEM_stage_inst_dmem_n13484, MEM_stage_inst_dmem_n13483, MEM_stage_inst_dmem_n13482, MEM_stage_inst_dmem_n13481, MEM_stage_inst_dmem_n13480, MEM_stage_inst_dmem_n13479, MEM_stage_inst_dmem_n13478, MEM_stage_inst_dmem_n13477, MEM_stage_inst_dmem_n13476, MEM_stage_inst_dmem_n13475, MEM_stage_inst_dmem_n13474, MEM_stage_inst_dmem_n13473, MEM_stage_inst_dmem_n13472, MEM_stage_inst_dmem_n13471, MEM_stage_inst_dmem_n13470, MEM_stage_inst_dmem_n13469, MEM_stage_inst_dmem_n13468, MEM_stage_inst_dmem_n13467, MEM_stage_inst_dmem_n13466, MEM_stage_inst_dmem_n13465, MEM_stage_inst_dmem_n13464, MEM_stage_inst_dmem_n13463, MEM_stage_inst_dmem_n13462, MEM_stage_inst_dmem_n13461, MEM_stage_inst_dmem_n13460, MEM_stage_inst_dmem_n13459, MEM_stage_inst_dmem_n13458, MEM_stage_inst_dmem_n13457, MEM_stage_inst_dmem_n13456, MEM_stage_inst_dmem_n13455, MEM_stage_inst_dmem_n13454, MEM_stage_inst_dmem_n13453, MEM_stage_inst_dmem_n13452, MEM_stage_inst_dmem_n13451, MEM_stage_inst_dmem_n13450, MEM_stage_inst_dmem_n13449, MEM_stage_inst_dmem_n13448, MEM_stage_inst_dmem_n13447, MEM_stage_inst_dmem_n13446, MEM_stage_inst_dmem_n13445, MEM_stage_inst_dmem_n13444, MEM_stage_inst_dmem_n13443, MEM_stage_inst_dmem_n13442, MEM_stage_inst_dmem_n13441, MEM_stage_inst_dmem_n13440, MEM_stage_inst_dmem_n13439, MEM_stage_inst_dmem_n13438, MEM_stage_inst_dmem_n13437, MEM_stage_inst_dmem_n13436, MEM_stage_inst_dmem_n13435, MEM_stage_inst_dmem_n13434, MEM_stage_inst_dmem_n13433, MEM_stage_inst_dmem_n13432, MEM_stage_inst_dmem_n13431, MEM_stage_inst_dmem_n13430, MEM_stage_inst_dmem_n13429, MEM_stage_inst_dmem_n13428, MEM_stage_inst_dmem_n13427, MEM_stage_inst_dmem_n13426, MEM_stage_inst_dmem_n13425, MEM_stage_inst_dmem_n13424, MEM_stage_inst_dmem_n13423, MEM_stage_inst_dmem_n13422, MEM_stage_inst_dmem_n13421, MEM_stage_inst_dmem_n13420, MEM_stage_inst_dmem_n13419, MEM_stage_inst_dmem_n13418, MEM_stage_inst_dmem_n13417, MEM_stage_inst_dmem_n13416, MEM_stage_inst_dmem_n13415, MEM_stage_inst_dmem_n13414, MEM_stage_inst_dmem_n13413, MEM_stage_inst_dmem_n13412, MEM_stage_inst_dmem_n13411, MEM_stage_inst_dmem_n13410, MEM_stage_inst_dmem_n13409, MEM_stage_inst_dmem_n13408, MEM_stage_inst_dmem_n13407, MEM_stage_inst_dmem_n13406, MEM_stage_inst_dmem_n13405, MEM_stage_inst_dmem_n13404, MEM_stage_inst_dmem_n13403, MEM_stage_inst_dmem_n13402, MEM_stage_inst_dmem_n13401, MEM_stage_inst_dmem_n13400, MEM_stage_inst_dmem_n13399, MEM_stage_inst_dmem_n13398, MEM_stage_inst_dmem_n13397, MEM_stage_inst_dmem_n13396, MEM_stage_inst_dmem_n13395, MEM_stage_inst_dmem_n13394, MEM_stage_inst_dmem_n13393, MEM_stage_inst_dmem_n13392, MEM_stage_inst_dmem_n13391, MEM_stage_inst_dmem_n13390, MEM_stage_inst_dmem_n13389, MEM_stage_inst_dmem_n13388, MEM_stage_inst_dmem_n13387, MEM_stage_inst_dmem_n13386, MEM_stage_inst_dmem_n13385, MEM_stage_inst_dmem_n13384, MEM_stage_inst_dmem_n13383, MEM_stage_inst_dmem_n13382, MEM_stage_inst_dmem_n13381, MEM_stage_inst_dmem_n13380, MEM_stage_inst_dmem_n13379, MEM_stage_inst_dmem_n13378, MEM_stage_inst_dmem_n13377, MEM_stage_inst_dmem_n13376, MEM_stage_inst_dmem_n13375, MEM_stage_inst_dmem_n13374, MEM_stage_inst_dmem_n13373, MEM_stage_inst_dmem_n13372, MEM_stage_inst_dmem_n13371, MEM_stage_inst_dmem_n13370, MEM_stage_inst_dmem_n13369, MEM_stage_inst_dmem_n13368, MEM_stage_inst_dmem_n13367, MEM_stage_inst_dmem_n13366, MEM_stage_inst_dmem_n13365, MEM_stage_inst_dmem_n13364, MEM_stage_inst_dmem_n13363, MEM_stage_inst_dmem_n13362, MEM_stage_inst_dmem_n13361, MEM_stage_inst_dmem_n13360, MEM_stage_inst_dmem_n13359, MEM_stage_inst_dmem_n13358, MEM_stage_inst_dmem_n13357, MEM_stage_inst_dmem_n13356, MEM_stage_inst_dmem_n13355, MEM_stage_inst_dmem_n13354, MEM_stage_inst_dmem_n13353, MEM_stage_inst_dmem_n13352, MEM_stage_inst_dmem_n13351, MEM_stage_inst_dmem_n13350, MEM_stage_inst_dmem_n13349, MEM_stage_inst_dmem_n13348, MEM_stage_inst_dmem_n13347, MEM_stage_inst_dmem_n13346, MEM_stage_inst_dmem_n13345, MEM_stage_inst_dmem_n13344, MEM_stage_inst_dmem_n13343, MEM_stage_inst_dmem_n13342, MEM_stage_inst_dmem_n13341, MEM_stage_inst_dmem_n13340, MEM_stage_inst_dmem_n13339, MEM_stage_inst_dmem_n13338, MEM_stage_inst_dmem_n13337, MEM_stage_inst_dmem_n13336, MEM_stage_inst_dmem_n13335, MEM_stage_inst_dmem_n13334, MEM_stage_inst_dmem_n13333, MEM_stage_inst_dmem_n13332, MEM_stage_inst_dmem_n13331, MEM_stage_inst_dmem_n13330, MEM_stage_inst_dmem_n13329, MEM_stage_inst_dmem_n13328, MEM_stage_inst_dmem_n13327, MEM_stage_inst_dmem_n13326, MEM_stage_inst_dmem_n13325, MEM_stage_inst_dmem_n13324, MEM_stage_inst_dmem_n13323, MEM_stage_inst_dmem_n13322, MEM_stage_inst_dmem_n13321, MEM_stage_inst_dmem_n13320, MEM_stage_inst_dmem_n13319, MEM_stage_inst_dmem_n13318, MEM_stage_inst_dmem_n13317, MEM_stage_inst_dmem_n13316, MEM_stage_inst_dmem_n13315, MEM_stage_inst_dmem_n13314, MEM_stage_inst_dmem_n13313, MEM_stage_inst_dmem_n13312, MEM_stage_inst_dmem_n13311, MEM_stage_inst_dmem_n13310, MEM_stage_inst_dmem_n13309, MEM_stage_inst_dmem_n13308, MEM_stage_inst_dmem_n13307, MEM_stage_inst_dmem_n13306, MEM_stage_inst_dmem_n13305, MEM_stage_inst_dmem_n13304, MEM_stage_inst_dmem_n13303, MEM_stage_inst_dmem_n13302, MEM_stage_inst_dmem_n13301, MEM_stage_inst_dmem_n13300, MEM_stage_inst_dmem_n13299, MEM_stage_inst_dmem_n13298, MEM_stage_inst_dmem_n13297, MEM_stage_inst_dmem_n13296, MEM_stage_inst_dmem_n13295, MEM_stage_inst_dmem_n13294, MEM_stage_inst_dmem_n13293, MEM_stage_inst_dmem_n13292, MEM_stage_inst_dmem_n13291, MEM_stage_inst_dmem_n13290, MEM_stage_inst_dmem_n13289, MEM_stage_inst_dmem_n13288, MEM_stage_inst_dmem_n13287, MEM_stage_inst_dmem_n13286, MEM_stage_inst_dmem_n13285, MEM_stage_inst_dmem_n13284, MEM_stage_inst_dmem_n13283, MEM_stage_inst_dmem_n13282, MEM_stage_inst_dmem_n13281, MEM_stage_inst_dmem_n13280, MEM_stage_inst_dmem_n13279, MEM_stage_inst_dmem_n13278, MEM_stage_inst_dmem_n13277, MEM_stage_inst_dmem_n13276, MEM_stage_inst_dmem_n13275, MEM_stage_inst_dmem_n13274, MEM_stage_inst_dmem_n13273, MEM_stage_inst_dmem_n13272, MEM_stage_inst_dmem_n13271, MEM_stage_inst_dmem_n13270, MEM_stage_inst_dmem_n13269, MEM_stage_inst_dmem_n13268, MEM_stage_inst_dmem_n13267, MEM_stage_inst_dmem_n13266, MEM_stage_inst_dmem_n13265, MEM_stage_inst_dmem_n13264, MEM_stage_inst_dmem_n13263, MEM_stage_inst_dmem_n13262, MEM_stage_inst_dmem_n13261, MEM_stage_inst_dmem_n13260, MEM_stage_inst_dmem_n13259, MEM_stage_inst_dmem_n13258, MEM_stage_inst_dmem_n13257, MEM_stage_inst_dmem_n13256, MEM_stage_inst_dmem_n13255, MEM_stage_inst_dmem_n13254, MEM_stage_inst_dmem_n13253, MEM_stage_inst_dmem_n13252, MEM_stage_inst_dmem_n13251, MEM_stage_inst_dmem_n13250, MEM_stage_inst_dmem_n13249, MEM_stage_inst_dmem_n13248, MEM_stage_inst_dmem_n13247, MEM_stage_inst_dmem_n13246, MEM_stage_inst_dmem_n13245, MEM_stage_inst_dmem_n13244, MEM_stage_inst_dmem_n13243, MEM_stage_inst_dmem_n13242, MEM_stage_inst_dmem_n13241, MEM_stage_inst_dmem_n13240, MEM_stage_inst_dmem_n13239, MEM_stage_inst_dmem_n13238, MEM_stage_inst_dmem_n13237, MEM_stage_inst_dmem_n13236, MEM_stage_inst_dmem_n13235, MEM_stage_inst_dmem_n13234, MEM_stage_inst_dmem_n13233, MEM_stage_inst_dmem_n13232, MEM_stage_inst_dmem_n13231, MEM_stage_inst_dmem_n13230, MEM_stage_inst_dmem_n13229, MEM_stage_inst_dmem_n13228, MEM_stage_inst_dmem_n13227, MEM_stage_inst_dmem_n13226, MEM_stage_inst_dmem_n13225, MEM_stage_inst_dmem_n13224, MEM_stage_inst_dmem_n13223, MEM_stage_inst_dmem_n13222, MEM_stage_inst_dmem_n13221, MEM_stage_inst_dmem_n13220, MEM_stage_inst_dmem_n13219, MEM_stage_inst_dmem_n13218, MEM_stage_inst_dmem_n13217, MEM_stage_inst_dmem_n13216, MEM_stage_inst_dmem_n13215, MEM_stage_inst_dmem_n13214, MEM_stage_inst_dmem_n13213, MEM_stage_inst_dmem_n13212, MEM_stage_inst_dmem_n13211, MEM_stage_inst_dmem_n13210, MEM_stage_inst_dmem_n13209, MEM_stage_inst_dmem_n13208, MEM_stage_inst_dmem_n13207, MEM_stage_inst_dmem_n13206, MEM_stage_inst_dmem_n13205, MEM_stage_inst_dmem_n13204, MEM_stage_inst_dmem_n13203, MEM_stage_inst_dmem_n13202, MEM_stage_inst_dmem_n13201, MEM_stage_inst_dmem_n13200, MEM_stage_inst_dmem_n13199, MEM_stage_inst_dmem_n13198, MEM_stage_inst_dmem_n13197, MEM_stage_inst_dmem_n13196, MEM_stage_inst_dmem_n13195, MEM_stage_inst_dmem_n13194, MEM_stage_inst_dmem_n13193, MEM_stage_inst_dmem_n13192, MEM_stage_inst_dmem_n13191, MEM_stage_inst_dmem_n13190, MEM_stage_inst_dmem_n13189, MEM_stage_inst_dmem_n13188, MEM_stage_inst_dmem_n13187, MEM_stage_inst_dmem_n13186, MEM_stage_inst_dmem_n13185, MEM_stage_inst_dmem_n13184, MEM_stage_inst_dmem_n13183, MEM_stage_inst_dmem_n13182, MEM_stage_inst_dmem_n13181, MEM_stage_inst_dmem_n13180, MEM_stage_inst_dmem_n13179, MEM_stage_inst_dmem_n13178, MEM_stage_inst_dmem_n13177, MEM_stage_inst_dmem_n13176, MEM_stage_inst_dmem_n13175, MEM_stage_inst_dmem_n13174, MEM_stage_inst_dmem_n13173, MEM_stage_inst_dmem_n13172, MEM_stage_inst_dmem_n13171, MEM_stage_inst_dmem_n13170, MEM_stage_inst_dmem_n13169, MEM_stage_inst_dmem_n13168, MEM_stage_inst_dmem_n13167, MEM_stage_inst_dmem_n13166, MEM_stage_inst_dmem_n13165, MEM_stage_inst_dmem_n13164, MEM_stage_inst_dmem_n13163, MEM_stage_inst_dmem_n13162, MEM_stage_inst_dmem_n13161, MEM_stage_inst_dmem_n13160, MEM_stage_inst_dmem_n13159, MEM_stage_inst_dmem_n13158, MEM_stage_inst_dmem_n13157, MEM_stage_inst_dmem_n13156, MEM_stage_inst_dmem_n13155, MEM_stage_inst_dmem_n13154, MEM_stage_inst_dmem_n13153, MEM_stage_inst_dmem_n13152, MEM_stage_inst_dmem_n13151, MEM_stage_inst_dmem_n13150, MEM_stage_inst_dmem_n13149, MEM_stage_inst_dmem_n13148, MEM_stage_inst_dmem_n13147, MEM_stage_inst_dmem_n13146, MEM_stage_inst_dmem_n13145, MEM_stage_inst_dmem_n13144, MEM_stage_inst_dmem_n13143, MEM_stage_inst_dmem_n13142, MEM_stage_inst_dmem_n13141, MEM_stage_inst_dmem_n13140, MEM_stage_inst_dmem_n13139, MEM_stage_inst_dmem_n13138, MEM_stage_inst_dmem_n13137, MEM_stage_inst_dmem_n13136, MEM_stage_inst_dmem_n13135, MEM_stage_inst_dmem_n13134, MEM_stage_inst_dmem_n13133, MEM_stage_inst_dmem_n13132, MEM_stage_inst_dmem_n13131, MEM_stage_inst_dmem_n13130, MEM_stage_inst_dmem_n13129, MEM_stage_inst_dmem_n13128, MEM_stage_inst_dmem_n13127, MEM_stage_inst_dmem_n13126, MEM_stage_inst_dmem_n13125, MEM_stage_inst_dmem_n13124, MEM_stage_inst_dmem_n13123, MEM_stage_inst_dmem_n13122, MEM_stage_inst_dmem_n13121, MEM_stage_inst_dmem_n13120, MEM_stage_inst_dmem_n13119, MEM_stage_inst_dmem_n13118, MEM_stage_inst_dmem_n13117, MEM_stage_inst_dmem_n13116, MEM_stage_inst_dmem_n13115, MEM_stage_inst_dmem_n13114, MEM_stage_inst_dmem_n13113, MEM_stage_inst_dmem_n13112, MEM_stage_inst_dmem_n13111, MEM_stage_inst_dmem_n13110, MEM_stage_inst_dmem_n13109, MEM_stage_inst_dmem_n13108, MEM_stage_inst_dmem_n13107, MEM_stage_inst_dmem_n13106, MEM_stage_inst_dmem_n13105, MEM_stage_inst_dmem_n13104, MEM_stage_inst_dmem_n13103, MEM_stage_inst_dmem_n13102, MEM_stage_inst_dmem_n13101, MEM_stage_inst_dmem_n13100, MEM_stage_inst_dmem_n13099, MEM_stage_inst_dmem_n13098, MEM_stage_inst_dmem_n13097, MEM_stage_inst_dmem_n13096, MEM_stage_inst_dmem_n13095, MEM_stage_inst_dmem_n13094, MEM_stage_inst_dmem_n13093, MEM_stage_inst_dmem_n13092, MEM_stage_inst_dmem_n13091, MEM_stage_inst_dmem_n13090, MEM_stage_inst_dmem_n13089, MEM_stage_inst_dmem_n13088, MEM_stage_inst_dmem_n13087, MEM_stage_inst_dmem_n13086, MEM_stage_inst_dmem_n13085, MEM_stage_inst_dmem_n13084, MEM_stage_inst_dmem_n13083, MEM_stage_inst_dmem_n13082, MEM_stage_inst_dmem_n13081, MEM_stage_inst_dmem_n13080, MEM_stage_inst_dmem_n13079, MEM_stage_inst_dmem_n13078, MEM_stage_inst_dmem_n13077, MEM_stage_inst_dmem_n13076, MEM_stage_inst_dmem_n13075, MEM_stage_inst_dmem_n13074, MEM_stage_inst_dmem_n13073, MEM_stage_inst_dmem_n13072, MEM_stage_inst_dmem_n13071, MEM_stage_inst_dmem_n13070, MEM_stage_inst_dmem_n13068, MEM_stage_inst_dmem_n13067, MEM_stage_inst_dmem_n13066, MEM_stage_inst_dmem_n13065, MEM_stage_inst_dmem_n13064, MEM_stage_inst_dmem_n13063, MEM_stage_inst_dmem_n13062, MEM_stage_inst_dmem_n13061, MEM_stage_inst_dmem_n13060, MEM_stage_inst_dmem_n13059, MEM_stage_inst_dmem_n13058, MEM_stage_inst_dmem_n13057, MEM_stage_inst_dmem_n13056, MEM_stage_inst_dmem_n13055, MEM_stage_inst_dmem_n13054, MEM_stage_inst_dmem_n13053, MEM_stage_inst_dmem_n13052, MEM_stage_inst_dmem_n13051, MEM_stage_inst_dmem_n13050, MEM_stage_inst_dmem_n13049, MEM_stage_inst_dmem_n13048, MEM_stage_inst_dmem_n13047, MEM_stage_inst_dmem_n13046, MEM_stage_inst_dmem_n13045, MEM_stage_inst_dmem_n13044, MEM_stage_inst_dmem_n13043, MEM_stage_inst_dmem_n13042, MEM_stage_inst_dmem_n13041, MEM_stage_inst_dmem_n13040, MEM_stage_inst_dmem_n13039, MEM_stage_inst_dmem_n13038, MEM_stage_inst_dmem_n13037, MEM_stage_inst_dmem_n13036, MEM_stage_inst_dmem_n13035, MEM_stage_inst_dmem_n13034, MEM_stage_inst_dmem_n13033, MEM_stage_inst_dmem_n13032, MEM_stage_inst_dmem_n13031, MEM_stage_inst_dmem_n13030, MEM_stage_inst_dmem_n13029, MEM_stage_inst_dmem_n13028, MEM_stage_inst_dmem_n13027, MEM_stage_inst_dmem_n13026, MEM_stage_inst_dmem_n13025, MEM_stage_inst_dmem_n13024, MEM_stage_inst_dmem_n13023, MEM_stage_inst_dmem_n13022, MEM_stage_inst_dmem_n13021, MEM_stage_inst_dmem_n13020, MEM_stage_inst_dmem_n13019, MEM_stage_inst_dmem_n13018, MEM_stage_inst_dmem_n13017, MEM_stage_inst_dmem_n13016, MEM_stage_inst_dmem_n13015, MEM_stage_inst_dmem_n13014, MEM_stage_inst_dmem_n13013, MEM_stage_inst_dmem_n13012, MEM_stage_inst_dmem_n13011, MEM_stage_inst_dmem_n13010, MEM_stage_inst_dmem_n13009, MEM_stage_inst_dmem_n13008, MEM_stage_inst_dmem_n13007, MEM_stage_inst_dmem_n13006, MEM_stage_inst_dmem_n13005, MEM_stage_inst_dmem_n13004, MEM_stage_inst_dmem_n13003, MEM_stage_inst_dmem_n13002, MEM_stage_inst_dmem_n13001, MEM_stage_inst_dmem_n13000, MEM_stage_inst_dmem_n12999, MEM_stage_inst_dmem_n12998, MEM_stage_inst_dmem_n12997, MEM_stage_inst_dmem_n12996, MEM_stage_inst_dmem_n12995, MEM_stage_inst_dmem_n12994, MEM_stage_inst_dmem_n12993, MEM_stage_inst_dmem_n12992, MEM_stage_inst_dmem_n12991, MEM_stage_inst_dmem_n12990, MEM_stage_inst_dmem_n12989, MEM_stage_inst_dmem_n12988, MEM_stage_inst_dmem_n12987, MEM_stage_inst_dmem_n12986, MEM_stage_inst_dmem_n12985, MEM_stage_inst_dmem_n12984, MEM_stage_inst_dmem_n12983, MEM_stage_inst_dmem_n12982, MEM_stage_inst_dmem_n12981, MEM_stage_inst_dmem_n12980, MEM_stage_inst_dmem_n12979, MEM_stage_inst_dmem_n12978, MEM_stage_inst_dmem_n12977, MEM_stage_inst_dmem_n12976, MEM_stage_inst_dmem_n12975, MEM_stage_inst_dmem_n12974, MEM_stage_inst_dmem_n12973, MEM_stage_inst_dmem_n12972, MEM_stage_inst_dmem_n12971, MEM_stage_inst_dmem_n12970, MEM_stage_inst_dmem_n12969, MEM_stage_inst_dmem_n12968, MEM_stage_inst_dmem_n12967, MEM_stage_inst_dmem_n12966, MEM_stage_inst_dmem_n12965, MEM_stage_inst_dmem_n12964, MEM_stage_inst_dmem_n12963, MEM_stage_inst_dmem_n12962, MEM_stage_inst_dmem_n12961, MEM_stage_inst_dmem_n12960, MEM_stage_inst_dmem_n12959, MEM_stage_inst_dmem_n12958, MEM_stage_inst_dmem_n12957, MEM_stage_inst_dmem_n12956, MEM_stage_inst_dmem_n12955, MEM_stage_inst_dmem_n12954, MEM_stage_inst_dmem_n12953, MEM_stage_inst_dmem_n12952, MEM_stage_inst_dmem_n12951, MEM_stage_inst_dmem_n12950, MEM_stage_inst_dmem_n12949, MEM_stage_inst_dmem_n12948, MEM_stage_inst_dmem_n12947, MEM_stage_inst_dmem_n12946, MEM_stage_inst_dmem_n12945, MEM_stage_inst_dmem_n12944, MEM_stage_inst_dmem_n12943, MEM_stage_inst_dmem_n12942, MEM_stage_inst_dmem_n12941, MEM_stage_inst_dmem_n12940, MEM_stage_inst_dmem_n12939, MEM_stage_inst_dmem_n12938, MEM_stage_inst_dmem_n12937, MEM_stage_inst_dmem_n12936, MEM_stage_inst_dmem_n12935, MEM_stage_inst_dmem_n12934, MEM_stage_inst_dmem_n12933, MEM_stage_inst_dmem_n12932, MEM_stage_inst_dmem_n12931, MEM_stage_inst_dmem_n12930, MEM_stage_inst_dmem_n12929, MEM_stage_inst_dmem_n12928, MEM_stage_inst_dmem_n12927, MEM_stage_inst_dmem_n12926, MEM_stage_inst_dmem_n12925, MEM_stage_inst_dmem_n12924, MEM_stage_inst_dmem_n12923, MEM_stage_inst_dmem_n12922, MEM_stage_inst_dmem_n12921, MEM_stage_inst_dmem_n12920, MEM_stage_inst_dmem_n12919, MEM_stage_inst_dmem_n12918, MEM_stage_inst_dmem_n12917, MEM_stage_inst_dmem_n12916, MEM_stage_inst_dmem_n12915, MEM_stage_inst_dmem_n12914, MEM_stage_inst_dmem_n12913, MEM_stage_inst_dmem_n12912, MEM_stage_inst_dmem_n12911, MEM_stage_inst_dmem_n12910, MEM_stage_inst_dmem_n12909, MEM_stage_inst_dmem_n12908, MEM_stage_inst_dmem_n12907, MEM_stage_inst_dmem_n12906, MEM_stage_inst_dmem_n12905, MEM_stage_inst_dmem_n12904, MEM_stage_inst_dmem_n12903, MEM_stage_inst_dmem_n12902, MEM_stage_inst_dmem_n12901, MEM_stage_inst_dmem_n12900, MEM_stage_inst_dmem_n12899, MEM_stage_inst_dmem_n12898, MEM_stage_inst_dmem_n12897, MEM_stage_inst_dmem_n12896, MEM_stage_inst_dmem_n12895, MEM_stage_inst_dmem_n12894, MEM_stage_inst_dmem_n12893, MEM_stage_inst_dmem_n12892, MEM_stage_inst_dmem_n12891, MEM_stage_inst_dmem_n12890, MEM_stage_inst_dmem_n12889, MEM_stage_inst_dmem_n12888, MEM_stage_inst_dmem_n12887, MEM_stage_inst_dmem_n12886, MEM_stage_inst_dmem_n12885, MEM_stage_inst_dmem_n12884, MEM_stage_inst_dmem_n12883, MEM_stage_inst_dmem_n12882, MEM_stage_inst_dmem_n12881, MEM_stage_inst_dmem_n12880, MEM_stage_inst_dmem_n12879, MEM_stage_inst_dmem_n12878, MEM_stage_inst_dmem_n12877, MEM_stage_inst_dmem_n12876, MEM_stage_inst_dmem_n12875, MEM_stage_inst_dmem_n12874, MEM_stage_inst_dmem_n12873, MEM_stage_inst_dmem_n12872, MEM_stage_inst_dmem_n12871, MEM_stage_inst_dmem_n12870, MEM_stage_inst_dmem_n12869, MEM_stage_inst_dmem_n12868, MEM_stage_inst_dmem_n12867, MEM_stage_inst_dmem_n12866, MEM_stage_inst_dmem_n12865, MEM_stage_inst_dmem_n12864, MEM_stage_inst_dmem_n12863, MEM_stage_inst_dmem_n12862, MEM_stage_inst_dmem_n12861, MEM_stage_inst_dmem_n12860, MEM_stage_inst_dmem_n12859, MEM_stage_inst_dmem_n8762, MEM_stage_inst_dmem_n8761, MEM_stage_inst_dmem_n8760, MEM_stage_inst_dmem_n8759, MEM_stage_inst_dmem_n8758, MEM_stage_inst_dmem_n8757, MEM_stage_inst_dmem_n8756, MEM_stage_inst_dmem_n8755, MEM_stage_inst_dmem_n8754, MEM_stage_inst_dmem_n8753, MEM_stage_inst_dmem_n8752, MEM_stage_inst_dmem_n8751, MEM_stage_inst_dmem_n8750, MEM_stage_inst_dmem_n8749, MEM_stage_inst_dmem_n8748, MEM_stage_inst_dmem_n8747, MEM_stage_inst_dmem_n8746, MEM_stage_inst_dmem_n8745, MEM_stage_inst_dmem_n8744, MEM_stage_inst_dmem_n8743, MEM_stage_inst_dmem_n8742, MEM_stage_inst_dmem_n8741, MEM_stage_inst_dmem_n8740, MEM_stage_inst_dmem_n8739, MEM_stage_inst_dmem_n8738, MEM_stage_inst_dmem_n8737, MEM_stage_inst_dmem_n8736, MEM_stage_inst_dmem_n8735, MEM_stage_inst_dmem_n8734, MEM_stage_inst_dmem_n8733, MEM_stage_inst_dmem_n8732, MEM_stage_inst_dmem_n8731, MEM_stage_inst_dmem_n8730, MEM_stage_inst_dmem_n8729, MEM_stage_inst_dmem_n8728, MEM_stage_inst_dmem_n8727, MEM_stage_inst_dmem_n8726, MEM_stage_inst_dmem_n8725, MEM_stage_inst_dmem_n8724, MEM_stage_inst_dmem_n8723, MEM_stage_inst_dmem_n8722, MEM_stage_inst_dmem_n8721, MEM_stage_inst_dmem_n8720, MEM_stage_inst_dmem_n8719, MEM_stage_inst_dmem_n8718, MEM_stage_inst_dmem_n8717, MEM_stage_inst_dmem_n8716, MEM_stage_inst_dmem_n8715, MEM_stage_inst_dmem_n8714, MEM_stage_inst_dmem_n8713, MEM_stage_inst_dmem_n8712, MEM_stage_inst_dmem_n8711, MEM_stage_inst_dmem_n8710, MEM_stage_inst_dmem_n8709, MEM_stage_inst_dmem_n8708, MEM_stage_inst_dmem_n8707, MEM_stage_inst_dmem_n8706, MEM_stage_inst_dmem_n8705, MEM_stage_inst_dmem_n8704, MEM_stage_inst_dmem_n8703, MEM_stage_inst_dmem_n8702, MEM_stage_inst_dmem_n8701, MEM_stage_inst_dmem_n8700, MEM_stage_inst_dmem_n8699, MEM_stage_inst_dmem_n8698, MEM_stage_inst_dmem_n8697, MEM_stage_inst_dmem_n8696, MEM_stage_inst_dmem_n8695, MEM_stage_inst_dmem_n8694, MEM_stage_inst_dmem_n8693, MEM_stage_inst_dmem_n8692, MEM_stage_inst_dmem_n8691, MEM_stage_inst_dmem_n8690, MEM_stage_inst_dmem_n8689, MEM_stage_inst_dmem_n8688, MEM_stage_inst_dmem_n8687, MEM_stage_inst_dmem_n8686, MEM_stage_inst_dmem_n8685, MEM_stage_inst_dmem_n8684, MEM_stage_inst_dmem_n8683, MEM_stage_inst_dmem_n8682, MEM_stage_inst_dmem_n8681, MEM_stage_inst_dmem_n8680, MEM_stage_inst_dmem_n8679, MEM_stage_inst_dmem_n8678, MEM_stage_inst_dmem_n8677, MEM_stage_inst_dmem_n8676, MEM_stage_inst_dmem_n8675, MEM_stage_inst_dmem_n8674, MEM_stage_inst_dmem_n8673, MEM_stage_inst_dmem_n8672, MEM_stage_inst_dmem_n8671, MEM_stage_inst_dmem_n8670, MEM_stage_inst_dmem_n8669, MEM_stage_inst_dmem_n8668, MEM_stage_inst_dmem_n8667, MEM_stage_inst_dmem_n8666, MEM_stage_inst_dmem_n8665, MEM_stage_inst_dmem_n8664, MEM_stage_inst_dmem_n8663, MEM_stage_inst_dmem_n8662, MEM_stage_inst_dmem_n8661, MEM_stage_inst_dmem_n8660, MEM_stage_inst_dmem_n8659, MEM_stage_inst_dmem_n8658, MEM_stage_inst_dmem_n8657, MEM_stage_inst_dmem_n8656, MEM_stage_inst_dmem_n8655, MEM_stage_inst_dmem_n8654, MEM_stage_inst_dmem_n8653, MEM_stage_inst_dmem_n8652, MEM_stage_inst_dmem_n8651, MEM_stage_inst_dmem_n8650, MEM_stage_inst_dmem_n8649, MEM_stage_inst_dmem_n8648, MEM_stage_inst_dmem_n8647, MEM_stage_inst_dmem_n8646, MEM_stage_inst_dmem_n8645, MEM_stage_inst_dmem_n8644, MEM_stage_inst_dmem_n8643, MEM_stage_inst_dmem_n8642, MEM_stage_inst_dmem_n8641, MEM_stage_inst_dmem_n8640, MEM_stage_inst_dmem_n8639, MEM_stage_inst_dmem_n8638, MEM_stage_inst_dmem_n8637, MEM_stage_inst_dmem_n8636, MEM_stage_inst_dmem_n8635, MEM_stage_inst_dmem_n8634, MEM_stage_inst_dmem_n8633, MEM_stage_inst_dmem_n8632, MEM_stage_inst_dmem_n8631, MEM_stage_inst_dmem_n8630, MEM_stage_inst_dmem_n8629, MEM_stage_inst_dmem_n8628, MEM_stage_inst_dmem_n8627, MEM_stage_inst_dmem_n8626, MEM_stage_inst_dmem_n8625, MEM_stage_inst_dmem_n8624, MEM_stage_inst_dmem_n8623, MEM_stage_inst_dmem_n8622, MEM_stage_inst_dmem_n8621, MEM_stage_inst_dmem_n8620, MEM_stage_inst_dmem_n8619, MEM_stage_inst_dmem_n8618, MEM_stage_inst_dmem_n8617, MEM_stage_inst_dmem_n8616, MEM_stage_inst_dmem_n8615, MEM_stage_inst_dmem_n8614, MEM_stage_inst_dmem_n8613, MEM_stage_inst_dmem_n8612, MEM_stage_inst_dmem_n8611, MEM_stage_inst_dmem_n8610, MEM_stage_inst_dmem_n8609, MEM_stage_inst_dmem_n8608, MEM_stage_inst_dmem_n8607, MEM_stage_inst_dmem_n8606, MEM_stage_inst_dmem_n8605, MEM_stage_inst_dmem_n8604, MEM_stage_inst_dmem_n8603, MEM_stage_inst_dmem_n8602, MEM_stage_inst_dmem_n8601, MEM_stage_inst_dmem_n8600, MEM_stage_inst_dmem_n8599, MEM_stage_inst_dmem_n8598, MEM_stage_inst_dmem_n8597, MEM_stage_inst_dmem_n8596, MEM_stage_inst_dmem_n8595, MEM_stage_inst_dmem_n8594, MEM_stage_inst_dmem_n8593, MEM_stage_inst_dmem_n8592, MEM_stage_inst_dmem_n8591, MEM_stage_inst_dmem_n8590, MEM_stage_inst_dmem_n8589, MEM_stage_inst_dmem_n8588, MEM_stage_inst_dmem_n8587, MEM_stage_inst_dmem_n8586, MEM_stage_inst_dmem_n8585, MEM_stage_inst_dmem_n8584, MEM_stage_inst_dmem_n8583, MEM_stage_inst_dmem_n8582, MEM_stage_inst_dmem_n8581, MEM_stage_inst_dmem_n8580, MEM_stage_inst_dmem_n8579, MEM_stage_inst_dmem_n8578, MEM_stage_inst_dmem_n8577, MEM_stage_inst_dmem_n8576, MEM_stage_inst_dmem_n8575, MEM_stage_inst_dmem_n8574, MEM_stage_inst_dmem_n8573, MEM_stage_inst_dmem_n8572, MEM_stage_inst_dmem_n8571, MEM_stage_inst_dmem_n8570, MEM_stage_inst_dmem_n8569, MEM_stage_inst_dmem_n8568, MEM_stage_inst_dmem_n8567, MEM_stage_inst_dmem_n8566, MEM_stage_inst_dmem_n8565, MEM_stage_inst_dmem_n8564, MEM_stage_inst_dmem_n8563, MEM_stage_inst_dmem_n8562, MEM_stage_inst_dmem_n8561, MEM_stage_inst_dmem_n8560, MEM_stage_inst_dmem_n8559, MEM_stage_inst_dmem_n8558, MEM_stage_inst_dmem_n8557, MEM_stage_inst_dmem_n8556, MEM_stage_inst_dmem_n8555, MEM_stage_inst_dmem_n8554, MEM_stage_inst_dmem_n8553, MEM_stage_inst_dmem_n8552, MEM_stage_inst_dmem_n8551, MEM_stage_inst_dmem_n8550, MEM_stage_inst_dmem_n8549, MEM_stage_inst_dmem_n8548, MEM_stage_inst_dmem_n8547, MEM_stage_inst_dmem_n8546, MEM_stage_inst_dmem_n8545, MEM_stage_inst_dmem_n8544, MEM_stage_inst_dmem_n8543, MEM_stage_inst_dmem_n8542, MEM_stage_inst_dmem_n8541, MEM_stage_inst_dmem_n8540, MEM_stage_inst_dmem_n8539, MEM_stage_inst_dmem_n8538, MEM_stage_inst_dmem_n8537, MEM_stage_inst_dmem_n8536, MEM_stage_inst_dmem_n8535, MEM_stage_inst_dmem_n8534, MEM_stage_inst_dmem_n8533, MEM_stage_inst_dmem_n8532, MEM_stage_inst_dmem_n8531, MEM_stage_inst_dmem_n8530, MEM_stage_inst_dmem_n8529, MEM_stage_inst_dmem_n8528, MEM_stage_inst_dmem_n8527, MEM_stage_inst_dmem_n8526, MEM_stage_inst_dmem_n8525, MEM_stage_inst_dmem_n8524, MEM_stage_inst_dmem_n8523, MEM_stage_inst_dmem_n8522, MEM_stage_inst_dmem_n8521, MEM_stage_inst_dmem_n8520, MEM_stage_inst_dmem_n8519, MEM_stage_inst_dmem_n8518, MEM_stage_inst_dmem_n8517, MEM_stage_inst_dmem_n8516, MEM_stage_inst_dmem_n8515, MEM_stage_inst_dmem_n8514, MEM_stage_inst_dmem_n8513, MEM_stage_inst_dmem_n8512, MEM_stage_inst_dmem_n8511, MEM_stage_inst_dmem_n8510, MEM_stage_inst_dmem_n8509, MEM_stage_inst_dmem_n8508, MEM_stage_inst_dmem_n8507, MEM_stage_inst_dmem_n8506, MEM_stage_inst_dmem_n8505, MEM_stage_inst_dmem_n8504, MEM_stage_inst_dmem_n8503, MEM_stage_inst_dmem_n8502, MEM_stage_inst_dmem_n8501, MEM_stage_inst_dmem_n8500, MEM_stage_inst_dmem_n8499, MEM_stage_inst_dmem_n8498, MEM_stage_inst_dmem_n8497, MEM_stage_inst_dmem_n8496, MEM_stage_inst_dmem_n8495, MEM_stage_inst_dmem_n8494, MEM_stage_inst_dmem_n8493, MEM_stage_inst_dmem_n8492, MEM_stage_inst_dmem_n8491, MEM_stage_inst_dmem_n8490, MEM_stage_inst_dmem_n8489, MEM_stage_inst_dmem_n8488, MEM_stage_inst_dmem_n8487, MEM_stage_inst_dmem_n8486, MEM_stage_inst_dmem_n8485, MEM_stage_inst_dmem_n8484, MEM_stage_inst_dmem_n8483, MEM_stage_inst_dmem_n8482, MEM_stage_inst_dmem_n8481, MEM_stage_inst_dmem_n8480, MEM_stage_inst_dmem_n8479, MEM_stage_inst_dmem_n8478, MEM_stage_inst_dmem_n8477, MEM_stage_inst_dmem_n8476, MEM_stage_inst_dmem_n8475, MEM_stage_inst_dmem_n8474, MEM_stage_inst_dmem_n8473, MEM_stage_inst_dmem_n8472, MEM_stage_inst_dmem_n8471, MEM_stage_inst_dmem_n8470, MEM_stage_inst_dmem_n8469, MEM_stage_inst_dmem_n8468, MEM_stage_inst_dmem_n8467, MEM_stage_inst_dmem_n8466, MEM_stage_inst_dmem_n8465, MEM_stage_inst_dmem_n8464, MEM_stage_inst_dmem_n8463, MEM_stage_inst_dmem_n8462, MEM_stage_inst_dmem_n8461, MEM_stage_inst_dmem_n8460, MEM_stage_inst_dmem_n8459, MEM_stage_inst_dmem_n8458, MEM_stage_inst_dmem_n8457, MEM_stage_inst_dmem_n8456, MEM_stage_inst_dmem_n8455, MEM_stage_inst_dmem_n8454, MEM_stage_inst_dmem_n8453, MEM_stage_inst_dmem_n8452, MEM_stage_inst_dmem_n8451, MEM_stage_inst_dmem_n8450, MEM_stage_inst_dmem_n8449, MEM_stage_inst_dmem_n8448, MEM_stage_inst_dmem_n8447, MEM_stage_inst_dmem_n8446, MEM_stage_inst_dmem_n8445, MEM_stage_inst_dmem_n8444, MEM_stage_inst_dmem_n8443, MEM_stage_inst_dmem_n8442, MEM_stage_inst_dmem_n8441, MEM_stage_inst_dmem_n8440, MEM_stage_inst_dmem_n8439, MEM_stage_inst_dmem_n8438, MEM_stage_inst_dmem_n8437, MEM_stage_inst_dmem_n8436, MEM_stage_inst_dmem_n8435, MEM_stage_inst_dmem_n8434, MEM_stage_inst_dmem_n8433, MEM_stage_inst_dmem_n8432, MEM_stage_inst_dmem_n8431, MEM_stage_inst_dmem_n8430, MEM_stage_inst_dmem_n8429, MEM_stage_inst_dmem_n8428, MEM_stage_inst_dmem_n8427, MEM_stage_inst_dmem_n8426, MEM_stage_inst_dmem_n8425, MEM_stage_inst_dmem_n8424, MEM_stage_inst_dmem_n8423, MEM_stage_inst_dmem_n8422, MEM_stage_inst_dmem_n8421, MEM_stage_inst_dmem_n8420, MEM_stage_inst_dmem_n8419, MEM_stage_inst_dmem_n8418, MEM_stage_inst_dmem_n8417, MEM_stage_inst_dmem_n8416, MEM_stage_inst_dmem_n8415, MEM_stage_inst_dmem_n8414, MEM_stage_inst_dmem_n8413, MEM_stage_inst_dmem_n8412, MEM_stage_inst_dmem_n8411, MEM_stage_inst_dmem_n8410, MEM_stage_inst_dmem_n8409, MEM_stage_inst_dmem_n8408, MEM_stage_inst_dmem_n8407, MEM_stage_inst_dmem_n8406, MEM_stage_inst_dmem_n8405, MEM_stage_inst_dmem_n8404, MEM_stage_inst_dmem_n8403, MEM_stage_inst_dmem_n8402, MEM_stage_inst_dmem_n8401, MEM_stage_inst_dmem_n8400, MEM_stage_inst_dmem_n8399, MEM_stage_inst_dmem_n8398, MEM_stage_inst_dmem_n8397, MEM_stage_inst_dmem_n8396, MEM_stage_inst_dmem_n8395, MEM_stage_inst_dmem_n8394, MEM_stage_inst_dmem_n8393, MEM_stage_inst_dmem_n8392, MEM_stage_inst_dmem_n8391, MEM_stage_inst_dmem_n8390, MEM_stage_inst_dmem_n8389, MEM_stage_inst_dmem_n8388, MEM_stage_inst_dmem_n8387, MEM_stage_inst_dmem_n8386, MEM_stage_inst_dmem_n8385, MEM_stage_inst_dmem_n8384, MEM_stage_inst_dmem_n8383, MEM_stage_inst_dmem_n8382, MEM_stage_inst_dmem_n8381, MEM_stage_inst_dmem_n8380, MEM_stage_inst_dmem_n8379, MEM_stage_inst_dmem_n8378, MEM_stage_inst_dmem_n8377, MEM_stage_inst_dmem_n8376, MEM_stage_inst_dmem_n8375, MEM_stage_inst_dmem_n8374, MEM_stage_inst_dmem_n8373, MEM_stage_inst_dmem_n8372, MEM_stage_inst_dmem_n8371, MEM_stage_inst_dmem_n8370, MEM_stage_inst_dmem_n8369, MEM_stage_inst_dmem_n8368, MEM_stage_inst_dmem_n8367, MEM_stage_inst_dmem_n8366, MEM_stage_inst_dmem_n8365, MEM_stage_inst_dmem_n8364, MEM_stage_inst_dmem_n8363, MEM_stage_inst_dmem_n8362, MEM_stage_inst_dmem_n8361, MEM_stage_inst_dmem_n8360, MEM_stage_inst_dmem_n8359, MEM_stage_inst_dmem_n8358, MEM_stage_inst_dmem_n8357, MEM_stage_inst_dmem_n8356, MEM_stage_inst_dmem_n8355, MEM_stage_inst_dmem_n8354, MEM_stage_inst_dmem_n8353, MEM_stage_inst_dmem_n8352, MEM_stage_inst_dmem_n8351, MEM_stage_inst_dmem_n8350, MEM_stage_inst_dmem_n8349, MEM_stage_inst_dmem_n8348, MEM_stage_inst_dmem_n8347, MEM_stage_inst_dmem_n8346, MEM_stage_inst_dmem_n8345, MEM_stage_inst_dmem_n8344, MEM_stage_inst_dmem_n8343, MEM_stage_inst_dmem_n8342, MEM_stage_inst_dmem_n8341, MEM_stage_inst_dmem_n8340, MEM_stage_inst_dmem_n8339, MEM_stage_inst_dmem_n8338, MEM_stage_inst_dmem_n8337, MEM_stage_inst_dmem_n8336, MEM_stage_inst_dmem_n8335, MEM_stage_inst_dmem_n8334, MEM_stage_inst_dmem_n8333, MEM_stage_inst_dmem_n8332, MEM_stage_inst_dmem_n8331, MEM_stage_inst_dmem_n8330, MEM_stage_inst_dmem_n8329, MEM_stage_inst_dmem_n8328, MEM_stage_inst_dmem_n8327, MEM_stage_inst_dmem_n8326, MEM_stage_inst_dmem_n8325, MEM_stage_inst_dmem_n8324, MEM_stage_inst_dmem_n8323, MEM_stage_inst_dmem_n8322, MEM_stage_inst_dmem_n8321, MEM_stage_inst_dmem_n8320, MEM_stage_inst_dmem_n8319, MEM_stage_inst_dmem_n8318, MEM_stage_inst_dmem_n8317, MEM_stage_inst_dmem_n8316, MEM_stage_inst_dmem_n8315, MEM_stage_inst_dmem_n8314, MEM_stage_inst_dmem_n8313, MEM_stage_inst_dmem_n8312, MEM_stage_inst_dmem_n8311, MEM_stage_inst_dmem_n8310, MEM_stage_inst_dmem_n8309, MEM_stage_inst_dmem_n8308, MEM_stage_inst_dmem_n8307, MEM_stage_inst_dmem_n8306, MEM_stage_inst_dmem_n8305, MEM_stage_inst_dmem_n8304, MEM_stage_inst_dmem_n8303, MEM_stage_inst_dmem_n8302, MEM_stage_inst_dmem_n8301, MEM_stage_inst_dmem_n8300, MEM_stage_inst_dmem_n8299, MEM_stage_inst_dmem_n8298, MEM_stage_inst_dmem_n8297, MEM_stage_inst_dmem_n8296, MEM_stage_inst_dmem_n8295, MEM_stage_inst_dmem_n8294, MEM_stage_inst_dmem_n8293, MEM_stage_inst_dmem_n8292, MEM_stage_inst_dmem_n8291, MEM_stage_inst_dmem_n8290, MEM_stage_inst_dmem_n8289, MEM_stage_inst_dmem_n8288, MEM_stage_inst_dmem_n8287, MEM_stage_inst_dmem_n8286, MEM_stage_inst_dmem_n8285, MEM_stage_inst_dmem_n8284, MEM_stage_inst_dmem_n8283, MEM_stage_inst_dmem_n8282, MEM_stage_inst_dmem_n8281, MEM_stage_inst_dmem_n8280, MEM_stage_inst_dmem_n8279, MEM_stage_inst_dmem_n8278, MEM_stage_inst_dmem_n8277, MEM_stage_inst_dmem_n8276, MEM_stage_inst_dmem_n8275, MEM_stage_inst_dmem_n8274, MEM_stage_inst_dmem_n8273, MEM_stage_inst_dmem_n8272, MEM_stage_inst_dmem_n8271, MEM_stage_inst_dmem_n8270, MEM_stage_inst_dmem_n8269, MEM_stage_inst_dmem_n8268, MEM_stage_inst_dmem_n8267, MEM_stage_inst_dmem_n8266, MEM_stage_inst_dmem_n8265, MEM_stage_inst_dmem_n8264, MEM_stage_inst_dmem_n8263, MEM_stage_inst_dmem_n8262, MEM_stage_inst_dmem_n8261, MEM_stage_inst_dmem_n8260, MEM_stage_inst_dmem_n8259, MEM_stage_inst_dmem_n8258, MEM_stage_inst_dmem_n8257, MEM_stage_inst_dmem_n8256, MEM_stage_inst_dmem_n8255, MEM_stage_inst_dmem_n8254, MEM_stage_inst_dmem_n8253, MEM_stage_inst_dmem_n8252, MEM_stage_inst_dmem_n8251, MEM_stage_inst_dmem_n8250, MEM_stage_inst_dmem_n8249, MEM_stage_inst_dmem_n8248, MEM_stage_inst_dmem_n8247, MEM_stage_inst_dmem_n8246, MEM_stage_inst_dmem_n8245, MEM_stage_inst_dmem_n8244, MEM_stage_inst_dmem_n8243, MEM_stage_inst_dmem_n8242, MEM_stage_inst_dmem_n8241, MEM_stage_inst_dmem_n8240, MEM_stage_inst_dmem_n8239, MEM_stage_inst_dmem_n8238, MEM_stage_inst_dmem_n8237, MEM_stage_inst_dmem_n8236, MEM_stage_inst_dmem_n8235, MEM_stage_inst_dmem_n8234, MEM_stage_inst_dmem_n8233, MEM_stage_inst_dmem_n8232, MEM_stage_inst_dmem_n8231, MEM_stage_inst_dmem_n8230, MEM_stage_inst_dmem_n8229, MEM_stage_inst_dmem_n8228, MEM_stage_inst_dmem_n8227, MEM_stage_inst_dmem_n8226, MEM_stage_inst_dmem_n8225, MEM_stage_inst_dmem_n8224, MEM_stage_inst_dmem_n8223, MEM_stage_inst_dmem_n8222, MEM_stage_inst_dmem_n8221, MEM_stage_inst_dmem_n8220, MEM_stage_inst_dmem_n8219, MEM_stage_inst_dmem_n8218, MEM_stage_inst_dmem_n8217, MEM_stage_inst_dmem_n8216, MEM_stage_inst_dmem_n8215, MEM_stage_inst_dmem_n8214, MEM_stage_inst_dmem_n8213, MEM_stage_inst_dmem_n8212, MEM_stage_inst_dmem_n8211, MEM_stage_inst_dmem_n8210, MEM_stage_inst_dmem_n8209, MEM_stage_inst_dmem_n8208, MEM_stage_inst_dmem_n8207, MEM_stage_inst_dmem_n8206, MEM_stage_inst_dmem_n8205, MEM_stage_inst_dmem_n8204, MEM_stage_inst_dmem_n8203, MEM_stage_inst_dmem_n8202, MEM_stage_inst_dmem_n8201, MEM_stage_inst_dmem_n8200, MEM_stage_inst_dmem_n8199, MEM_stage_inst_dmem_n8198, MEM_stage_inst_dmem_n8197, MEM_stage_inst_dmem_n8196, MEM_stage_inst_dmem_n8195, MEM_stage_inst_dmem_n8194, MEM_stage_inst_dmem_n8193, MEM_stage_inst_dmem_n8192, MEM_stage_inst_dmem_n8191, MEM_stage_inst_dmem_n8190, MEM_stage_inst_dmem_n8189, MEM_stage_inst_dmem_n8188, MEM_stage_inst_dmem_n8187, MEM_stage_inst_dmem_n8186, MEM_stage_inst_dmem_n8185, MEM_stage_inst_dmem_n8184, MEM_stage_inst_dmem_n8183, MEM_stage_inst_dmem_n8182, MEM_stage_inst_dmem_n8181, MEM_stage_inst_dmem_n8180, MEM_stage_inst_dmem_n8179, MEM_stage_inst_dmem_n8178, MEM_stage_inst_dmem_n8177, MEM_stage_inst_dmem_n8176, MEM_stage_inst_dmem_n8175, MEM_stage_inst_dmem_n8174, MEM_stage_inst_dmem_n8173, MEM_stage_inst_dmem_n8172, MEM_stage_inst_dmem_n8171, MEM_stage_inst_dmem_n8170, MEM_stage_inst_dmem_n8169, MEM_stage_inst_dmem_n8168, MEM_stage_inst_dmem_n8167, MEM_stage_inst_dmem_n8166, MEM_stage_inst_dmem_n8165, MEM_stage_inst_dmem_n8164, MEM_stage_inst_dmem_n8163, MEM_stage_inst_dmem_n8162, MEM_stage_inst_dmem_n8161, MEM_stage_inst_dmem_n8160, MEM_stage_inst_dmem_n8159, MEM_stage_inst_dmem_n8158, MEM_stage_inst_dmem_n8157, MEM_stage_inst_dmem_n8156, MEM_stage_inst_dmem_n8155, MEM_stage_inst_dmem_n8154, MEM_stage_inst_dmem_n8153, MEM_stage_inst_dmem_n8152, MEM_stage_inst_dmem_n8151, MEM_stage_inst_dmem_n8150, MEM_stage_inst_dmem_n8149, MEM_stage_inst_dmem_n8148, MEM_stage_inst_dmem_n8147, MEM_stage_inst_dmem_n8146, MEM_stage_inst_dmem_n8145, MEM_stage_inst_dmem_n8144, MEM_stage_inst_dmem_n8143, MEM_stage_inst_dmem_n8142, MEM_stage_inst_dmem_n8141, MEM_stage_inst_dmem_n8140, MEM_stage_inst_dmem_n8139, MEM_stage_inst_dmem_n8138, MEM_stage_inst_dmem_n8137, MEM_stage_inst_dmem_n8136, MEM_stage_inst_dmem_n8135, MEM_stage_inst_dmem_n8134, MEM_stage_inst_dmem_n8133, MEM_stage_inst_dmem_n8132, MEM_stage_inst_dmem_n8131, MEM_stage_inst_dmem_n8130, MEM_stage_inst_dmem_n8129, MEM_stage_inst_dmem_n8128, MEM_stage_inst_dmem_n8127, MEM_stage_inst_dmem_n8126, MEM_stage_inst_dmem_n8125, MEM_stage_inst_dmem_n8124, MEM_stage_inst_dmem_n8123, MEM_stage_inst_dmem_n8122, MEM_stage_inst_dmem_n8121, MEM_stage_inst_dmem_n8120, MEM_stage_inst_dmem_n8119, MEM_stage_inst_dmem_n8118, MEM_stage_inst_dmem_n8117, MEM_stage_inst_dmem_n8116, MEM_stage_inst_dmem_n8115, MEM_stage_inst_dmem_n8114, MEM_stage_inst_dmem_n8113, MEM_stage_inst_dmem_n8112, MEM_stage_inst_dmem_n8111, MEM_stage_inst_dmem_n8110, MEM_stage_inst_dmem_n8109, MEM_stage_inst_dmem_n8108, MEM_stage_inst_dmem_n8107, MEM_stage_inst_dmem_n8106, MEM_stage_inst_dmem_n8105, MEM_stage_inst_dmem_n8104, MEM_stage_inst_dmem_n8103, MEM_stage_inst_dmem_n8102, MEM_stage_inst_dmem_n8101, MEM_stage_inst_dmem_n8100, MEM_stage_inst_dmem_n8099, MEM_stage_inst_dmem_n8098, MEM_stage_inst_dmem_n8097, MEM_stage_inst_dmem_n8096, MEM_stage_inst_dmem_n8095, MEM_stage_inst_dmem_n8094, MEM_stage_inst_dmem_n8093, MEM_stage_inst_dmem_n8092, MEM_stage_inst_dmem_n8091, MEM_stage_inst_dmem_n8090, MEM_stage_inst_dmem_n8089, MEM_stage_inst_dmem_n8088, MEM_stage_inst_dmem_n8087, MEM_stage_inst_dmem_n8086, MEM_stage_inst_dmem_n8085, MEM_stage_inst_dmem_n8084, MEM_stage_inst_dmem_n8083, MEM_stage_inst_dmem_n8082, MEM_stage_inst_dmem_n8081, MEM_stage_inst_dmem_n8080, MEM_stage_inst_dmem_n8079, MEM_stage_inst_dmem_n8078, MEM_stage_inst_dmem_n8077, MEM_stage_inst_dmem_n8076, MEM_stage_inst_dmem_n8075, MEM_stage_inst_dmem_n8074, MEM_stage_inst_dmem_n8073, MEM_stage_inst_dmem_n8072, MEM_stage_inst_dmem_n8071, MEM_stage_inst_dmem_n8070, MEM_stage_inst_dmem_n8069, MEM_stage_inst_dmem_n8068, MEM_stage_inst_dmem_n8067, MEM_stage_inst_dmem_n8066, MEM_stage_inst_dmem_n8065, MEM_stage_inst_dmem_n8064, MEM_stage_inst_dmem_n8063, MEM_stage_inst_dmem_n8062, MEM_stage_inst_dmem_n8061, MEM_stage_inst_dmem_n8060, MEM_stage_inst_dmem_n8059, MEM_stage_inst_dmem_n8058, MEM_stage_inst_dmem_n8057, MEM_stage_inst_dmem_n8056, MEM_stage_inst_dmem_n8055, MEM_stage_inst_dmem_n8054, MEM_stage_inst_dmem_n8053, MEM_stage_inst_dmem_n8052, MEM_stage_inst_dmem_n8051, MEM_stage_inst_dmem_n8050, MEM_stage_inst_dmem_n8049, MEM_stage_inst_dmem_n8048, MEM_stage_inst_dmem_n8047, MEM_stage_inst_dmem_n8046, MEM_stage_inst_dmem_n8045, MEM_stage_inst_dmem_n8044, MEM_stage_inst_dmem_n8043, MEM_stage_inst_dmem_n8042, MEM_stage_inst_dmem_n8041, MEM_stage_inst_dmem_n8040, MEM_stage_inst_dmem_n8039, MEM_stage_inst_dmem_n8038, MEM_stage_inst_dmem_n8037, MEM_stage_inst_dmem_n8036, MEM_stage_inst_dmem_n8035, MEM_stage_inst_dmem_n8034, MEM_stage_inst_dmem_n8033, MEM_stage_inst_dmem_n8032, MEM_stage_inst_dmem_n8031, MEM_stage_inst_dmem_n8030, MEM_stage_inst_dmem_n8029, MEM_stage_inst_dmem_n8028, MEM_stage_inst_dmem_n8027, MEM_stage_inst_dmem_n8026, MEM_stage_inst_dmem_n8025, MEM_stage_inst_dmem_n8024, MEM_stage_inst_dmem_n8023, MEM_stage_inst_dmem_n8022, MEM_stage_inst_dmem_n8021, MEM_stage_inst_dmem_n8020, MEM_stage_inst_dmem_n8019, MEM_stage_inst_dmem_n8018, MEM_stage_inst_dmem_n8017, MEM_stage_inst_dmem_n8016, MEM_stage_inst_dmem_n8015, MEM_stage_inst_dmem_n8014, MEM_stage_inst_dmem_n8013, MEM_stage_inst_dmem_n8012, MEM_stage_inst_dmem_n8011, MEM_stage_inst_dmem_n8010, MEM_stage_inst_dmem_n8009, MEM_stage_inst_dmem_n8008, MEM_stage_inst_dmem_n8007, MEM_stage_inst_dmem_n8006, MEM_stage_inst_dmem_n8005, MEM_stage_inst_dmem_n8004, MEM_stage_inst_dmem_n8003, MEM_stage_inst_dmem_n8002, MEM_stage_inst_dmem_n8001, MEM_stage_inst_dmem_n8000, MEM_stage_inst_dmem_n7999, MEM_stage_inst_dmem_n7998, MEM_stage_inst_dmem_n7997, MEM_stage_inst_dmem_n7996, MEM_stage_inst_dmem_n7995, MEM_stage_inst_dmem_n7994, MEM_stage_inst_dmem_n7993, MEM_stage_inst_dmem_n7992, MEM_stage_inst_dmem_n7991, MEM_stage_inst_dmem_n7990, MEM_stage_inst_dmem_n7989, MEM_stage_inst_dmem_n7988, MEM_stage_inst_dmem_n7987, MEM_stage_inst_dmem_n7986, MEM_stage_inst_dmem_n7985, MEM_stage_inst_dmem_n7984, MEM_stage_inst_dmem_n7983, MEM_stage_inst_dmem_n7982, MEM_stage_inst_dmem_n7981, MEM_stage_inst_dmem_n7980, MEM_stage_inst_dmem_n7979, MEM_stage_inst_dmem_n7978, MEM_stage_inst_dmem_n7977, MEM_stage_inst_dmem_n7976, MEM_stage_inst_dmem_n7975, MEM_stage_inst_dmem_n7974, MEM_stage_inst_dmem_n7973, MEM_stage_inst_dmem_n7972, MEM_stage_inst_dmem_n7971, MEM_stage_inst_dmem_n7970, MEM_stage_inst_dmem_n7969, MEM_stage_inst_dmem_n7968, MEM_stage_inst_dmem_n7967, MEM_stage_inst_dmem_n7966, MEM_stage_inst_dmem_n7965, MEM_stage_inst_dmem_n7964, MEM_stage_inst_dmem_n7963, MEM_stage_inst_dmem_n7962, MEM_stage_inst_dmem_n7961, MEM_stage_inst_dmem_n7960, MEM_stage_inst_dmem_n7959, MEM_stage_inst_dmem_n7958, MEM_stage_inst_dmem_n7957, MEM_stage_inst_dmem_n7956, MEM_stage_inst_dmem_n7955, MEM_stage_inst_dmem_n7954, MEM_stage_inst_dmem_n7953, MEM_stage_inst_dmem_n7952, MEM_stage_inst_dmem_n7951, MEM_stage_inst_dmem_n7950, MEM_stage_inst_dmem_n7949, MEM_stage_inst_dmem_n7948, MEM_stage_inst_dmem_n7947, MEM_stage_inst_dmem_n7946, MEM_stage_inst_dmem_n7945, MEM_stage_inst_dmem_n7944, MEM_stage_inst_dmem_n7943, MEM_stage_inst_dmem_n7942, MEM_stage_inst_dmem_n7941, MEM_stage_inst_dmem_n7940, MEM_stage_inst_dmem_n7939, MEM_stage_inst_dmem_n7938, MEM_stage_inst_dmem_n7937, MEM_stage_inst_dmem_n7936, MEM_stage_inst_dmem_n7935, MEM_stage_inst_dmem_n7934, MEM_stage_inst_dmem_n7933, MEM_stage_inst_dmem_n7932, MEM_stage_inst_dmem_n7931, MEM_stage_inst_dmem_n7930, MEM_stage_inst_dmem_n7929, MEM_stage_inst_dmem_n7928, MEM_stage_inst_dmem_n7927, MEM_stage_inst_dmem_n7926, MEM_stage_inst_dmem_n7925, MEM_stage_inst_dmem_n7924, MEM_stage_inst_dmem_n7923, MEM_stage_inst_dmem_n7922, MEM_stage_inst_dmem_n7921, MEM_stage_inst_dmem_n7920, MEM_stage_inst_dmem_n7919, MEM_stage_inst_dmem_n7918, MEM_stage_inst_dmem_n7917, MEM_stage_inst_dmem_n7916, MEM_stage_inst_dmem_n7915, MEM_stage_inst_dmem_n7914, MEM_stage_inst_dmem_n7913, MEM_stage_inst_dmem_n7912, MEM_stage_inst_dmem_n7911, MEM_stage_inst_dmem_n7910, MEM_stage_inst_dmem_n7909, MEM_stage_inst_dmem_n7908, MEM_stage_inst_dmem_n7907, MEM_stage_inst_dmem_n7906, MEM_stage_inst_dmem_n7905, MEM_stage_inst_dmem_n7904, MEM_stage_inst_dmem_n7903, MEM_stage_inst_dmem_n7902, MEM_stage_inst_dmem_n7901, MEM_stage_inst_dmem_n7900, MEM_stage_inst_dmem_n7899, MEM_stage_inst_dmem_n7898, MEM_stage_inst_dmem_n7897, MEM_stage_inst_dmem_n7896, MEM_stage_inst_dmem_n7895, MEM_stage_inst_dmem_n7894, MEM_stage_inst_dmem_n7893, MEM_stage_inst_dmem_n7892, MEM_stage_inst_dmem_n7891, MEM_stage_inst_dmem_n7890, MEM_stage_inst_dmem_n7889, MEM_stage_inst_dmem_n7888, MEM_stage_inst_dmem_n7887, MEM_stage_inst_dmem_n7886, MEM_stage_inst_dmem_n7885, MEM_stage_inst_dmem_n7884, MEM_stage_inst_dmem_n7883, MEM_stage_inst_dmem_n7882, MEM_stage_inst_dmem_n7881, MEM_stage_inst_dmem_n7880, MEM_stage_inst_dmem_n7879, MEM_stage_inst_dmem_n7878, MEM_stage_inst_dmem_n7877, MEM_stage_inst_dmem_n7876, MEM_stage_inst_dmem_n7875, MEM_stage_inst_dmem_n7874, MEM_stage_inst_dmem_n7873, MEM_stage_inst_dmem_n7872, MEM_stage_inst_dmem_n7871, MEM_stage_inst_dmem_n7870, MEM_stage_inst_dmem_n7869, MEM_stage_inst_dmem_n7868, MEM_stage_inst_dmem_n7867, MEM_stage_inst_dmem_n7866, MEM_stage_inst_dmem_n7865, MEM_stage_inst_dmem_n7864, MEM_stage_inst_dmem_n7863, MEM_stage_inst_dmem_n7862, MEM_stage_inst_dmem_n7861, MEM_stage_inst_dmem_n7860, MEM_stage_inst_dmem_n7859, MEM_stage_inst_dmem_n7858, MEM_stage_inst_dmem_n7857, MEM_stage_inst_dmem_n7856, MEM_stage_inst_dmem_n7855, MEM_stage_inst_dmem_n7854, MEM_stage_inst_dmem_n7853, MEM_stage_inst_dmem_n7852, MEM_stage_inst_dmem_n7851, MEM_stage_inst_dmem_n7850, MEM_stage_inst_dmem_n7849, MEM_stage_inst_dmem_n7848, MEM_stage_inst_dmem_n7847, MEM_stage_inst_dmem_n7846, MEM_stage_inst_dmem_n7845, MEM_stage_inst_dmem_n7844, MEM_stage_inst_dmem_n7843, MEM_stage_inst_dmem_n7842, MEM_stage_inst_dmem_n7841, MEM_stage_inst_dmem_n7840, MEM_stage_inst_dmem_n7839, MEM_stage_inst_dmem_n7838, MEM_stage_inst_dmem_n7837, MEM_stage_inst_dmem_n7836, MEM_stage_inst_dmem_n7835, MEM_stage_inst_dmem_n7834, MEM_stage_inst_dmem_n7833, MEM_stage_inst_dmem_n7832, MEM_stage_inst_dmem_n7831, MEM_stage_inst_dmem_n7830, MEM_stage_inst_dmem_n7829, MEM_stage_inst_dmem_n7828, MEM_stage_inst_dmem_n7827, MEM_stage_inst_dmem_n7826, MEM_stage_inst_dmem_n7825, MEM_stage_inst_dmem_n7824, MEM_stage_inst_dmem_n7823, MEM_stage_inst_dmem_n7822, MEM_stage_inst_dmem_n7821, MEM_stage_inst_dmem_n7820, MEM_stage_inst_dmem_n7819, MEM_stage_inst_dmem_n7818, MEM_stage_inst_dmem_n7817, MEM_stage_inst_dmem_n7816, MEM_stage_inst_dmem_n7815, MEM_stage_inst_dmem_n7814, MEM_stage_inst_dmem_n7813, MEM_stage_inst_dmem_n7812, MEM_stage_inst_dmem_n7811, MEM_stage_inst_dmem_n7810, MEM_stage_inst_dmem_n7809, MEM_stage_inst_dmem_n7808, MEM_stage_inst_dmem_n7807, MEM_stage_inst_dmem_n7806, MEM_stage_inst_dmem_n7805, MEM_stage_inst_dmem_n7804, MEM_stage_inst_dmem_n7803, MEM_stage_inst_dmem_n7802, MEM_stage_inst_dmem_n7801, MEM_stage_inst_dmem_n7800, MEM_stage_inst_dmem_n7799, MEM_stage_inst_dmem_n7798, MEM_stage_inst_dmem_n7797, MEM_stage_inst_dmem_n7796, MEM_stage_inst_dmem_n7795, MEM_stage_inst_dmem_n7794, MEM_stage_inst_dmem_n7793, MEM_stage_inst_dmem_n7792, MEM_stage_inst_dmem_n7791, MEM_stage_inst_dmem_n7790, MEM_stage_inst_dmem_n7789, MEM_stage_inst_dmem_n7788, MEM_stage_inst_dmem_n7787, MEM_stage_inst_dmem_n7786, MEM_stage_inst_dmem_n7785, MEM_stage_inst_dmem_n7784, MEM_stage_inst_dmem_n7783, MEM_stage_inst_dmem_n7782, MEM_stage_inst_dmem_n7781, MEM_stage_inst_dmem_n7780, MEM_stage_inst_dmem_n7779, MEM_stage_inst_dmem_n7778, MEM_stage_inst_dmem_n7777, MEM_stage_inst_dmem_n7776, MEM_stage_inst_dmem_n7775, MEM_stage_inst_dmem_n7774, MEM_stage_inst_dmem_n7773, MEM_stage_inst_dmem_n7772, MEM_stage_inst_dmem_n7771, MEM_stage_inst_dmem_n7770, MEM_stage_inst_dmem_n7769, MEM_stage_inst_dmem_n7768, MEM_stage_inst_dmem_n7767, MEM_stage_inst_dmem_n7766, MEM_stage_inst_dmem_n7765, MEM_stage_inst_dmem_n7764, MEM_stage_inst_dmem_n7763, MEM_stage_inst_dmem_n7762, MEM_stage_inst_dmem_n7761, MEM_stage_inst_dmem_n7760, MEM_stage_inst_dmem_n7759, MEM_stage_inst_dmem_n7758, MEM_stage_inst_dmem_n7757, MEM_stage_inst_dmem_n7756, MEM_stage_inst_dmem_n7755, MEM_stage_inst_dmem_n7754, MEM_stage_inst_dmem_n7753, MEM_stage_inst_dmem_n7752, MEM_stage_inst_dmem_n7751, MEM_stage_inst_dmem_n7750, MEM_stage_inst_dmem_n7749, MEM_stage_inst_dmem_n7748, MEM_stage_inst_dmem_n7747, MEM_stage_inst_dmem_n7746, MEM_stage_inst_dmem_n7745, MEM_stage_inst_dmem_n7744, MEM_stage_inst_dmem_n7743, MEM_stage_inst_dmem_n7742, MEM_stage_inst_dmem_n7741, MEM_stage_inst_dmem_n7740, MEM_stage_inst_dmem_n7739, MEM_stage_inst_dmem_n7738, MEM_stage_inst_dmem_n7737, MEM_stage_inst_dmem_n7736, MEM_stage_inst_dmem_n7735, MEM_stage_inst_dmem_n7734, MEM_stage_inst_dmem_n7733, MEM_stage_inst_dmem_n7732, MEM_stage_inst_dmem_n7731, MEM_stage_inst_dmem_n7730, MEM_stage_inst_dmem_n7729, MEM_stage_inst_dmem_n7728, MEM_stage_inst_dmem_n7727, MEM_stage_inst_dmem_n7726, MEM_stage_inst_dmem_n7725, MEM_stage_inst_dmem_n7724, MEM_stage_inst_dmem_n7723, MEM_stage_inst_dmem_n7722, MEM_stage_inst_dmem_n7721, MEM_stage_inst_dmem_n7720, MEM_stage_inst_dmem_n7719, MEM_stage_inst_dmem_n7718, MEM_stage_inst_dmem_n7717, MEM_stage_inst_dmem_n7716, MEM_stage_inst_dmem_n7715, MEM_stage_inst_dmem_n7714, MEM_stage_inst_dmem_n7713, MEM_stage_inst_dmem_n7712, MEM_stage_inst_dmem_n7711, MEM_stage_inst_dmem_n7710, MEM_stage_inst_dmem_n7709, MEM_stage_inst_dmem_n7708, MEM_stage_inst_dmem_n7707, MEM_stage_inst_dmem_n7706, MEM_stage_inst_dmem_n7705, MEM_stage_inst_dmem_n7704, MEM_stage_inst_dmem_n7703, MEM_stage_inst_dmem_n7702, MEM_stage_inst_dmem_n7701, MEM_stage_inst_dmem_n7700, MEM_stage_inst_dmem_n7699, MEM_stage_inst_dmem_n7698, MEM_stage_inst_dmem_n7697, MEM_stage_inst_dmem_n7696, MEM_stage_inst_dmem_n7695, MEM_stage_inst_dmem_n7694, MEM_stage_inst_dmem_n7693, MEM_stage_inst_dmem_n7692, MEM_stage_inst_dmem_n7691, MEM_stage_inst_dmem_n7690, MEM_stage_inst_dmem_n7689, MEM_stage_inst_dmem_n7688, MEM_stage_inst_dmem_n7687, MEM_stage_inst_dmem_n7686, MEM_stage_inst_dmem_n7685, MEM_stage_inst_dmem_n7684, MEM_stage_inst_dmem_n7683, MEM_stage_inst_dmem_n7682, MEM_stage_inst_dmem_n7681, MEM_stage_inst_dmem_n7680, MEM_stage_inst_dmem_n7679, MEM_stage_inst_dmem_n7678, MEM_stage_inst_dmem_n7677, MEM_stage_inst_dmem_n7676, MEM_stage_inst_dmem_n7675, MEM_stage_inst_dmem_n7674, MEM_stage_inst_dmem_n7673, MEM_stage_inst_dmem_n7672, MEM_stage_inst_dmem_n7671, MEM_stage_inst_dmem_n7670, MEM_stage_inst_dmem_n7669, MEM_stage_inst_dmem_n7668, MEM_stage_inst_dmem_n7667, MEM_stage_inst_dmem_n7666, MEM_stage_inst_dmem_n7665, MEM_stage_inst_dmem_n7664, MEM_stage_inst_dmem_n7663, MEM_stage_inst_dmem_n7662, MEM_stage_inst_dmem_n7661, MEM_stage_inst_dmem_n7660, MEM_stage_inst_dmem_n7659, MEM_stage_inst_dmem_n7658, MEM_stage_inst_dmem_n7657, MEM_stage_inst_dmem_n7656, MEM_stage_inst_dmem_n7655, MEM_stage_inst_dmem_n7654, MEM_stage_inst_dmem_n7653, MEM_stage_inst_dmem_n7652, MEM_stage_inst_dmem_n7651, MEM_stage_inst_dmem_n7650, MEM_stage_inst_dmem_n7649, MEM_stage_inst_dmem_n7648, MEM_stage_inst_dmem_n7647, MEM_stage_inst_dmem_n7646, MEM_stage_inst_dmem_n7645, MEM_stage_inst_dmem_n7644, MEM_stage_inst_dmem_n7643, MEM_stage_inst_dmem_n7642, MEM_stage_inst_dmem_n7641, MEM_stage_inst_dmem_n7640, MEM_stage_inst_dmem_n7639, MEM_stage_inst_dmem_n7638, MEM_stage_inst_dmem_n7637, MEM_stage_inst_dmem_n7636, MEM_stage_inst_dmem_n7635, MEM_stage_inst_dmem_n7634, MEM_stage_inst_dmem_n7633, MEM_stage_inst_dmem_n7632, MEM_stage_inst_dmem_n7631, MEM_stage_inst_dmem_n7630, MEM_stage_inst_dmem_n7629, MEM_stage_inst_dmem_n7628, MEM_stage_inst_dmem_n7627, MEM_stage_inst_dmem_n7626, MEM_stage_inst_dmem_n7625, MEM_stage_inst_dmem_n7624, MEM_stage_inst_dmem_n7623, MEM_stage_inst_dmem_n7622, MEM_stage_inst_dmem_n7621, MEM_stage_inst_dmem_n7620, MEM_stage_inst_dmem_n7619, MEM_stage_inst_dmem_n7618, MEM_stage_inst_dmem_n7617, MEM_stage_inst_dmem_n7616, MEM_stage_inst_dmem_n7615, MEM_stage_inst_dmem_n7614, MEM_stage_inst_dmem_n7613, MEM_stage_inst_dmem_n7612, MEM_stage_inst_dmem_n7611, MEM_stage_inst_dmem_n7610, MEM_stage_inst_dmem_n7609, MEM_stage_inst_dmem_n7608, MEM_stage_inst_dmem_n7607, MEM_stage_inst_dmem_n7606, MEM_stage_inst_dmem_n7605, MEM_stage_inst_dmem_n7604, MEM_stage_inst_dmem_n7603, MEM_stage_inst_dmem_n7602, MEM_stage_inst_dmem_n7601, MEM_stage_inst_dmem_n7600, MEM_stage_inst_dmem_n7599, MEM_stage_inst_dmem_n7598, MEM_stage_inst_dmem_n7597, MEM_stage_inst_dmem_n7596, MEM_stage_inst_dmem_n7595, MEM_stage_inst_dmem_n7594, MEM_stage_inst_dmem_n7593, MEM_stage_inst_dmem_n7592, MEM_stage_inst_dmem_n7591, MEM_stage_inst_dmem_n7590, MEM_stage_inst_dmem_n7589, MEM_stage_inst_dmem_n7588, MEM_stage_inst_dmem_n7587, MEM_stage_inst_dmem_n7586, MEM_stage_inst_dmem_n7585, MEM_stage_inst_dmem_n7584, MEM_stage_inst_dmem_n7583, MEM_stage_inst_dmem_n7582, MEM_stage_inst_dmem_n7581, MEM_stage_inst_dmem_n7580, MEM_stage_inst_dmem_n7579, MEM_stage_inst_dmem_n7578, MEM_stage_inst_dmem_n7577, MEM_stage_inst_dmem_n7576, MEM_stage_inst_dmem_n7575, MEM_stage_inst_dmem_n7574, MEM_stage_inst_dmem_n7573, MEM_stage_inst_dmem_n7572, MEM_stage_inst_dmem_n7571, MEM_stage_inst_dmem_n7570, MEM_stage_inst_dmem_n7569, MEM_stage_inst_dmem_n7568, MEM_stage_inst_dmem_n7567, MEM_stage_inst_dmem_n7566, MEM_stage_inst_dmem_n7565, MEM_stage_inst_dmem_n7564, MEM_stage_inst_dmem_n7563, MEM_stage_inst_dmem_n7562, MEM_stage_inst_dmem_n7561, MEM_stage_inst_dmem_n7560, MEM_stage_inst_dmem_n7559, MEM_stage_inst_dmem_n7558, MEM_stage_inst_dmem_n7557, MEM_stage_inst_dmem_n7556, MEM_stage_inst_dmem_n7555, MEM_stage_inst_dmem_n7554, MEM_stage_inst_dmem_n7553, MEM_stage_inst_dmem_n7552, MEM_stage_inst_dmem_n7551, MEM_stage_inst_dmem_n7550, MEM_stage_inst_dmem_n7549, MEM_stage_inst_dmem_n7548, MEM_stage_inst_dmem_n7547, MEM_stage_inst_dmem_n7546, MEM_stage_inst_dmem_n7545, MEM_stage_inst_dmem_n7544, MEM_stage_inst_dmem_n7543, MEM_stage_inst_dmem_n7542, MEM_stage_inst_dmem_n7541, MEM_stage_inst_dmem_n7540, MEM_stage_inst_dmem_n7539, MEM_stage_inst_dmem_n7538, MEM_stage_inst_dmem_n7537, MEM_stage_inst_dmem_n7536, MEM_stage_inst_dmem_n7535, MEM_stage_inst_dmem_n7534, MEM_stage_inst_dmem_n7533, MEM_stage_inst_dmem_n7532, MEM_stage_inst_dmem_n7531, MEM_stage_inst_dmem_n7530, MEM_stage_inst_dmem_n7529, MEM_stage_inst_dmem_n7528, MEM_stage_inst_dmem_n7527, MEM_stage_inst_dmem_n7526, MEM_stage_inst_dmem_n7525, MEM_stage_inst_dmem_n7524, MEM_stage_inst_dmem_n7523, MEM_stage_inst_dmem_n7522, MEM_stage_inst_dmem_n7521, MEM_stage_inst_dmem_n7520, MEM_stage_inst_dmem_n7519, MEM_stage_inst_dmem_n7518, MEM_stage_inst_dmem_n7517, MEM_stage_inst_dmem_n7516, MEM_stage_inst_dmem_n7515, MEM_stage_inst_dmem_n7514, MEM_stage_inst_dmem_n7513, MEM_stage_inst_dmem_n7512, MEM_stage_inst_dmem_n7511, MEM_stage_inst_dmem_n7510, MEM_stage_inst_dmem_n7509, MEM_stage_inst_dmem_n7508, MEM_stage_inst_dmem_n7507, MEM_stage_inst_dmem_n7506, MEM_stage_inst_dmem_n7505, MEM_stage_inst_dmem_n7504, MEM_stage_inst_dmem_n7503, MEM_stage_inst_dmem_n7502, MEM_stage_inst_dmem_n7501, MEM_stage_inst_dmem_n7500, MEM_stage_inst_dmem_n7499, MEM_stage_inst_dmem_n7498, MEM_stage_inst_dmem_n7497, MEM_stage_inst_dmem_n7496, MEM_stage_inst_dmem_n7495, MEM_stage_inst_dmem_n7494, MEM_stage_inst_dmem_n7493, MEM_stage_inst_dmem_n7492, MEM_stage_inst_dmem_n7491, MEM_stage_inst_dmem_n7490, MEM_stage_inst_dmem_n7489, MEM_stage_inst_dmem_n7488, MEM_stage_inst_dmem_n7487, MEM_stage_inst_dmem_n7486, MEM_stage_inst_dmem_n7485, MEM_stage_inst_dmem_n7484, MEM_stage_inst_dmem_n7483, MEM_stage_inst_dmem_n7482, MEM_stage_inst_dmem_n7481, MEM_stage_inst_dmem_n7480, MEM_stage_inst_dmem_n7479, MEM_stage_inst_dmem_n7478, MEM_stage_inst_dmem_n7477, MEM_stage_inst_dmem_n7476, MEM_stage_inst_dmem_n7475, MEM_stage_inst_dmem_n7474, MEM_stage_inst_dmem_n7473, MEM_stage_inst_dmem_n7472, MEM_stage_inst_dmem_n7471, MEM_stage_inst_dmem_n7470, MEM_stage_inst_dmem_n7469, MEM_stage_inst_dmem_n7468, MEM_stage_inst_dmem_n7467, MEM_stage_inst_dmem_n7466, MEM_stage_inst_dmem_n7465, MEM_stage_inst_dmem_n7464, MEM_stage_inst_dmem_n7463, MEM_stage_inst_dmem_n7462, MEM_stage_inst_dmem_n7461, MEM_stage_inst_dmem_n7460, MEM_stage_inst_dmem_n7459, MEM_stage_inst_dmem_n7458, MEM_stage_inst_dmem_n7457, MEM_stage_inst_dmem_n7456, MEM_stage_inst_dmem_n7455, MEM_stage_inst_dmem_n7454, MEM_stage_inst_dmem_n7453, MEM_stage_inst_dmem_n7452, MEM_stage_inst_dmem_n7451, MEM_stage_inst_dmem_n7450, MEM_stage_inst_dmem_n7449, MEM_stage_inst_dmem_n7448, MEM_stage_inst_dmem_n7447, MEM_stage_inst_dmem_n7446, MEM_stage_inst_dmem_n7445, MEM_stage_inst_dmem_n7444, MEM_stage_inst_dmem_n7443, MEM_stage_inst_dmem_n7442, MEM_stage_inst_dmem_n7441, MEM_stage_inst_dmem_n7440, MEM_stage_inst_dmem_n7439, MEM_stage_inst_dmem_n7438, MEM_stage_inst_dmem_n7437, MEM_stage_inst_dmem_n7436, MEM_stage_inst_dmem_n7435, MEM_stage_inst_dmem_n7434, MEM_stage_inst_dmem_n7433, MEM_stage_inst_dmem_n7432, MEM_stage_inst_dmem_n7431, MEM_stage_inst_dmem_n7430, MEM_stage_inst_dmem_n7429, MEM_stage_inst_dmem_n7428, MEM_stage_inst_dmem_n7427, MEM_stage_inst_dmem_n7426, MEM_stage_inst_dmem_n7425, MEM_stage_inst_dmem_n7424, MEM_stage_inst_dmem_n7423, MEM_stage_inst_dmem_n7422, MEM_stage_inst_dmem_n7421, MEM_stage_inst_dmem_n7420, MEM_stage_inst_dmem_n7419, MEM_stage_inst_dmem_n7418, MEM_stage_inst_dmem_n7417, MEM_stage_inst_dmem_n7416, MEM_stage_inst_dmem_n7415, MEM_stage_inst_dmem_n7414, MEM_stage_inst_dmem_n7413, MEM_stage_inst_dmem_n7412, MEM_stage_inst_dmem_n7411, MEM_stage_inst_dmem_n7410, MEM_stage_inst_dmem_n7409, MEM_stage_inst_dmem_n7408, MEM_stage_inst_dmem_n7407, MEM_stage_inst_dmem_n7406, MEM_stage_inst_dmem_n7405, MEM_stage_inst_dmem_n7404, MEM_stage_inst_dmem_n7403, MEM_stage_inst_dmem_n7402, MEM_stage_inst_dmem_n7401, MEM_stage_inst_dmem_n7400, MEM_stage_inst_dmem_n7399, MEM_stage_inst_dmem_n7398, MEM_stage_inst_dmem_n7397, MEM_stage_inst_dmem_n7396, MEM_stage_inst_dmem_n7395, MEM_stage_inst_dmem_n7394, MEM_stage_inst_dmem_n7393, MEM_stage_inst_dmem_n7392, MEM_stage_inst_dmem_n7391, MEM_stage_inst_dmem_n7390, MEM_stage_inst_dmem_n7389, MEM_stage_inst_dmem_n7388, MEM_stage_inst_dmem_n7387, MEM_stage_inst_dmem_n7386, MEM_stage_inst_dmem_n7385, MEM_stage_inst_dmem_n7384, MEM_stage_inst_dmem_n7383, MEM_stage_inst_dmem_n7382, MEM_stage_inst_dmem_n7381, MEM_stage_inst_dmem_n7380, MEM_stage_inst_dmem_n7379, MEM_stage_inst_dmem_n7378, MEM_stage_inst_dmem_n7377, MEM_stage_inst_dmem_n7376, MEM_stage_inst_dmem_n7375, MEM_stage_inst_dmem_n7374, MEM_stage_inst_dmem_n7373, MEM_stage_inst_dmem_n7372, MEM_stage_inst_dmem_n7371, MEM_stage_inst_dmem_n7370, MEM_stage_inst_dmem_n7369, MEM_stage_inst_dmem_n7368, MEM_stage_inst_dmem_n7367, MEM_stage_inst_dmem_n7366, MEM_stage_inst_dmem_n7365, MEM_stage_inst_dmem_n7364, MEM_stage_inst_dmem_n7363, MEM_stage_inst_dmem_n7362, MEM_stage_inst_dmem_n7361, MEM_stage_inst_dmem_n7360, MEM_stage_inst_dmem_n7359, MEM_stage_inst_dmem_n7358, MEM_stage_inst_dmem_n7357, MEM_stage_inst_dmem_n7356, MEM_stage_inst_dmem_n7355, MEM_stage_inst_dmem_n7354, MEM_stage_inst_dmem_n7353, MEM_stage_inst_dmem_n7352, MEM_stage_inst_dmem_n7351, MEM_stage_inst_dmem_n7350, MEM_stage_inst_dmem_n7349, MEM_stage_inst_dmem_n7348, MEM_stage_inst_dmem_n7347, MEM_stage_inst_dmem_n7346, MEM_stage_inst_dmem_n7345, MEM_stage_inst_dmem_n7344, MEM_stage_inst_dmem_n7343, MEM_stage_inst_dmem_n7342, MEM_stage_inst_dmem_n7341, MEM_stage_inst_dmem_n7340, MEM_stage_inst_dmem_n7339, MEM_stage_inst_dmem_n7338, MEM_stage_inst_dmem_n7337, MEM_stage_inst_dmem_n7336, MEM_stage_inst_dmem_n7335, MEM_stage_inst_dmem_n7334, MEM_stage_inst_dmem_n7333, MEM_stage_inst_dmem_n7332, MEM_stage_inst_dmem_n7331, MEM_stage_inst_dmem_n7330, MEM_stage_inst_dmem_n7329, MEM_stage_inst_dmem_n7328, MEM_stage_inst_dmem_n7327, MEM_stage_inst_dmem_n7326, MEM_stage_inst_dmem_n7325, MEM_stage_inst_dmem_n7324, MEM_stage_inst_dmem_n7323, MEM_stage_inst_dmem_n7322, MEM_stage_inst_dmem_n7321, MEM_stage_inst_dmem_n7320, MEM_stage_inst_dmem_n7319, MEM_stage_inst_dmem_n7318, MEM_stage_inst_dmem_n7317, MEM_stage_inst_dmem_n7316, MEM_stage_inst_dmem_n7315, MEM_stage_inst_dmem_n7314, MEM_stage_inst_dmem_n7313, MEM_stage_inst_dmem_n7312, MEM_stage_inst_dmem_n7311, MEM_stage_inst_dmem_n7310, MEM_stage_inst_dmem_n7309, MEM_stage_inst_dmem_n7308, MEM_stage_inst_dmem_n7307, MEM_stage_inst_dmem_n7306, MEM_stage_inst_dmem_n7305, MEM_stage_inst_dmem_n7304, MEM_stage_inst_dmem_n7303, MEM_stage_inst_dmem_n7302, MEM_stage_inst_dmem_n7301, MEM_stage_inst_dmem_n7300, MEM_stage_inst_dmem_n7299, MEM_stage_inst_dmem_n7298, MEM_stage_inst_dmem_n7297, MEM_stage_inst_dmem_n7296, MEM_stage_inst_dmem_n7295, MEM_stage_inst_dmem_n7294, MEM_stage_inst_dmem_n7293, MEM_stage_inst_dmem_n7292, MEM_stage_inst_dmem_n7291, MEM_stage_inst_dmem_n7290, MEM_stage_inst_dmem_n7289, MEM_stage_inst_dmem_n7288, MEM_stage_inst_dmem_n7287, MEM_stage_inst_dmem_n7286, MEM_stage_inst_dmem_n7285, MEM_stage_inst_dmem_n7284, MEM_stage_inst_dmem_n7283, MEM_stage_inst_dmem_n7282, MEM_stage_inst_dmem_n7281, MEM_stage_inst_dmem_n7280, MEM_stage_inst_dmem_n7279, MEM_stage_inst_dmem_n7278, MEM_stage_inst_dmem_n7277, MEM_stage_inst_dmem_n7276, MEM_stage_inst_dmem_n7275, MEM_stage_inst_dmem_n7274, MEM_stage_inst_dmem_n7273, MEM_stage_inst_dmem_n7272, MEM_stage_inst_dmem_n7271, MEM_stage_inst_dmem_n7270, MEM_stage_inst_dmem_n7269, MEM_stage_inst_dmem_n7268, MEM_stage_inst_dmem_n7267, MEM_stage_inst_dmem_n7266, MEM_stage_inst_dmem_n7265, MEM_stage_inst_dmem_n7264, MEM_stage_inst_dmem_n7263, MEM_stage_inst_dmem_n7262, MEM_stage_inst_dmem_n7261, MEM_stage_inst_dmem_n7260, MEM_stage_inst_dmem_n7259, MEM_stage_inst_dmem_n7258, MEM_stage_inst_dmem_n7257, MEM_stage_inst_dmem_n7256, MEM_stage_inst_dmem_n7255, MEM_stage_inst_dmem_n7254, MEM_stage_inst_dmem_n7253, MEM_stage_inst_dmem_n7252, MEM_stage_inst_dmem_n7251, MEM_stage_inst_dmem_n7250, MEM_stage_inst_dmem_n7249, MEM_stage_inst_dmem_n7248, MEM_stage_inst_dmem_n7247, MEM_stage_inst_dmem_n7246, MEM_stage_inst_dmem_n7245, MEM_stage_inst_dmem_n7244, MEM_stage_inst_dmem_n7243, MEM_stage_inst_dmem_n7242, MEM_stage_inst_dmem_n7241, MEM_stage_inst_dmem_n7240, MEM_stage_inst_dmem_n7239, MEM_stage_inst_dmem_n7238, MEM_stage_inst_dmem_n7237, MEM_stage_inst_dmem_n7236, MEM_stage_inst_dmem_n7235, MEM_stage_inst_dmem_n7234, MEM_stage_inst_dmem_n7233, MEM_stage_inst_dmem_n7232, MEM_stage_inst_dmem_n7231, MEM_stage_inst_dmem_n7230, MEM_stage_inst_dmem_n7229, MEM_stage_inst_dmem_n7228, MEM_stage_inst_dmem_n7227, MEM_stage_inst_dmem_n7226, MEM_stage_inst_dmem_n7225, MEM_stage_inst_dmem_n7224, MEM_stage_inst_dmem_n7223, MEM_stage_inst_dmem_n7222, MEM_stage_inst_dmem_n7221, MEM_stage_inst_dmem_n7220, MEM_stage_inst_dmem_n7219, MEM_stage_inst_dmem_n7218, MEM_stage_inst_dmem_n7217, MEM_stage_inst_dmem_n7216, MEM_stage_inst_dmem_n7215, MEM_stage_inst_dmem_n7214, MEM_stage_inst_dmem_n7213, MEM_stage_inst_dmem_n7212, MEM_stage_inst_dmem_n7211, MEM_stage_inst_dmem_n7210, MEM_stage_inst_dmem_n7209, MEM_stage_inst_dmem_n7208, MEM_stage_inst_dmem_n7207, MEM_stage_inst_dmem_n7206, MEM_stage_inst_dmem_n7205, MEM_stage_inst_dmem_n7204, MEM_stage_inst_dmem_n7203, MEM_stage_inst_dmem_n7202, MEM_stage_inst_dmem_n7201, MEM_stage_inst_dmem_n7200, MEM_stage_inst_dmem_n7199, MEM_stage_inst_dmem_n7198, MEM_stage_inst_dmem_n7197, MEM_stage_inst_dmem_n7196, MEM_stage_inst_dmem_n7195, MEM_stage_inst_dmem_n7194, MEM_stage_inst_dmem_n7193, MEM_stage_inst_dmem_n7192, MEM_stage_inst_dmem_n7191, MEM_stage_inst_dmem_n7190, MEM_stage_inst_dmem_n7189, MEM_stage_inst_dmem_n7188, MEM_stage_inst_dmem_n7187, MEM_stage_inst_dmem_n7186, MEM_stage_inst_dmem_n7185, MEM_stage_inst_dmem_n7184, MEM_stage_inst_dmem_n7183, MEM_stage_inst_dmem_n7182, MEM_stage_inst_dmem_n7181, MEM_stage_inst_dmem_n7180, MEM_stage_inst_dmem_n7179, MEM_stage_inst_dmem_n7178, MEM_stage_inst_dmem_n7177, MEM_stage_inst_dmem_n7176, MEM_stage_inst_dmem_n7175, MEM_stage_inst_dmem_n7174, MEM_stage_inst_dmem_n7173, MEM_stage_inst_dmem_n7172, MEM_stage_inst_dmem_n7171, MEM_stage_inst_dmem_n7170, MEM_stage_inst_dmem_n7169, MEM_stage_inst_dmem_n7168, MEM_stage_inst_dmem_n7167, MEM_stage_inst_dmem_n7166, MEM_stage_inst_dmem_n7165, MEM_stage_inst_dmem_n7164, MEM_stage_inst_dmem_n7163, MEM_stage_inst_dmem_n7162, MEM_stage_inst_dmem_n7161, MEM_stage_inst_dmem_n7160, MEM_stage_inst_dmem_n7159, MEM_stage_inst_dmem_n7158, MEM_stage_inst_dmem_n7157, MEM_stage_inst_dmem_n7156, MEM_stage_inst_dmem_n7155, MEM_stage_inst_dmem_n7154, MEM_stage_inst_dmem_n7153, MEM_stage_inst_dmem_n7152, MEM_stage_inst_dmem_n7151, MEM_stage_inst_dmem_n7150, MEM_stage_inst_dmem_n7149, MEM_stage_inst_dmem_n7148, MEM_stage_inst_dmem_n7147, MEM_stage_inst_dmem_n7146, MEM_stage_inst_dmem_n7145, MEM_stage_inst_dmem_n7144, MEM_stage_inst_dmem_n7143, MEM_stage_inst_dmem_n7142, MEM_stage_inst_dmem_n7141, MEM_stage_inst_dmem_n7140, MEM_stage_inst_dmem_n7139, MEM_stage_inst_dmem_n7138, MEM_stage_inst_dmem_n7137, MEM_stage_inst_dmem_n7136, MEM_stage_inst_dmem_n7135, MEM_stage_inst_dmem_n7134, MEM_stage_inst_dmem_n7133, MEM_stage_inst_dmem_n7132, MEM_stage_inst_dmem_n7131, MEM_stage_inst_dmem_n7130, MEM_stage_inst_dmem_n7129, MEM_stage_inst_dmem_n7128, MEM_stage_inst_dmem_n7127, MEM_stage_inst_dmem_n7126, MEM_stage_inst_dmem_n7125, MEM_stage_inst_dmem_n7124, MEM_stage_inst_dmem_n7123, MEM_stage_inst_dmem_n7122, MEM_stage_inst_dmem_n7121, MEM_stage_inst_dmem_n7120, MEM_stage_inst_dmem_n7119, MEM_stage_inst_dmem_n7118, MEM_stage_inst_dmem_n7117, MEM_stage_inst_dmem_n7116, MEM_stage_inst_dmem_n7115, MEM_stage_inst_dmem_n7114, MEM_stage_inst_dmem_n7113, MEM_stage_inst_dmem_n7112, MEM_stage_inst_dmem_n7111, MEM_stage_inst_dmem_n7110, MEM_stage_inst_dmem_n7109, MEM_stage_inst_dmem_n7108, MEM_stage_inst_dmem_n7107, MEM_stage_inst_dmem_n7106, MEM_stage_inst_dmem_n7105, MEM_stage_inst_dmem_n7104, MEM_stage_inst_dmem_n7103, MEM_stage_inst_dmem_n7102, MEM_stage_inst_dmem_n7101, MEM_stage_inst_dmem_n7100, MEM_stage_inst_dmem_n7099, MEM_stage_inst_dmem_n7098, MEM_stage_inst_dmem_n7097, MEM_stage_inst_dmem_n7096, MEM_stage_inst_dmem_n7095, MEM_stage_inst_dmem_n7094, MEM_stage_inst_dmem_n7093, MEM_stage_inst_dmem_n7092, MEM_stage_inst_dmem_n7091, MEM_stage_inst_dmem_n7090, MEM_stage_inst_dmem_n7089, MEM_stage_inst_dmem_n7088, MEM_stage_inst_dmem_n7087, MEM_stage_inst_dmem_n7086, MEM_stage_inst_dmem_n7085, MEM_stage_inst_dmem_n7084, MEM_stage_inst_dmem_n7083, MEM_stage_inst_dmem_n7082, MEM_stage_inst_dmem_n7081, MEM_stage_inst_dmem_n7080, MEM_stage_inst_dmem_n7079, MEM_stage_inst_dmem_n7078, MEM_stage_inst_dmem_n7077, MEM_stage_inst_dmem_n7076, MEM_stage_inst_dmem_n7075, MEM_stage_inst_dmem_n7074, MEM_stage_inst_dmem_n7073, MEM_stage_inst_dmem_n7072, MEM_stage_inst_dmem_n7071, MEM_stage_inst_dmem_n7070, MEM_stage_inst_dmem_n7069, MEM_stage_inst_dmem_n7068, MEM_stage_inst_dmem_n7067, MEM_stage_inst_dmem_n7066, MEM_stage_inst_dmem_n7065, MEM_stage_inst_dmem_n7064, MEM_stage_inst_dmem_n7063, MEM_stage_inst_dmem_n7062, MEM_stage_inst_dmem_n7061, MEM_stage_inst_dmem_n7060, MEM_stage_inst_dmem_n7059, MEM_stage_inst_dmem_n7058, MEM_stage_inst_dmem_n7057, MEM_stage_inst_dmem_n7056, MEM_stage_inst_dmem_n7055, MEM_stage_inst_dmem_n7054, MEM_stage_inst_dmem_n7053, MEM_stage_inst_dmem_n7052, MEM_stage_inst_dmem_n7051, MEM_stage_inst_dmem_n7050, MEM_stage_inst_dmem_n7049, MEM_stage_inst_dmem_n7048, MEM_stage_inst_dmem_n7047, MEM_stage_inst_dmem_n7046, MEM_stage_inst_dmem_n7045, MEM_stage_inst_dmem_n7044, MEM_stage_inst_dmem_n7043, MEM_stage_inst_dmem_n7042, MEM_stage_inst_dmem_n7041, MEM_stage_inst_dmem_n7040, MEM_stage_inst_dmem_n7039, MEM_stage_inst_dmem_n7038, MEM_stage_inst_dmem_n7037, MEM_stage_inst_dmem_n7036, MEM_stage_inst_dmem_n7035, MEM_stage_inst_dmem_n7034, MEM_stage_inst_dmem_n7033, MEM_stage_inst_dmem_n7032, MEM_stage_inst_dmem_n7031, MEM_stage_inst_dmem_n7030, MEM_stage_inst_dmem_n7029, MEM_stage_inst_dmem_n7028, MEM_stage_inst_dmem_n7027, MEM_stage_inst_dmem_n7026, MEM_stage_inst_dmem_n7025, MEM_stage_inst_dmem_n7024, MEM_stage_inst_dmem_n7023, MEM_stage_inst_dmem_n7022, MEM_stage_inst_dmem_n7021, MEM_stage_inst_dmem_n7020, MEM_stage_inst_dmem_n7019, MEM_stage_inst_dmem_n7018, MEM_stage_inst_dmem_n7017, MEM_stage_inst_dmem_n7016, MEM_stage_inst_dmem_n7015, MEM_stage_inst_dmem_n7014, MEM_stage_inst_dmem_n7013, MEM_stage_inst_dmem_n7012, MEM_stage_inst_dmem_n7011, MEM_stage_inst_dmem_n7010, MEM_stage_inst_dmem_n7009, MEM_stage_inst_dmem_n7008, MEM_stage_inst_dmem_n7007, MEM_stage_inst_dmem_n7006, MEM_stage_inst_dmem_n7005, MEM_stage_inst_dmem_n7004, MEM_stage_inst_dmem_n7003, MEM_stage_inst_dmem_n7002, MEM_stage_inst_dmem_n7001, MEM_stage_inst_dmem_n7000, MEM_stage_inst_dmem_n6999, MEM_stage_inst_dmem_n6998, MEM_stage_inst_dmem_n6997, MEM_stage_inst_dmem_n6996, MEM_stage_inst_dmem_n6995, MEM_stage_inst_dmem_n6994, MEM_stage_inst_dmem_n6993, MEM_stage_inst_dmem_n6992, MEM_stage_inst_dmem_n6991, MEM_stage_inst_dmem_n6990, MEM_stage_inst_dmem_n6989, MEM_stage_inst_dmem_n6988, MEM_stage_inst_dmem_n6987, MEM_stage_inst_dmem_n6986, MEM_stage_inst_dmem_n6985, MEM_stage_inst_dmem_n6984, MEM_stage_inst_dmem_n6983, MEM_stage_inst_dmem_n6982, MEM_stage_inst_dmem_n6981, MEM_stage_inst_dmem_n6980, MEM_stage_inst_dmem_n6979, MEM_stage_inst_dmem_n6978, MEM_stage_inst_dmem_n6977, MEM_stage_inst_dmem_n6976, MEM_stage_inst_dmem_n6975, MEM_stage_inst_dmem_n6974, MEM_stage_inst_dmem_n6973, MEM_stage_inst_dmem_n6972, MEM_stage_inst_dmem_n6971, MEM_stage_inst_dmem_n6970, MEM_stage_inst_dmem_n6969, MEM_stage_inst_dmem_n6968, MEM_stage_inst_dmem_n6967, MEM_stage_inst_dmem_n6966, MEM_stage_inst_dmem_n6965, MEM_stage_inst_dmem_n6964, MEM_stage_inst_dmem_n6963, MEM_stage_inst_dmem_n6962, MEM_stage_inst_dmem_n6961, MEM_stage_inst_dmem_n6960, MEM_stage_inst_dmem_n6959, MEM_stage_inst_dmem_n6958, MEM_stage_inst_dmem_n6957, MEM_stage_inst_dmem_n6956, MEM_stage_inst_dmem_n6955, MEM_stage_inst_dmem_n6954, MEM_stage_inst_dmem_n6953, MEM_stage_inst_dmem_n6952, MEM_stage_inst_dmem_n6951, MEM_stage_inst_dmem_n6950, MEM_stage_inst_dmem_n6949, MEM_stage_inst_dmem_n6948, MEM_stage_inst_dmem_n6947, MEM_stage_inst_dmem_n6946, MEM_stage_inst_dmem_n6945, MEM_stage_inst_dmem_n6944, MEM_stage_inst_dmem_n6943, MEM_stage_inst_dmem_n6942, MEM_stage_inst_dmem_n6941, MEM_stage_inst_dmem_n6940, MEM_stage_inst_dmem_n6939, MEM_stage_inst_dmem_n6938, MEM_stage_inst_dmem_n6937, MEM_stage_inst_dmem_n6936, MEM_stage_inst_dmem_n6935, MEM_stage_inst_dmem_n6934, MEM_stage_inst_dmem_n6933, MEM_stage_inst_dmem_n6932, MEM_stage_inst_dmem_n6931, MEM_stage_inst_dmem_n6930, MEM_stage_inst_dmem_n6929, MEM_stage_inst_dmem_n6928, MEM_stage_inst_dmem_n6927, MEM_stage_inst_dmem_n6926, MEM_stage_inst_dmem_n6925, MEM_stage_inst_dmem_n6924, MEM_stage_inst_dmem_n6923, MEM_stage_inst_dmem_n6922, MEM_stage_inst_dmem_n6921, MEM_stage_inst_dmem_n6920, MEM_stage_inst_dmem_n6919, MEM_stage_inst_dmem_n6918, MEM_stage_inst_dmem_n6917, MEM_stage_inst_dmem_n6916, MEM_stage_inst_dmem_n6915, MEM_stage_inst_dmem_n6914, MEM_stage_inst_dmem_n6913, MEM_stage_inst_dmem_n6912, MEM_stage_inst_dmem_n6911, MEM_stage_inst_dmem_n6910, MEM_stage_inst_dmem_n6909, MEM_stage_inst_dmem_n6908, MEM_stage_inst_dmem_n6907, MEM_stage_inst_dmem_n6906, MEM_stage_inst_dmem_n6905, MEM_stage_inst_dmem_n6904, MEM_stage_inst_dmem_n6903, MEM_stage_inst_dmem_n6902, MEM_stage_inst_dmem_n6901, MEM_stage_inst_dmem_n6900, MEM_stage_inst_dmem_n6899, MEM_stage_inst_dmem_n6898, MEM_stage_inst_dmem_n6897, MEM_stage_inst_dmem_n6896, MEM_stage_inst_dmem_n6895, MEM_stage_inst_dmem_n6894, MEM_stage_inst_dmem_n6893, MEM_stage_inst_dmem_n6892, MEM_stage_inst_dmem_n6891, MEM_stage_inst_dmem_n6890, MEM_stage_inst_dmem_n6889, MEM_stage_inst_dmem_n6888, MEM_stage_inst_dmem_n6887, MEM_stage_inst_dmem_n6886, MEM_stage_inst_dmem_n6885, MEM_stage_inst_dmem_n6884, MEM_stage_inst_dmem_n6883, MEM_stage_inst_dmem_n6882, MEM_stage_inst_dmem_n6881, MEM_stage_inst_dmem_n6880, MEM_stage_inst_dmem_n6879, MEM_stage_inst_dmem_n6878, MEM_stage_inst_dmem_n6877, MEM_stage_inst_dmem_n6876, MEM_stage_inst_dmem_n6875, MEM_stage_inst_dmem_n6874, MEM_stage_inst_dmem_n6873, MEM_stage_inst_dmem_n6872, MEM_stage_inst_dmem_n6871, MEM_stage_inst_dmem_n6870, MEM_stage_inst_dmem_n6869, MEM_stage_inst_dmem_n6868, MEM_stage_inst_dmem_n6867, MEM_stage_inst_dmem_n6866, MEM_stage_inst_dmem_n6865, MEM_stage_inst_dmem_n6864, MEM_stage_inst_dmem_n6863, MEM_stage_inst_dmem_n6862, MEM_stage_inst_dmem_n6861, MEM_stage_inst_dmem_n6860, MEM_stage_inst_dmem_n6859, MEM_stage_inst_dmem_n6858, MEM_stage_inst_dmem_n6857, MEM_stage_inst_dmem_n6856, MEM_stage_inst_dmem_n6855, MEM_stage_inst_dmem_n6854, MEM_stage_inst_dmem_n6853, MEM_stage_inst_dmem_n6852, MEM_stage_inst_dmem_n6851, MEM_stage_inst_dmem_n6850, MEM_stage_inst_dmem_n6849, MEM_stage_inst_dmem_n6848, MEM_stage_inst_dmem_n6847, MEM_stage_inst_dmem_n6846, MEM_stage_inst_dmem_n6845, MEM_stage_inst_dmem_n6844, MEM_stage_inst_dmem_n6843, MEM_stage_inst_dmem_n6842, MEM_stage_inst_dmem_n6841, MEM_stage_inst_dmem_n6840, MEM_stage_inst_dmem_n6839, MEM_stage_inst_dmem_n6838, MEM_stage_inst_dmem_n6837, MEM_stage_inst_dmem_n6836, MEM_stage_inst_dmem_n6835, MEM_stage_inst_dmem_n6834, MEM_stage_inst_dmem_n6833, MEM_stage_inst_dmem_n6832, MEM_stage_inst_dmem_n6831, MEM_stage_inst_dmem_n6830, MEM_stage_inst_dmem_n6829, MEM_stage_inst_dmem_n6828, MEM_stage_inst_dmem_n6827, MEM_stage_inst_dmem_n6826, MEM_stage_inst_dmem_n6825, MEM_stage_inst_dmem_n6824, MEM_stage_inst_dmem_n6823, MEM_stage_inst_dmem_n6822, MEM_stage_inst_dmem_n6821, MEM_stage_inst_dmem_n6820, MEM_stage_inst_dmem_n6819, MEM_stage_inst_dmem_n6818, MEM_stage_inst_dmem_n6817, MEM_stage_inst_dmem_n6816, MEM_stage_inst_dmem_n6815, MEM_stage_inst_dmem_n6814, MEM_stage_inst_dmem_n6813, MEM_stage_inst_dmem_n6812, MEM_stage_inst_dmem_n6811, MEM_stage_inst_dmem_n6810, MEM_stage_inst_dmem_n6809, MEM_stage_inst_dmem_n6808, MEM_stage_inst_dmem_n6807, MEM_stage_inst_dmem_n6806, MEM_stage_inst_dmem_n6805, MEM_stage_inst_dmem_n6804, MEM_stage_inst_dmem_n6803, MEM_stage_inst_dmem_n6802, MEM_stage_inst_dmem_n6801, MEM_stage_inst_dmem_n6800, MEM_stage_inst_dmem_n6799, MEM_stage_inst_dmem_n6798, MEM_stage_inst_dmem_n6797, MEM_stage_inst_dmem_n6796, MEM_stage_inst_dmem_n6795, MEM_stage_inst_dmem_n6794, MEM_stage_inst_dmem_n6793, MEM_stage_inst_dmem_n6792, MEM_stage_inst_dmem_n6791, MEM_stage_inst_dmem_n6790, MEM_stage_inst_dmem_n6789, MEM_stage_inst_dmem_n6788, MEM_stage_inst_dmem_n6787, MEM_stage_inst_dmem_n6786, MEM_stage_inst_dmem_n6785, MEM_stage_inst_dmem_n6784, MEM_stage_inst_dmem_n6783, MEM_stage_inst_dmem_n6782, MEM_stage_inst_dmem_n6781, MEM_stage_inst_dmem_n6780, MEM_stage_inst_dmem_n6779, MEM_stage_inst_dmem_n6778, MEM_stage_inst_dmem_n6777, MEM_stage_inst_dmem_n6776, MEM_stage_inst_dmem_n6775, MEM_stage_inst_dmem_n6774, MEM_stage_inst_dmem_n6773, MEM_stage_inst_dmem_n6772, MEM_stage_inst_dmem_n6771, MEM_stage_inst_dmem_n6770, MEM_stage_inst_dmem_n6769, MEM_stage_inst_dmem_n6768, MEM_stage_inst_dmem_n6767, MEM_stage_inst_dmem_n6766, MEM_stage_inst_dmem_n6765, MEM_stage_inst_dmem_n6764, MEM_stage_inst_dmem_n6763, MEM_stage_inst_dmem_n6762, MEM_stage_inst_dmem_n6761, MEM_stage_inst_dmem_n6760, MEM_stage_inst_dmem_n6759, MEM_stage_inst_dmem_n6758, MEM_stage_inst_dmem_n6757, MEM_stage_inst_dmem_n6756, MEM_stage_inst_dmem_n6755, MEM_stage_inst_dmem_n6754, MEM_stage_inst_dmem_n6753, MEM_stage_inst_dmem_n6752, MEM_stage_inst_dmem_n6751, MEM_stage_inst_dmem_n6750, MEM_stage_inst_dmem_n6749, MEM_stage_inst_dmem_n6748, MEM_stage_inst_dmem_n6747, MEM_stage_inst_dmem_n6746, MEM_stage_inst_dmem_n6745, MEM_stage_inst_dmem_n6744, MEM_stage_inst_dmem_n6743, MEM_stage_inst_dmem_n6742, MEM_stage_inst_dmem_n6741, MEM_stage_inst_dmem_n6740, MEM_stage_inst_dmem_n6739, MEM_stage_inst_dmem_n6738, MEM_stage_inst_dmem_n6737, MEM_stage_inst_dmem_n6736, MEM_stage_inst_dmem_n6735, MEM_stage_inst_dmem_n6734, MEM_stage_inst_dmem_n6733, MEM_stage_inst_dmem_n6732, MEM_stage_inst_dmem_n6731, MEM_stage_inst_dmem_n6730, MEM_stage_inst_dmem_n6729, MEM_stage_inst_dmem_n6728, MEM_stage_inst_dmem_n6727, MEM_stage_inst_dmem_n6726, MEM_stage_inst_dmem_n6725, MEM_stage_inst_dmem_n6724, MEM_stage_inst_dmem_n6723, MEM_stage_inst_dmem_n6722, MEM_stage_inst_dmem_n6721, MEM_stage_inst_dmem_n6720, MEM_stage_inst_dmem_n6719, MEM_stage_inst_dmem_n6718, MEM_stage_inst_dmem_n6717, MEM_stage_inst_dmem_n6716, MEM_stage_inst_dmem_n6715, MEM_stage_inst_dmem_n6714, MEM_stage_inst_dmem_n6713, MEM_stage_inst_dmem_n6712, MEM_stage_inst_dmem_n6711, MEM_stage_inst_dmem_n6710, MEM_stage_inst_dmem_n6709, MEM_stage_inst_dmem_n6708, MEM_stage_inst_dmem_n6707, MEM_stage_inst_dmem_n6706, MEM_stage_inst_dmem_n6705, MEM_stage_inst_dmem_n6704, MEM_stage_inst_dmem_n6703, MEM_stage_inst_dmem_n6702, MEM_stage_inst_dmem_n6701, MEM_stage_inst_dmem_n6700, MEM_stage_inst_dmem_n6699, MEM_stage_inst_dmem_n6698, MEM_stage_inst_dmem_n6697, MEM_stage_inst_dmem_n6696, MEM_stage_inst_dmem_n6695, MEM_stage_inst_dmem_n6694, MEM_stage_inst_dmem_n6693, MEM_stage_inst_dmem_n6692, MEM_stage_inst_dmem_n6691, MEM_stage_inst_dmem_n6690, MEM_stage_inst_dmem_n6689, MEM_stage_inst_dmem_n6688, MEM_stage_inst_dmem_n6687, MEM_stage_inst_dmem_n6686, MEM_stage_inst_dmem_n6685, MEM_stage_inst_dmem_n6684, MEM_stage_inst_dmem_n6683, MEM_stage_inst_dmem_n6682, MEM_stage_inst_dmem_n6681, MEM_stage_inst_dmem_n6680, MEM_stage_inst_dmem_n6679, MEM_stage_inst_dmem_n6678, MEM_stage_inst_dmem_n6677, MEM_stage_inst_dmem_n6676, MEM_stage_inst_dmem_n6675, MEM_stage_inst_dmem_n6674, MEM_stage_inst_dmem_n6673, MEM_stage_inst_dmem_n6672, MEM_stage_inst_dmem_n6671, MEM_stage_inst_dmem_n6670, MEM_stage_inst_dmem_n6669, MEM_stage_inst_dmem_n6668, MEM_stage_inst_dmem_n6667, MEM_stage_inst_dmem_n6666, MEM_stage_inst_dmem_n6665, MEM_stage_inst_dmem_n6664, MEM_stage_inst_dmem_n6663, MEM_stage_inst_dmem_n6662, MEM_stage_inst_dmem_n6661, MEM_stage_inst_dmem_n6660, MEM_stage_inst_dmem_n6659, MEM_stage_inst_dmem_n6658, MEM_stage_inst_dmem_n6657, MEM_stage_inst_dmem_n6656, MEM_stage_inst_dmem_n6655, MEM_stage_inst_dmem_n6654, MEM_stage_inst_dmem_n6653, MEM_stage_inst_dmem_n6652, MEM_stage_inst_dmem_n6651, MEM_stage_inst_dmem_n6650, MEM_stage_inst_dmem_n6649, MEM_stage_inst_dmem_n6648, MEM_stage_inst_dmem_n6647, MEM_stage_inst_dmem_n6646, MEM_stage_inst_dmem_n6645, MEM_stage_inst_dmem_n6644, MEM_stage_inst_dmem_n6643, MEM_stage_inst_dmem_n6642, MEM_stage_inst_dmem_n6641, MEM_stage_inst_dmem_n6640, MEM_stage_inst_dmem_n6639, MEM_stage_inst_dmem_n6638, MEM_stage_inst_dmem_n6637, MEM_stage_inst_dmem_n6636, MEM_stage_inst_dmem_n6635, MEM_stage_inst_dmem_n6634, MEM_stage_inst_dmem_n6633, MEM_stage_inst_dmem_n6632, MEM_stage_inst_dmem_n6631, MEM_stage_inst_dmem_n6630, MEM_stage_inst_dmem_n6629, MEM_stage_inst_dmem_n6628, MEM_stage_inst_dmem_n6627, MEM_stage_inst_dmem_n6626, MEM_stage_inst_dmem_n6625, MEM_stage_inst_dmem_n6624, MEM_stage_inst_dmem_n6623, MEM_stage_inst_dmem_n6622, MEM_stage_inst_dmem_n6621, MEM_stage_inst_dmem_n6620, MEM_stage_inst_dmem_n6619, MEM_stage_inst_dmem_n6618, MEM_stage_inst_dmem_n6617, MEM_stage_inst_dmem_n6616, MEM_stage_inst_dmem_n6615, MEM_stage_inst_dmem_n6614, MEM_stage_inst_dmem_n6613, MEM_stage_inst_dmem_n6612, MEM_stage_inst_dmem_n6611, MEM_stage_inst_dmem_n6610, MEM_stage_inst_dmem_n6609, MEM_stage_inst_dmem_n6608, MEM_stage_inst_dmem_n6607, MEM_stage_inst_dmem_n6606, MEM_stage_inst_dmem_n6605, MEM_stage_inst_dmem_n6604, MEM_stage_inst_dmem_n6603, MEM_stage_inst_dmem_n6602, MEM_stage_inst_dmem_n6601, MEM_stage_inst_dmem_n6600, MEM_stage_inst_dmem_n6599, MEM_stage_inst_dmem_n6598, MEM_stage_inst_dmem_n6597, MEM_stage_inst_dmem_n6596, MEM_stage_inst_dmem_n6595, MEM_stage_inst_dmem_n6594, MEM_stage_inst_dmem_n6593, MEM_stage_inst_dmem_n6592, MEM_stage_inst_dmem_n6591, MEM_stage_inst_dmem_n6590, MEM_stage_inst_dmem_n6589, MEM_stage_inst_dmem_n6588, MEM_stage_inst_dmem_n6587, MEM_stage_inst_dmem_n6586, MEM_stage_inst_dmem_n6585, MEM_stage_inst_dmem_n6584, MEM_stage_inst_dmem_n6583, MEM_stage_inst_dmem_n6582, MEM_stage_inst_dmem_n6581, MEM_stage_inst_dmem_n6580, MEM_stage_inst_dmem_n6579, MEM_stage_inst_dmem_n6578, MEM_stage_inst_dmem_n6577, MEM_stage_inst_dmem_n6576, MEM_stage_inst_dmem_n6575, MEM_stage_inst_dmem_n6574, MEM_stage_inst_dmem_n6573, MEM_stage_inst_dmem_n6572, MEM_stage_inst_dmem_n6571, MEM_stage_inst_dmem_n6570, MEM_stage_inst_dmem_n6569, MEM_stage_inst_dmem_n6568, MEM_stage_inst_dmem_n6567, MEM_stage_inst_dmem_n6566, MEM_stage_inst_dmem_n6565, MEM_stage_inst_dmem_n6564, MEM_stage_inst_dmem_n6563, MEM_stage_inst_dmem_n6562, MEM_stage_inst_dmem_n6561, MEM_stage_inst_dmem_n6560, MEM_stage_inst_dmem_n6559, MEM_stage_inst_dmem_n6558, MEM_stage_inst_dmem_n6557, MEM_stage_inst_dmem_n6556, MEM_stage_inst_dmem_n6555, MEM_stage_inst_dmem_n6554, MEM_stage_inst_dmem_n6553, MEM_stage_inst_dmem_n6552, MEM_stage_inst_dmem_n6551, MEM_stage_inst_dmem_n6550, MEM_stage_inst_dmem_n6549, MEM_stage_inst_dmem_n6548, MEM_stage_inst_dmem_n6547, MEM_stage_inst_dmem_n6546, MEM_stage_inst_dmem_n6545, MEM_stage_inst_dmem_n6544, MEM_stage_inst_dmem_n6543, MEM_stage_inst_dmem_n6542, MEM_stage_inst_dmem_n6541, MEM_stage_inst_dmem_n6540, MEM_stage_inst_dmem_n6539, MEM_stage_inst_dmem_n6538, MEM_stage_inst_dmem_n6537, MEM_stage_inst_dmem_n6536, MEM_stage_inst_dmem_n6535, MEM_stage_inst_dmem_n6534, MEM_stage_inst_dmem_n6533, MEM_stage_inst_dmem_n6532, MEM_stage_inst_dmem_n6531, MEM_stage_inst_dmem_n6530, MEM_stage_inst_dmem_n6529, MEM_stage_inst_dmem_n6528, MEM_stage_inst_dmem_n6527, MEM_stage_inst_dmem_n6526, MEM_stage_inst_dmem_n6525, MEM_stage_inst_dmem_n6524, MEM_stage_inst_dmem_n6523, MEM_stage_inst_dmem_n6522, MEM_stage_inst_dmem_n6521, MEM_stage_inst_dmem_n6520, MEM_stage_inst_dmem_n6519, MEM_stage_inst_dmem_n6518, MEM_stage_inst_dmem_n6517, MEM_stage_inst_dmem_n6516, MEM_stage_inst_dmem_n6515, MEM_stage_inst_dmem_n6514, MEM_stage_inst_dmem_n6513, MEM_stage_inst_dmem_n6512, MEM_stage_inst_dmem_n6511, MEM_stage_inst_dmem_n6510, MEM_stage_inst_dmem_n6509, MEM_stage_inst_dmem_n6508, MEM_stage_inst_dmem_n6507, MEM_stage_inst_dmem_n6506, MEM_stage_inst_dmem_n6505, MEM_stage_inst_dmem_n6504, MEM_stage_inst_dmem_n6503, MEM_stage_inst_dmem_n6502, MEM_stage_inst_dmem_n6501, MEM_stage_inst_dmem_n6500, MEM_stage_inst_dmem_n6499, MEM_stage_inst_dmem_n6498, MEM_stage_inst_dmem_n6497, MEM_stage_inst_dmem_n6496, MEM_stage_inst_dmem_n6495, MEM_stage_inst_dmem_n6494, MEM_stage_inst_dmem_n6493, MEM_stage_inst_dmem_n6492, MEM_stage_inst_dmem_n6491, MEM_stage_inst_dmem_n6490, MEM_stage_inst_dmem_n6489, MEM_stage_inst_dmem_n6488, MEM_stage_inst_dmem_n6487, MEM_stage_inst_dmem_n6486, MEM_stage_inst_dmem_n6485, MEM_stage_inst_dmem_n6484, MEM_stage_inst_dmem_n6483, MEM_stage_inst_dmem_n6482, MEM_stage_inst_dmem_n6481, MEM_stage_inst_dmem_n6480, MEM_stage_inst_dmem_n6479, MEM_stage_inst_dmem_n6478, MEM_stage_inst_dmem_n6477, MEM_stage_inst_dmem_n6476, MEM_stage_inst_dmem_n6475, MEM_stage_inst_dmem_n6474, MEM_stage_inst_dmem_n6473, MEM_stage_inst_dmem_n6472, MEM_stage_inst_dmem_n6471, MEM_stage_inst_dmem_n6470, MEM_stage_inst_dmem_n6469, MEM_stage_inst_dmem_n6468, MEM_stage_inst_dmem_n6467, MEM_stage_inst_dmem_n6466, MEM_stage_inst_dmem_n6465, MEM_stage_inst_dmem_n6464, MEM_stage_inst_dmem_n6463, MEM_stage_inst_dmem_n6462, MEM_stage_inst_dmem_n6461, MEM_stage_inst_dmem_n6460, MEM_stage_inst_dmem_n6459, MEM_stage_inst_dmem_n6458, MEM_stage_inst_dmem_n6457, MEM_stage_inst_dmem_n6456, MEM_stage_inst_dmem_n6455, MEM_stage_inst_dmem_n6454, MEM_stage_inst_dmem_n6453, MEM_stage_inst_dmem_n6452, MEM_stage_inst_dmem_n6451, MEM_stage_inst_dmem_n6450, MEM_stage_inst_dmem_n6449, MEM_stage_inst_dmem_n6448, MEM_stage_inst_dmem_n6447, MEM_stage_inst_dmem_n6446, MEM_stage_inst_dmem_n6445, MEM_stage_inst_dmem_n6444, MEM_stage_inst_dmem_n6443, MEM_stage_inst_dmem_n6442, MEM_stage_inst_dmem_n6441, MEM_stage_inst_dmem_n6440, MEM_stage_inst_dmem_n6439, MEM_stage_inst_dmem_n6438, MEM_stage_inst_dmem_n6437, MEM_stage_inst_dmem_n6436, MEM_stage_inst_dmem_n6435, MEM_stage_inst_dmem_n6434, MEM_stage_inst_dmem_n6433, MEM_stage_inst_dmem_n6432, MEM_stage_inst_dmem_n6431, MEM_stage_inst_dmem_n6430, MEM_stage_inst_dmem_n6429, MEM_stage_inst_dmem_n6428, MEM_stage_inst_dmem_n6427, MEM_stage_inst_dmem_n6426, MEM_stage_inst_dmem_n6425, MEM_stage_inst_dmem_n6424, MEM_stage_inst_dmem_n6423, MEM_stage_inst_dmem_n6422, MEM_stage_inst_dmem_n6421, MEM_stage_inst_dmem_n6420, MEM_stage_inst_dmem_n6419, MEM_stage_inst_dmem_n6418, MEM_stage_inst_dmem_n6417, MEM_stage_inst_dmem_n6416, MEM_stage_inst_dmem_n6415, MEM_stage_inst_dmem_n6414, MEM_stage_inst_dmem_n6413, MEM_stage_inst_dmem_n6412, MEM_stage_inst_dmem_n6411, MEM_stage_inst_dmem_n6410, MEM_stage_inst_dmem_n6409, MEM_stage_inst_dmem_n6408, MEM_stage_inst_dmem_n6407, MEM_stage_inst_dmem_n6406, MEM_stage_inst_dmem_n6405, MEM_stage_inst_dmem_n6404, MEM_stage_inst_dmem_n6403, MEM_stage_inst_dmem_n6402, MEM_stage_inst_dmem_n6401, MEM_stage_inst_dmem_n6400, MEM_stage_inst_dmem_n6399, MEM_stage_inst_dmem_n6398, MEM_stage_inst_dmem_n6397, MEM_stage_inst_dmem_n6396, MEM_stage_inst_dmem_n6395, MEM_stage_inst_dmem_n6394, MEM_stage_inst_dmem_n6393, MEM_stage_inst_dmem_n6392, MEM_stage_inst_dmem_n6391, MEM_stage_inst_dmem_n6390, MEM_stage_inst_dmem_n6389, MEM_stage_inst_dmem_n6388, MEM_stage_inst_dmem_n6387, MEM_stage_inst_dmem_n6386, MEM_stage_inst_dmem_n6385, MEM_stage_inst_dmem_n6384, MEM_stage_inst_dmem_n6383, MEM_stage_inst_dmem_n6382, MEM_stage_inst_dmem_n6381, MEM_stage_inst_dmem_n6380, MEM_stage_inst_dmem_n6379, MEM_stage_inst_dmem_n6378, MEM_stage_inst_dmem_n6377, MEM_stage_inst_dmem_n6376, MEM_stage_inst_dmem_n6375, MEM_stage_inst_dmem_n6374, MEM_stage_inst_dmem_n6373, MEM_stage_inst_dmem_n6372, MEM_stage_inst_dmem_n6371, MEM_stage_inst_dmem_n6370, MEM_stage_inst_dmem_n6369, MEM_stage_inst_dmem_n6368, MEM_stage_inst_dmem_n6367, MEM_stage_inst_dmem_n6366, MEM_stage_inst_dmem_n6365, MEM_stage_inst_dmem_n6364, MEM_stage_inst_dmem_n6363, MEM_stage_inst_dmem_n6362, MEM_stage_inst_dmem_n6361, MEM_stage_inst_dmem_n6360, MEM_stage_inst_dmem_n6359, MEM_stage_inst_dmem_n6358, MEM_stage_inst_dmem_n6357, MEM_stage_inst_dmem_n6356, MEM_stage_inst_dmem_n6355, MEM_stage_inst_dmem_n6354, MEM_stage_inst_dmem_n6353, MEM_stage_inst_dmem_n6352, MEM_stage_inst_dmem_n6351, MEM_stage_inst_dmem_n6350, MEM_stage_inst_dmem_n6349, MEM_stage_inst_dmem_n6348, MEM_stage_inst_dmem_n6347, MEM_stage_inst_dmem_n6346, MEM_stage_inst_dmem_n6345, MEM_stage_inst_dmem_n6344, MEM_stage_inst_dmem_n6343, MEM_stage_inst_dmem_n6342, MEM_stage_inst_dmem_n6341, MEM_stage_inst_dmem_n6340, MEM_stage_inst_dmem_n6339, MEM_stage_inst_dmem_n6338, MEM_stage_inst_dmem_n6337, MEM_stage_inst_dmem_n6336, MEM_stage_inst_dmem_n6335, MEM_stage_inst_dmem_n6334, MEM_stage_inst_dmem_n6333, MEM_stage_inst_dmem_n6332, MEM_stage_inst_dmem_n6331, MEM_stage_inst_dmem_n6330, MEM_stage_inst_dmem_n6329, MEM_stage_inst_dmem_n6328, MEM_stage_inst_dmem_n6327, MEM_stage_inst_dmem_n6326, MEM_stage_inst_dmem_n6325, MEM_stage_inst_dmem_n6324, MEM_stage_inst_dmem_n6323, MEM_stage_inst_dmem_n6322, MEM_stage_inst_dmem_n6321, MEM_stage_inst_dmem_n6320, MEM_stage_inst_dmem_n6319, MEM_stage_inst_dmem_n6318, MEM_stage_inst_dmem_n6317, MEM_stage_inst_dmem_n6316, MEM_stage_inst_dmem_n6315, MEM_stage_inst_dmem_n6314, MEM_stage_inst_dmem_n6313, MEM_stage_inst_dmem_n6312, MEM_stage_inst_dmem_n6311, MEM_stage_inst_dmem_n6310, MEM_stage_inst_dmem_n6309, MEM_stage_inst_dmem_n6308, MEM_stage_inst_dmem_n6307, MEM_stage_inst_dmem_n6306, MEM_stage_inst_dmem_n6305, MEM_stage_inst_dmem_n6304, MEM_stage_inst_dmem_n6303, MEM_stage_inst_dmem_n6302, MEM_stage_inst_dmem_n6301, MEM_stage_inst_dmem_n6300, MEM_stage_inst_dmem_n6299, MEM_stage_inst_dmem_n6298, MEM_stage_inst_dmem_n6297, MEM_stage_inst_dmem_n6296, MEM_stage_inst_dmem_n6295, MEM_stage_inst_dmem_n6294, MEM_stage_inst_dmem_n6293, MEM_stage_inst_dmem_n6292, MEM_stage_inst_dmem_n6291, MEM_stage_inst_dmem_n6290, MEM_stage_inst_dmem_n6289, MEM_stage_inst_dmem_n6288, MEM_stage_inst_dmem_n6287, MEM_stage_inst_dmem_n6286, MEM_stage_inst_dmem_n6285, MEM_stage_inst_dmem_n6284, MEM_stage_inst_dmem_n6283, MEM_stage_inst_dmem_n6282, MEM_stage_inst_dmem_n6281, MEM_stage_inst_dmem_n6280, MEM_stage_inst_dmem_n6279, MEM_stage_inst_dmem_n6278, MEM_stage_inst_dmem_n6277, MEM_stage_inst_dmem_n6276, MEM_stage_inst_dmem_n6275, MEM_stage_inst_dmem_n6274, MEM_stage_inst_dmem_n6273, MEM_stage_inst_dmem_n6272, MEM_stage_inst_dmem_n6271, MEM_stage_inst_dmem_n6270, MEM_stage_inst_dmem_n6269, MEM_stage_inst_dmem_n6268, MEM_stage_inst_dmem_n6267, MEM_stage_inst_dmem_n6266, MEM_stage_inst_dmem_n6265, MEM_stage_inst_dmem_n6264, MEM_stage_inst_dmem_n6263, MEM_stage_inst_dmem_n6262, MEM_stage_inst_dmem_n6261, MEM_stage_inst_dmem_n6260, MEM_stage_inst_dmem_n6259, MEM_stage_inst_dmem_n6258, MEM_stage_inst_dmem_n6257, MEM_stage_inst_dmem_n6256, MEM_stage_inst_dmem_n6255, MEM_stage_inst_dmem_n6254, MEM_stage_inst_dmem_n6253, MEM_stage_inst_dmem_n6252, MEM_stage_inst_dmem_n6251, MEM_stage_inst_dmem_n6250, MEM_stage_inst_dmem_n6249, MEM_stage_inst_dmem_n6248, MEM_stage_inst_dmem_n6247, MEM_stage_inst_dmem_n6246, MEM_stage_inst_dmem_n6245, MEM_stage_inst_dmem_n6244, MEM_stage_inst_dmem_n6243, MEM_stage_inst_dmem_n6242, MEM_stage_inst_dmem_n6241, MEM_stage_inst_dmem_n6240, MEM_stage_inst_dmem_n6239, MEM_stage_inst_dmem_n6238, MEM_stage_inst_dmem_n6237, MEM_stage_inst_dmem_n6236, MEM_stage_inst_dmem_n6235, MEM_stage_inst_dmem_n6234, MEM_stage_inst_dmem_n6233, MEM_stage_inst_dmem_n6232, MEM_stage_inst_dmem_n6231, MEM_stage_inst_dmem_n6230, MEM_stage_inst_dmem_n6229, MEM_stage_inst_dmem_n6228, MEM_stage_inst_dmem_n6227, MEM_stage_inst_dmem_n6226, MEM_stage_inst_dmem_n6225, MEM_stage_inst_dmem_n6224, MEM_stage_inst_dmem_n6223, MEM_stage_inst_dmem_n6222, MEM_stage_inst_dmem_n6221, MEM_stage_inst_dmem_n6220, MEM_stage_inst_dmem_n6219, MEM_stage_inst_dmem_n6218, MEM_stage_inst_dmem_n6217, MEM_stage_inst_dmem_n6216, MEM_stage_inst_dmem_n6215, MEM_stage_inst_dmem_n6214, MEM_stage_inst_dmem_n6213, MEM_stage_inst_dmem_n6212, MEM_stage_inst_dmem_n6211, MEM_stage_inst_dmem_n6210, MEM_stage_inst_dmem_n6209, MEM_stage_inst_dmem_n6208, MEM_stage_inst_dmem_n6207, MEM_stage_inst_dmem_n6206, MEM_stage_inst_dmem_n6205, MEM_stage_inst_dmem_n6204, MEM_stage_inst_dmem_n6203, MEM_stage_inst_dmem_n6202, MEM_stage_inst_dmem_n6201, MEM_stage_inst_dmem_n6200, MEM_stage_inst_dmem_n6199, MEM_stage_inst_dmem_n6198, MEM_stage_inst_dmem_n6197, MEM_stage_inst_dmem_n6196, MEM_stage_inst_dmem_n6195, MEM_stage_inst_dmem_n6194, MEM_stage_inst_dmem_n6193, MEM_stage_inst_dmem_n6192, MEM_stage_inst_dmem_n6191, MEM_stage_inst_dmem_n6190, MEM_stage_inst_dmem_n6189, MEM_stage_inst_dmem_n6188, MEM_stage_inst_dmem_n6187, MEM_stage_inst_dmem_n6186, MEM_stage_inst_dmem_n6185, MEM_stage_inst_dmem_n6184, MEM_stage_inst_dmem_n6183, MEM_stage_inst_dmem_n6182, MEM_stage_inst_dmem_n6181, MEM_stage_inst_dmem_n6180, MEM_stage_inst_dmem_n6179, MEM_stage_inst_dmem_n6178, MEM_stage_inst_dmem_n6177, MEM_stage_inst_dmem_n6176, MEM_stage_inst_dmem_n6175, MEM_stage_inst_dmem_n6174, MEM_stage_inst_dmem_n6173, MEM_stage_inst_dmem_n6172, MEM_stage_inst_dmem_n6171, MEM_stage_inst_dmem_n6170, MEM_stage_inst_dmem_n6169, MEM_stage_inst_dmem_n6168, MEM_stage_inst_dmem_n6167, MEM_stage_inst_dmem_n6166, MEM_stage_inst_dmem_n6165, MEM_stage_inst_dmem_n6164, MEM_stage_inst_dmem_n6163, MEM_stage_inst_dmem_n6162, MEM_stage_inst_dmem_n6161, MEM_stage_inst_dmem_n6160, MEM_stage_inst_dmem_n6159, MEM_stage_inst_dmem_n6158, MEM_stage_inst_dmem_n6157, MEM_stage_inst_dmem_n6156, MEM_stage_inst_dmem_n6155, MEM_stage_inst_dmem_n6154, MEM_stage_inst_dmem_n6153, MEM_stage_inst_dmem_n6152, MEM_stage_inst_dmem_n6151, MEM_stage_inst_dmem_n6150, MEM_stage_inst_dmem_n6149, MEM_stage_inst_dmem_n6148, MEM_stage_inst_dmem_n6147, MEM_stage_inst_dmem_n6146, MEM_stage_inst_dmem_n6145, MEM_stage_inst_dmem_n6144, MEM_stage_inst_dmem_n6143, MEM_stage_inst_dmem_n6142, MEM_stage_inst_dmem_n6141, MEM_stage_inst_dmem_n6140, MEM_stage_inst_dmem_n6139, MEM_stage_inst_dmem_n6138, MEM_stage_inst_dmem_n6137, MEM_stage_inst_dmem_n6136, MEM_stage_inst_dmem_n6135, MEM_stage_inst_dmem_n6134, MEM_stage_inst_dmem_n6133, MEM_stage_inst_dmem_n6132, MEM_stage_inst_dmem_n6131, MEM_stage_inst_dmem_n6130, MEM_stage_inst_dmem_n6129, MEM_stage_inst_dmem_n6128, MEM_stage_inst_dmem_n6127, MEM_stage_inst_dmem_n6126, MEM_stage_inst_dmem_n6125, MEM_stage_inst_dmem_n6124, MEM_stage_inst_dmem_n6123, MEM_stage_inst_dmem_n6122, MEM_stage_inst_dmem_n6121, MEM_stage_inst_dmem_n6120, MEM_stage_inst_dmem_n6119, MEM_stage_inst_dmem_n6118, MEM_stage_inst_dmem_n6117, MEM_stage_inst_dmem_n6116, MEM_stage_inst_dmem_n6115, MEM_stage_inst_dmem_n6114, MEM_stage_inst_dmem_n6113, MEM_stage_inst_dmem_n6112, MEM_stage_inst_dmem_n6111, MEM_stage_inst_dmem_n6110, MEM_stage_inst_dmem_n6109, MEM_stage_inst_dmem_n6108, MEM_stage_inst_dmem_n6107, MEM_stage_inst_dmem_n6106, MEM_stage_inst_dmem_n6105, MEM_stage_inst_dmem_n6104, MEM_stage_inst_dmem_n6103, MEM_stage_inst_dmem_n6102, MEM_stage_inst_dmem_n6101, MEM_stage_inst_dmem_n6100, MEM_stage_inst_dmem_n6099, MEM_stage_inst_dmem_n6098, MEM_stage_inst_dmem_n6097, MEM_stage_inst_dmem_n6096, MEM_stage_inst_dmem_n6095, MEM_stage_inst_dmem_n6094, MEM_stage_inst_dmem_n6093, MEM_stage_inst_dmem_n6092, MEM_stage_inst_dmem_n6091, MEM_stage_inst_dmem_n6090, MEM_stage_inst_dmem_n6089, MEM_stage_inst_dmem_n6088, MEM_stage_inst_dmem_n6087, MEM_stage_inst_dmem_n6086, MEM_stage_inst_dmem_n6085, MEM_stage_inst_dmem_n6084, MEM_stage_inst_dmem_n6083, MEM_stage_inst_dmem_n6082, MEM_stage_inst_dmem_n6081, MEM_stage_inst_dmem_n6080, MEM_stage_inst_dmem_n6079, MEM_stage_inst_dmem_n6078, MEM_stage_inst_dmem_n6077, MEM_stage_inst_dmem_n6076, MEM_stage_inst_dmem_n6075, MEM_stage_inst_dmem_n6074, MEM_stage_inst_dmem_n6073, MEM_stage_inst_dmem_n6072, MEM_stage_inst_dmem_n6071, MEM_stage_inst_dmem_n6070, MEM_stage_inst_dmem_n6069, MEM_stage_inst_dmem_n6068, MEM_stage_inst_dmem_n6067, MEM_stage_inst_dmem_n6066, MEM_stage_inst_dmem_n6065, MEM_stage_inst_dmem_n6064, MEM_stage_inst_dmem_n6063, MEM_stage_inst_dmem_n6062, MEM_stage_inst_dmem_n6061, MEM_stage_inst_dmem_n6060, MEM_stage_inst_dmem_n6059, MEM_stage_inst_dmem_n6058, MEM_stage_inst_dmem_n6057, MEM_stage_inst_dmem_n6056, MEM_stage_inst_dmem_n6055, MEM_stage_inst_dmem_n6054, MEM_stage_inst_dmem_n6053, MEM_stage_inst_dmem_n6052, MEM_stage_inst_dmem_n6051, MEM_stage_inst_dmem_n6050, MEM_stage_inst_dmem_n6049, MEM_stage_inst_dmem_n6048, MEM_stage_inst_dmem_n6047, MEM_stage_inst_dmem_n6046, MEM_stage_inst_dmem_n6045, MEM_stage_inst_dmem_n6044, MEM_stage_inst_dmem_n6043, MEM_stage_inst_dmem_n6042, MEM_stage_inst_dmem_n6041, MEM_stage_inst_dmem_n6040, MEM_stage_inst_dmem_n6039, MEM_stage_inst_dmem_n6038, MEM_stage_inst_dmem_n6037, MEM_stage_inst_dmem_n6036, MEM_stage_inst_dmem_n6035, MEM_stage_inst_dmem_n6034, MEM_stage_inst_dmem_n6033, MEM_stage_inst_dmem_n6032, MEM_stage_inst_dmem_n6031, MEM_stage_inst_dmem_n6030, MEM_stage_inst_dmem_n6029, MEM_stage_inst_dmem_n6028, MEM_stage_inst_dmem_n6027, MEM_stage_inst_dmem_n6026, MEM_stage_inst_dmem_n6025, MEM_stage_inst_dmem_n6024, MEM_stage_inst_dmem_n6023, MEM_stage_inst_dmem_n6022, MEM_stage_inst_dmem_n6021, MEM_stage_inst_dmem_n6020, MEM_stage_inst_dmem_n6019, MEM_stage_inst_dmem_n6018, MEM_stage_inst_dmem_n6017, MEM_stage_inst_dmem_n6016, MEM_stage_inst_dmem_n6015, MEM_stage_inst_dmem_n6014, MEM_stage_inst_dmem_n6013, MEM_stage_inst_dmem_n6012, MEM_stage_inst_dmem_n6011, MEM_stage_inst_dmem_n6010, MEM_stage_inst_dmem_n6009, MEM_stage_inst_dmem_n6008, MEM_stage_inst_dmem_n6007, MEM_stage_inst_dmem_n6006, MEM_stage_inst_dmem_n6005, MEM_stage_inst_dmem_n6004, MEM_stage_inst_dmem_n6003, MEM_stage_inst_dmem_n6002, MEM_stage_inst_dmem_n6001, MEM_stage_inst_dmem_n6000, MEM_stage_inst_dmem_n5999, MEM_stage_inst_dmem_n5998, MEM_stage_inst_dmem_n5997, MEM_stage_inst_dmem_n5996, MEM_stage_inst_dmem_n5995, MEM_stage_inst_dmem_n5994, MEM_stage_inst_dmem_n5993, MEM_stage_inst_dmem_n5992, MEM_stage_inst_dmem_n5991, MEM_stage_inst_dmem_n5990, MEM_stage_inst_dmem_n5989, MEM_stage_inst_dmem_n5988, MEM_stage_inst_dmem_n5987, MEM_stage_inst_dmem_n5986, MEM_stage_inst_dmem_n5985, MEM_stage_inst_dmem_n5984, MEM_stage_inst_dmem_n5983, MEM_stage_inst_dmem_n5982, MEM_stage_inst_dmem_n5981, MEM_stage_inst_dmem_n5980, MEM_stage_inst_dmem_n5979, MEM_stage_inst_dmem_n5978, MEM_stage_inst_dmem_n5977, MEM_stage_inst_dmem_n5976, MEM_stage_inst_dmem_n5975, MEM_stage_inst_dmem_n5974, MEM_stage_inst_dmem_n5973, MEM_stage_inst_dmem_n5972, MEM_stage_inst_dmem_n5971, MEM_stage_inst_dmem_n5970, MEM_stage_inst_dmem_n5969, MEM_stage_inst_dmem_n5968, MEM_stage_inst_dmem_n5967, MEM_stage_inst_dmem_n5966, MEM_stage_inst_dmem_n5965, MEM_stage_inst_dmem_n5964, MEM_stage_inst_dmem_n5963, MEM_stage_inst_dmem_n5962, MEM_stage_inst_dmem_n5961, MEM_stage_inst_dmem_n5960, MEM_stage_inst_dmem_n5959, MEM_stage_inst_dmem_n5958, MEM_stage_inst_dmem_n5957, MEM_stage_inst_dmem_n5956, MEM_stage_inst_dmem_n5955, MEM_stage_inst_dmem_n5954, MEM_stage_inst_dmem_n5953, MEM_stage_inst_dmem_n5952, MEM_stage_inst_dmem_n5951, MEM_stage_inst_dmem_n5950, MEM_stage_inst_dmem_n5949, MEM_stage_inst_dmem_n5948, MEM_stage_inst_dmem_n5947, MEM_stage_inst_dmem_n5946, MEM_stage_inst_dmem_n5945, MEM_stage_inst_dmem_n5944, MEM_stage_inst_dmem_n5943, MEM_stage_inst_dmem_n5942, MEM_stage_inst_dmem_n5941, MEM_stage_inst_dmem_n5940, MEM_stage_inst_dmem_n5939, MEM_stage_inst_dmem_n5938, MEM_stage_inst_dmem_n5937, MEM_stage_inst_dmem_n5936, MEM_stage_inst_dmem_n5935, MEM_stage_inst_dmem_n5934, MEM_stage_inst_dmem_n5933, MEM_stage_inst_dmem_n5932, MEM_stage_inst_dmem_n5931, MEM_stage_inst_dmem_n5930, MEM_stage_inst_dmem_n5929, MEM_stage_inst_dmem_n5928, MEM_stage_inst_dmem_n5927, MEM_stage_inst_dmem_n5926, MEM_stage_inst_dmem_n5925, MEM_stage_inst_dmem_n5924, MEM_stage_inst_dmem_n5923, MEM_stage_inst_dmem_n5922, MEM_stage_inst_dmem_n5921, MEM_stage_inst_dmem_n5920, MEM_stage_inst_dmem_n5919, MEM_stage_inst_dmem_n5918, MEM_stage_inst_dmem_n5917, MEM_stage_inst_dmem_n5916, MEM_stage_inst_dmem_n5915, MEM_stage_inst_dmem_n5914, MEM_stage_inst_dmem_n5913, MEM_stage_inst_dmem_n5912, MEM_stage_inst_dmem_n5911, MEM_stage_inst_dmem_n5910, MEM_stage_inst_dmem_n5909, MEM_stage_inst_dmem_n5908, MEM_stage_inst_dmem_n5907, MEM_stage_inst_dmem_n5906, MEM_stage_inst_dmem_n5905, MEM_stage_inst_dmem_n5904, MEM_stage_inst_dmem_n5903, MEM_stage_inst_dmem_n5902, MEM_stage_inst_dmem_n5901, MEM_stage_inst_dmem_n5900, MEM_stage_inst_dmem_n5899, MEM_stage_inst_dmem_n5898, MEM_stage_inst_dmem_n5897, MEM_stage_inst_dmem_n5896, MEM_stage_inst_dmem_n5895, MEM_stage_inst_dmem_n5894, MEM_stage_inst_dmem_n5893, MEM_stage_inst_dmem_n5892, MEM_stage_inst_dmem_n5891, MEM_stage_inst_dmem_n5890, MEM_stage_inst_dmem_n5889, MEM_stage_inst_dmem_n5888, MEM_stage_inst_dmem_n5887, MEM_stage_inst_dmem_n5886, MEM_stage_inst_dmem_n5885, MEM_stage_inst_dmem_n5884, MEM_stage_inst_dmem_n5883, MEM_stage_inst_dmem_n5882, MEM_stage_inst_dmem_n5881, MEM_stage_inst_dmem_n5880, MEM_stage_inst_dmem_n5879, MEM_stage_inst_dmem_n5878, MEM_stage_inst_dmem_n5877, MEM_stage_inst_dmem_n5876, MEM_stage_inst_dmem_n5875, MEM_stage_inst_dmem_n5874, MEM_stage_inst_dmem_n5873, MEM_stage_inst_dmem_n5872, MEM_stage_inst_dmem_n5871, MEM_stage_inst_dmem_n5870, MEM_stage_inst_dmem_n5869, MEM_stage_inst_dmem_n5868, MEM_stage_inst_dmem_n5867, MEM_stage_inst_dmem_n5866, MEM_stage_inst_dmem_n5865, MEM_stage_inst_dmem_n5864, MEM_stage_inst_dmem_n5863, MEM_stage_inst_dmem_n5862, MEM_stage_inst_dmem_n5861, MEM_stage_inst_dmem_n5860, MEM_stage_inst_dmem_n5859, MEM_stage_inst_dmem_n5858, MEM_stage_inst_dmem_n5857, MEM_stage_inst_dmem_n5856, MEM_stage_inst_dmem_n5855, MEM_stage_inst_dmem_n5854, MEM_stage_inst_dmem_n5853, MEM_stage_inst_dmem_n5852, MEM_stage_inst_dmem_n5851, MEM_stage_inst_dmem_n5850, MEM_stage_inst_dmem_n5849, MEM_stage_inst_dmem_n5848, MEM_stage_inst_dmem_n5847, MEM_stage_inst_dmem_n5846, MEM_stage_inst_dmem_n5845, MEM_stage_inst_dmem_n5844, MEM_stage_inst_dmem_n5843, MEM_stage_inst_dmem_n5842, MEM_stage_inst_dmem_n5841, MEM_stage_inst_dmem_n5840, MEM_stage_inst_dmem_n5839, MEM_stage_inst_dmem_n5838, MEM_stage_inst_dmem_n5837, MEM_stage_inst_dmem_n5836, MEM_stage_inst_dmem_n5835, MEM_stage_inst_dmem_n5834, MEM_stage_inst_dmem_n5833, MEM_stage_inst_dmem_n5832, MEM_stage_inst_dmem_n5831, MEM_stage_inst_dmem_n5830, MEM_stage_inst_dmem_n5829, MEM_stage_inst_dmem_n5828, MEM_stage_inst_dmem_n5827, MEM_stage_inst_dmem_n5826, MEM_stage_inst_dmem_n5825, MEM_stage_inst_dmem_n5824, MEM_stage_inst_dmem_n5823, MEM_stage_inst_dmem_n5822, MEM_stage_inst_dmem_n5821, MEM_stage_inst_dmem_n5820, MEM_stage_inst_dmem_n5819, MEM_stage_inst_dmem_n5818, MEM_stage_inst_dmem_n5817, MEM_stage_inst_dmem_n5816, MEM_stage_inst_dmem_n5815, MEM_stage_inst_dmem_n5814, MEM_stage_inst_dmem_n5813, MEM_stage_inst_dmem_n5812, MEM_stage_inst_dmem_n5811, MEM_stage_inst_dmem_n5810, MEM_stage_inst_dmem_n5809, MEM_stage_inst_dmem_n5808, MEM_stage_inst_dmem_n5807, MEM_stage_inst_dmem_n5806, MEM_stage_inst_dmem_n5805, MEM_stage_inst_dmem_n5804, MEM_stage_inst_dmem_n5803, MEM_stage_inst_dmem_n5802, MEM_stage_inst_dmem_n5801, MEM_stage_inst_dmem_n5800, MEM_stage_inst_dmem_n5799, MEM_stage_inst_dmem_n5798, MEM_stage_inst_dmem_n5797, MEM_stage_inst_dmem_n5796, MEM_stage_inst_dmem_n5795, MEM_stage_inst_dmem_n5794, MEM_stage_inst_dmem_n5793, MEM_stage_inst_dmem_n5792, MEM_stage_inst_dmem_n5791, MEM_stage_inst_dmem_n5790, MEM_stage_inst_dmem_n5789, MEM_stage_inst_dmem_n5788, MEM_stage_inst_dmem_n5787, MEM_stage_inst_dmem_n5786, MEM_stage_inst_dmem_n5785, MEM_stage_inst_dmem_n5784, MEM_stage_inst_dmem_n5783, MEM_stage_inst_dmem_n5782, MEM_stage_inst_dmem_n5781, MEM_stage_inst_dmem_n5780, MEM_stage_inst_dmem_n5779, MEM_stage_inst_dmem_n5778, MEM_stage_inst_dmem_n5777, MEM_stage_inst_dmem_n5776, MEM_stage_inst_dmem_n5775, MEM_stage_inst_dmem_n5774, MEM_stage_inst_dmem_n5773, MEM_stage_inst_dmem_n5772, MEM_stage_inst_dmem_n5771, MEM_stage_inst_dmem_n5770, MEM_stage_inst_dmem_n5769, MEM_stage_inst_dmem_n5768, MEM_stage_inst_dmem_n5767, MEM_stage_inst_dmem_n5766, MEM_stage_inst_dmem_n5765, MEM_stage_inst_dmem_n5764, MEM_stage_inst_dmem_n5763, MEM_stage_inst_dmem_n5762, MEM_stage_inst_dmem_n5761, MEM_stage_inst_dmem_n5760, MEM_stage_inst_dmem_n5759, MEM_stage_inst_dmem_n5758, MEM_stage_inst_dmem_n5757, MEM_stage_inst_dmem_n5756, MEM_stage_inst_dmem_n5755, MEM_stage_inst_dmem_n5754, MEM_stage_inst_dmem_n5753, MEM_stage_inst_dmem_n5752, MEM_stage_inst_dmem_n5751, MEM_stage_inst_dmem_n5750, MEM_stage_inst_dmem_n5749, MEM_stage_inst_dmem_n5748, MEM_stage_inst_dmem_n5747, MEM_stage_inst_dmem_n5746, MEM_stage_inst_dmem_n5745, MEM_stage_inst_dmem_n5744, MEM_stage_inst_dmem_n5743, MEM_stage_inst_dmem_n5742, MEM_stage_inst_dmem_n5741, MEM_stage_inst_dmem_n5740, MEM_stage_inst_dmem_n5739, MEM_stage_inst_dmem_n5738, MEM_stage_inst_dmem_n5737, MEM_stage_inst_dmem_n5736, MEM_stage_inst_dmem_n5735, MEM_stage_inst_dmem_n5734, MEM_stage_inst_dmem_n5733, MEM_stage_inst_dmem_n5732, MEM_stage_inst_dmem_n5731, MEM_stage_inst_dmem_n5730, MEM_stage_inst_dmem_n5729, MEM_stage_inst_dmem_n5728, MEM_stage_inst_dmem_n5727, MEM_stage_inst_dmem_n5726, MEM_stage_inst_dmem_n5725, MEM_stage_inst_dmem_n5724, MEM_stage_inst_dmem_n5723, MEM_stage_inst_dmem_n5722, MEM_stage_inst_dmem_n5721, MEM_stage_inst_dmem_n5720, MEM_stage_inst_dmem_n5719, MEM_stage_inst_dmem_n5718, MEM_stage_inst_dmem_n5717, MEM_stage_inst_dmem_n5716, MEM_stage_inst_dmem_n5715, MEM_stage_inst_dmem_n5714, MEM_stage_inst_dmem_n5713, MEM_stage_inst_dmem_n5712, MEM_stage_inst_dmem_n5711, MEM_stage_inst_dmem_n5710, MEM_stage_inst_dmem_n5709, MEM_stage_inst_dmem_n5708, MEM_stage_inst_dmem_n5707, MEM_stage_inst_dmem_n5706, MEM_stage_inst_dmem_n5705, MEM_stage_inst_dmem_n5704, MEM_stage_inst_dmem_n5703, MEM_stage_inst_dmem_n5702, MEM_stage_inst_dmem_n5701, MEM_stage_inst_dmem_n5700, MEM_stage_inst_dmem_n5699, MEM_stage_inst_dmem_n5698, MEM_stage_inst_dmem_n5697, MEM_stage_inst_dmem_n5696, MEM_stage_inst_dmem_n5695, MEM_stage_inst_dmem_n5694, MEM_stage_inst_dmem_n5693, MEM_stage_inst_dmem_n5692, MEM_stage_inst_dmem_n5691, MEM_stage_inst_dmem_n5690, MEM_stage_inst_dmem_n5689, MEM_stage_inst_dmem_n5688, MEM_stage_inst_dmem_n5687, MEM_stage_inst_dmem_n5686, MEM_stage_inst_dmem_n5685, MEM_stage_inst_dmem_n5684, MEM_stage_inst_dmem_n5683, MEM_stage_inst_dmem_n5682, MEM_stage_inst_dmem_n5681, MEM_stage_inst_dmem_n5680, MEM_stage_inst_dmem_n5679, MEM_stage_inst_dmem_n5678, MEM_stage_inst_dmem_n5677, MEM_stage_inst_dmem_n5676, MEM_stage_inst_dmem_n5675, MEM_stage_inst_dmem_n5674, MEM_stage_inst_dmem_n5673, MEM_stage_inst_dmem_n5672, MEM_stage_inst_dmem_n5671, MEM_stage_inst_dmem_n5670, MEM_stage_inst_dmem_n5669, MEM_stage_inst_dmem_n5668, MEM_stage_inst_dmem_n5667, MEM_stage_inst_dmem_n5666, MEM_stage_inst_dmem_n5665, MEM_stage_inst_dmem_n5664, MEM_stage_inst_dmem_n5663, MEM_stage_inst_dmem_n5662, MEM_stage_inst_dmem_n5661, MEM_stage_inst_dmem_n5660, MEM_stage_inst_dmem_n5659, MEM_stage_inst_dmem_n5658, MEM_stage_inst_dmem_n5657, MEM_stage_inst_dmem_n5656, MEM_stage_inst_dmem_n5655, MEM_stage_inst_dmem_n5654, MEM_stage_inst_dmem_n5653, MEM_stage_inst_dmem_n5652, MEM_stage_inst_dmem_n5651, MEM_stage_inst_dmem_n5650, MEM_stage_inst_dmem_n5649, MEM_stage_inst_dmem_n5648, MEM_stage_inst_dmem_n5647, MEM_stage_inst_dmem_n5646, MEM_stage_inst_dmem_n5645, MEM_stage_inst_dmem_n5644, MEM_stage_inst_dmem_n5643, MEM_stage_inst_dmem_n5642, MEM_stage_inst_dmem_n5641, MEM_stage_inst_dmem_n5640, MEM_stage_inst_dmem_n5639, MEM_stage_inst_dmem_n5638, MEM_stage_inst_dmem_n5637, MEM_stage_inst_dmem_n5636, MEM_stage_inst_dmem_n5635, MEM_stage_inst_dmem_n5634, MEM_stage_inst_dmem_n5633, MEM_stage_inst_dmem_n5632, MEM_stage_inst_dmem_n5631, MEM_stage_inst_dmem_n5630, MEM_stage_inst_dmem_n5629, MEM_stage_inst_dmem_n5628, MEM_stage_inst_dmem_n5627, MEM_stage_inst_dmem_n5626, MEM_stage_inst_dmem_n5625, MEM_stage_inst_dmem_n5624, MEM_stage_inst_dmem_n5623, MEM_stage_inst_dmem_n5622, MEM_stage_inst_dmem_n5621, MEM_stage_inst_dmem_n5620, MEM_stage_inst_dmem_n5619, MEM_stage_inst_dmem_n5618, MEM_stage_inst_dmem_n5617, MEM_stage_inst_dmem_n5616, MEM_stage_inst_dmem_n5615, MEM_stage_inst_dmem_n5614, MEM_stage_inst_dmem_n5613, MEM_stage_inst_dmem_n5612, MEM_stage_inst_dmem_n5611, MEM_stage_inst_dmem_n5610, MEM_stage_inst_dmem_n5609, MEM_stage_inst_dmem_n5608, MEM_stage_inst_dmem_n5607, MEM_stage_inst_dmem_n5606, MEM_stage_inst_dmem_n5605, MEM_stage_inst_dmem_n5604, MEM_stage_inst_dmem_n5603, MEM_stage_inst_dmem_n5602, MEM_stage_inst_dmem_n5601, MEM_stage_inst_dmem_n5600, MEM_stage_inst_dmem_n5599, MEM_stage_inst_dmem_n5598, MEM_stage_inst_dmem_n5597, MEM_stage_inst_dmem_n5596, MEM_stage_inst_dmem_n5595, MEM_stage_inst_dmem_n5594, MEM_stage_inst_dmem_n5593, MEM_stage_inst_dmem_n5592, MEM_stage_inst_dmem_n5591, MEM_stage_inst_dmem_n5590, MEM_stage_inst_dmem_n5589, MEM_stage_inst_dmem_n5588, MEM_stage_inst_dmem_n5587, MEM_stage_inst_dmem_n5586, MEM_stage_inst_dmem_n5585, MEM_stage_inst_dmem_n5584, MEM_stage_inst_dmem_n5583, MEM_stage_inst_dmem_n5582, MEM_stage_inst_dmem_n5581, MEM_stage_inst_dmem_n5580, MEM_stage_inst_dmem_n5579, MEM_stage_inst_dmem_n5578, MEM_stage_inst_dmem_n5577, MEM_stage_inst_dmem_n5576, MEM_stage_inst_dmem_n5575, MEM_stage_inst_dmem_n5574, MEM_stage_inst_dmem_n5573, MEM_stage_inst_dmem_n5572, MEM_stage_inst_dmem_n5571, MEM_stage_inst_dmem_n5570, MEM_stage_inst_dmem_n5569, MEM_stage_inst_dmem_n5568, MEM_stage_inst_dmem_n5567, MEM_stage_inst_dmem_n5566, MEM_stage_inst_dmem_n5565, MEM_stage_inst_dmem_n5564, MEM_stage_inst_dmem_n5563, MEM_stage_inst_dmem_n5562, MEM_stage_inst_dmem_n5561, MEM_stage_inst_dmem_n5560, MEM_stage_inst_dmem_n5559, MEM_stage_inst_dmem_n5558, MEM_stage_inst_dmem_n5557, MEM_stage_inst_dmem_n5556, MEM_stage_inst_dmem_n5555, MEM_stage_inst_dmem_n5554, MEM_stage_inst_dmem_n5553, MEM_stage_inst_dmem_n5552, MEM_stage_inst_dmem_n5551, MEM_stage_inst_dmem_n5550, MEM_stage_inst_dmem_n5549, MEM_stage_inst_dmem_n5548, MEM_stage_inst_dmem_n5547, MEM_stage_inst_dmem_n5546, MEM_stage_inst_dmem_n5545, MEM_stage_inst_dmem_n5544, MEM_stage_inst_dmem_n5543, MEM_stage_inst_dmem_n5542, MEM_stage_inst_dmem_n5541, MEM_stage_inst_dmem_n5540, MEM_stage_inst_dmem_n5539, MEM_stage_inst_dmem_n5538, MEM_stage_inst_dmem_n5537, MEM_stage_inst_dmem_n5536, MEM_stage_inst_dmem_n5535, MEM_stage_inst_dmem_n5534, MEM_stage_inst_dmem_n5533, MEM_stage_inst_dmem_n5532, MEM_stage_inst_dmem_n5531, MEM_stage_inst_dmem_n5530, MEM_stage_inst_dmem_n5529, MEM_stage_inst_dmem_n5528, MEM_stage_inst_dmem_n5527, MEM_stage_inst_dmem_n5526, MEM_stage_inst_dmem_n5525, MEM_stage_inst_dmem_n5524, MEM_stage_inst_dmem_n5523, MEM_stage_inst_dmem_n5522, MEM_stage_inst_dmem_n5521, MEM_stage_inst_dmem_n5520, MEM_stage_inst_dmem_n5519, MEM_stage_inst_dmem_n5518, MEM_stage_inst_dmem_n5517, MEM_stage_inst_dmem_n5516, MEM_stage_inst_dmem_n5515, MEM_stage_inst_dmem_n5514, MEM_stage_inst_dmem_n5513, MEM_stage_inst_dmem_n5512, MEM_stage_inst_dmem_n5511, MEM_stage_inst_dmem_n5510, MEM_stage_inst_dmem_n5509, MEM_stage_inst_dmem_n5508, MEM_stage_inst_dmem_n5507, MEM_stage_inst_dmem_n5506, MEM_stage_inst_dmem_n5505, MEM_stage_inst_dmem_n5504, MEM_stage_inst_dmem_n5503, MEM_stage_inst_dmem_n5502, MEM_stage_inst_dmem_n5501, MEM_stage_inst_dmem_n5500, MEM_stage_inst_dmem_n5499, MEM_stage_inst_dmem_n5498, MEM_stage_inst_dmem_n5497, MEM_stage_inst_dmem_n5496, MEM_stage_inst_dmem_n5495, MEM_stage_inst_dmem_n5494, MEM_stage_inst_dmem_n5493, MEM_stage_inst_dmem_n5492, MEM_stage_inst_dmem_n5491, MEM_stage_inst_dmem_n5490, MEM_stage_inst_dmem_n5489, MEM_stage_inst_dmem_n5488, MEM_stage_inst_dmem_n5487, MEM_stage_inst_dmem_n5486, MEM_stage_inst_dmem_n5485, MEM_stage_inst_dmem_n5484, MEM_stage_inst_dmem_n5483, MEM_stage_inst_dmem_n5482, MEM_stage_inst_dmem_n5481, MEM_stage_inst_dmem_n5480, MEM_stage_inst_dmem_n5479, MEM_stage_inst_dmem_n5478, MEM_stage_inst_dmem_n5477, MEM_stage_inst_dmem_n5476, MEM_stage_inst_dmem_n5475, MEM_stage_inst_dmem_n5474, MEM_stage_inst_dmem_n5473, MEM_stage_inst_dmem_n5472, MEM_stage_inst_dmem_n5471, MEM_stage_inst_dmem_n5470, MEM_stage_inst_dmem_n5469, MEM_stage_inst_dmem_n5468, MEM_stage_inst_dmem_n5467, MEM_stage_inst_dmem_n5466, MEM_stage_inst_dmem_n5465, MEM_stage_inst_dmem_n5464, MEM_stage_inst_dmem_n5463, MEM_stage_inst_dmem_n5462, MEM_stage_inst_dmem_n5461, MEM_stage_inst_dmem_n5460, MEM_stage_inst_dmem_n5459, MEM_stage_inst_dmem_n5458, MEM_stage_inst_dmem_n5457, MEM_stage_inst_dmem_n5456, MEM_stage_inst_dmem_n5455, MEM_stage_inst_dmem_n5454, MEM_stage_inst_dmem_n5453, MEM_stage_inst_dmem_n5452, MEM_stage_inst_dmem_n5451, MEM_stage_inst_dmem_n5450, MEM_stage_inst_dmem_n5449, MEM_stage_inst_dmem_n5448, MEM_stage_inst_dmem_n5447, MEM_stage_inst_dmem_n5446, MEM_stage_inst_dmem_n5445, MEM_stage_inst_dmem_n5444, MEM_stage_inst_dmem_n5443, MEM_stage_inst_dmem_n5442, MEM_stage_inst_dmem_n5441, MEM_stage_inst_dmem_n5440, MEM_stage_inst_dmem_n5439, MEM_stage_inst_dmem_n5438, MEM_stage_inst_dmem_n5437, MEM_stage_inst_dmem_n5436, MEM_stage_inst_dmem_n5435, MEM_stage_inst_dmem_n5434, MEM_stage_inst_dmem_n5433, MEM_stage_inst_dmem_n5432, MEM_stage_inst_dmem_n5431, MEM_stage_inst_dmem_n5430, MEM_stage_inst_dmem_n5429, MEM_stage_inst_dmem_n5428, MEM_stage_inst_dmem_n5427, MEM_stage_inst_dmem_n5426, MEM_stage_inst_dmem_n5425, MEM_stage_inst_dmem_n5424, MEM_stage_inst_dmem_n5423, MEM_stage_inst_dmem_n5422, MEM_stage_inst_dmem_n5421, MEM_stage_inst_dmem_n5420, MEM_stage_inst_dmem_n5419, MEM_stage_inst_dmem_n5418, MEM_stage_inst_dmem_n5417, MEM_stage_inst_dmem_n5416, MEM_stage_inst_dmem_n5415, MEM_stage_inst_dmem_n5414, MEM_stage_inst_dmem_n5413, MEM_stage_inst_dmem_n5412, MEM_stage_inst_dmem_n5411, MEM_stage_inst_dmem_n5410, MEM_stage_inst_dmem_n5409, MEM_stage_inst_dmem_n5408, MEM_stage_inst_dmem_n5407, MEM_stage_inst_dmem_n5406, MEM_stage_inst_dmem_n5405, MEM_stage_inst_dmem_n5404, MEM_stage_inst_dmem_n5403, MEM_stage_inst_dmem_n5402, MEM_stage_inst_dmem_n5401, MEM_stage_inst_dmem_n5400, MEM_stage_inst_dmem_n5399, MEM_stage_inst_dmem_n5398, MEM_stage_inst_dmem_n5397, MEM_stage_inst_dmem_n5396, MEM_stage_inst_dmem_n5395, MEM_stage_inst_dmem_n5394, MEM_stage_inst_dmem_n5393, MEM_stage_inst_dmem_n5392, MEM_stage_inst_dmem_n5391, MEM_stage_inst_dmem_n5390, MEM_stage_inst_dmem_n5389, MEM_stage_inst_dmem_n5388, MEM_stage_inst_dmem_n5387, MEM_stage_inst_dmem_n5386, MEM_stage_inst_dmem_n5385, MEM_stage_inst_dmem_n5384, MEM_stage_inst_dmem_n5383, MEM_stage_inst_dmem_n5382, MEM_stage_inst_dmem_n5381, MEM_stage_inst_dmem_n5380, MEM_stage_inst_dmem_n5379, MEM_stage_inst_dmem_n5378, MEM_stage_inst_dmem_n5377, MEM_stage_inst_dmem_n5376, MEM_stage_inst_dmem_n5375, MEM_stage_inst_dmem_n5374, MEM_stage_inst_dmem_n5373, MEM_stage_inst_dmem_n5372, MEM_stage_inst_dmem_n5371, MEM_stage_inst_dmem_n5370, MEM_stage_inst_dmem_n5369, MEM_stage_inst_dmem_n5368, MEM_stage_inst_dmem_n5367, MEM_stage_inst_dmem_n5366, MEM_stage_inst_dmem_n5365, MEM_stage_inst_dmem_n5364, MEM_stage_inst_dmem_n5363, MEM_stage_inst_dmem_n5362, MEM_stage_inst_dmem_n5361, MEM_stage_inst_dmem_n5360, MEM_stage_inst_dmem_n5359, MEM_stage_inst_dmem_n5358, MEM_stage_inst_dmem_n5357, MEM_stage_inst_dmem_n5356, MEM_stage_inst_dmem_n5355, MEM_stage_inst_dmem_n5354, MEM_stage_inst_dmem_n5353, MEM_stage_inst_dmem_n5352, MEM_stage_inst_dmem_n5351, MEM_stage_inst_dmem_n5350, MEM_stage_inst_dmem_n5349, MEM_stage_inst_dmem_n5348, MEM_stage_inst_dmem_n5347, MEM_stage_inst_dmem_n5346, MEM_stage_inst_dmem_n5345, MEM_stage_inst_dmem_n5344, MEM_stage_inst_dmem_n5343, MEM_stage_inst_dmem_n5342, MEM_stage_inst_dmem_n5341, MEM_stage_inst_dmem_n5340, MEM_stage_inst_dmem_n5339, MEM_stage_inst_dmem_n5338, MEM_stage_inst_dmem_n5337, MEM_stage_inst_dmem_n5336, MEM_stage_inst_dmem_n5335, MEM_stage_inst_dmem_n5334, MEM_stage_inst_dmem_n5333, MEM_stage_inst_dmem_n5332, MEM_stage_inst_dmem_n5331, MEM_stage_inst_dmem_n5330, MEM_stage_inst_dmem_n5329, MEM_stage_inst_dmem_n5328, MEM_stage_inst_dmem_n5327, MEM_stage_inst_dmem_n5326, MEM_stage_inst_dmem_n5325, MEM_stage_inst_dmem_n5324, MEM_stage_inst_dmem_n5323, MEM_stage_inst_dmem_n5322, MEM_stage_inst_dmem_n5321, MEM_stage_inst_dmem_n5320, MEM_stage_inst_dmem_n5319, MEM_stage_inst_dmem_n5318, MEM_stage_inst_dmem_n5317, MEM_stage_inst_dmem_n5316, MEM_stage_inst_dmem_n5315, MEM_stage_inst_dmem_n5314, MEM_stage_inst_dmem_n5313, MEM_stage_inst_dmem_n5312, MEM_stage_inst_dmem_n5311, MEM_stage_inst_dmem_n5310, MEM_stage_inst_dmem_n5309, MEM_stage_inst_dmem_n5308, MEM_stage_inst_dmem_n5307, MEM_stage_inst_dmem_n5306, MEM_stage_inst_dmem_n5305, MEM_stage_inst_dmem_n5304, MEM_stage_inst_dmem_n5303, MEM_stage_inst_dmem_n5302, MEM_stage_inst_dmem_n5301, MEM_stage_inst_dmem_n5300, MEM_stage_inst_dmem_n5299, MEM_stage_inst_dmem_n5298, MEM_stage_inst_dmem_n5297, MEM_stage_inst_dmem_n5296, MEM_stage_inst_dmem_n5295, MEM_stage_inst_dmem_n5294, MEM_stage_inst_dmem_n5293, MEM_stage_inst_dmem_n5292, MEM_stage_inst_dmem_n5291, MEM_stage_inst_dmem_n5290, MEM_stage_inst_dmem_n5289, MEM_stage_inst_dmem_n5288, MEM_stage_inst_dmem_n5287, MEM_stage_inst_dmem_n5286, MEM_stage_inst_dmem_n5285, MEM_stage_inst_dmem_n5284, MEM_stage_inst_dmem_n5283, MEM_stage_inst_dmem_n5282, MEM_stage_inst_dmem_n5281, MEM_stage_inst_dmem_n5280, MEM_stage_inst_dmem_n5279, MEM_stage_inst_dmem_n5278, MEM_stage_inst_dmem_n5277, MEM_stage_inst_dmem_n5276, MEM_stage_inst_dmem_n5275, MEM_stage_inst_dmem_n5274, MEM_stage_inst_dmem_n5273, MEM_stage_inst_dmem_n5272, MEM_stage_inst_dmem_n5271, MEM_stage_inst_dmem_n5270, MEM_stage_inst_dmem_n5269, MEM_stage_inst_dmem_n5268, MEM_stage_inst_dmem_n5267, MEM_stage_inst_dmem_n5266, MEM_stage_inst_dmem_n5265, MEM_stage_inst_dmem_n5264, MEM_stage_inst_dmem_n5263, MEM_stage_inst_dmem_n5262, MEM_stage_inst_dmem_n5261, MEM_stage_inst_dmem_n5260, MEM_stage_inst_dmem_n5259, MEM_stage_inst_dmem_n5258, MEM_stage_inst_dmem_n5257, MEM_stage_inst_dmem_n5256, MEM_stage_inst_dmem_n5255, MEM_stage_inst_dmem_n5254, MEM_stage_inst_dmem_n5253, MEM_stage_inst_dmem_n5252, MEM_stage_inst_dmem_n5251, MEM_stage_inst_dmem_n5250, MEM_stage_inst_dmem_n5249, MEM_stage_inst_dmem_n5248, MEM_stage_inst_dmem_n5247, MEM_stage_inst_dmem_n5246, MEM_stage_inst_dmem_n5245, MEM_stage_inst_dmem_n5244, MEM_stage_inst_dmem_n5243, MEM_stage_inst_dmem_n5242, MEM_stage_inst_dmem_n5241, MEM_stage_inst_dmem_n5240, MEM_stage_inst_dmem_n5239, MEM_stage_inst_dmem_n5238, MEM_stage_inst_dmem_n5237, MEM_stage_inst_dmem_n5236, MEM_stage_inst_dmem_n5235, MEM_stage_inst_dmem_n5234, MEM_stage_inst_dmem_n5233, MEM_stage_inst_dmem_n5232, MEM_stage_inst_dmem_n5231, MEM_stage_inst_dmem_n5230, MEM_stage_inst_dmem_n5229, MEM_stage_inst_dmem_n5228, MEM_stage_inst_dmem_n5227, MEM_stage_inst_dmem_n5226, MEM_stage_inst_dmem_n5225, MEM_stage_inst_dmem_n5224, MEM_stage_inst_dmem_n5223, MEM_stage_inst_dmem_n5222, MEM_stage_inst_dmem_n5221, MEM_stage_inst_dmem_n5220, MEM_stage_inst_dmem_n5219, MEM_stage_inst_dmem_n5218, MEM_stage_inst_dmem_n5217, MEM_stage_inst_dmem_n5216, MEM_stage_inst_dmem_n5215, MEM_stage_inst_dmem_n5214, MEM_stage_inst_dmem_n5213, MEM_stage_inst_dmem_n5212, MEM_stage_inst_dmem_n5211, MEM_stage_inst_dmem_n5210, MEM_stage_inst_dmem_n5209, MEM_stage_inst_dmem_n5208, MEM_stage_inst_dmem_n5207, MEM_stage_inst_dmem_n5206, MEM_stage_inst_dmem_n5205, MEM_stage_inst_dmem_n5204, MEM_stage_inst_dmem_n5203, MEM_stage_inst_dmem_n5202, MEM_stage_inst_dmem_n5201, MEM_stage_inst_dmem_n5200, MEM_stage_inst_dmem_n5199, MEM_stage_inst_dmem_n5198, MEM_stage_inst_dmem_n5197, MEM_stage_inst_dmem_n5196, MEM_stage_inst_dmem_n5195, MEM_stage_inst_dmem_n5194, MEM_stage_inst_dmem_n5193, MEM_stage_inst_dmem_n5192, MEM_stage_inst_dmem_n5191, MEM_stage_inst_dmem_n5190, MEM_stage_inst_dmem_n5189, MEM_stage_inst_dmem_n5188, MEM_stage_inst_dmem_n5187, MEM_stage_inst_dmem_n5186, MEM_stage_inst_dmem_n5185, MEM_stage_inst_dmem_n5184, MEM_stage_inst_dmem_n5183, MEM_stage_inst_dmem_n5182, MEM_stage_inst_dmem_n5181, MEM_stage_inst_dmem_n5180, MEM_stage_inst_dmem_n5179, MEM_stage_inst_dmem_n5178, MEM_stage_inst_dmem_n5177, MEM_stage_inst_dmem_n5176, MEM_stage_inst_dmem_n5175, MEM_stage_inst_dmem_n5174, MEM_stage_inst_dmem_n5173, MEM_stage_inst_dmem_n5172, MEM_stage_inst_dmem_n5171, MEM_stage_inst_dmem_n5170, MEM_stage_inst_dmem_n5169, MEM_stage_inst_dmem_n5168, MEM_stage_inst_dmem_n5167, MEM_stage_inst_dmem_n5166, MEM_stage_inst_dmem_n5165, MEM_stage_inst_dmem_n5164, MEM_stage_inst_dmem_n5163, MEM_stage_inst_dmem_n5162, MEM_stage_inst_dmem_n5161, MEM_stage_inst_dmem_n5160, MEM_stage_inst_dmem_n5159, MEM_stage_inst_dmem_n5158, MEM_stage_inst_dmem_n5157, MEM_stage_inst_dmem_n5156, MEM_stage_inst_dmem_n5155, MEM_stage_inst_dmem_n5154, MEM_stage_inst_dmem_n5153, MEM_stage_inst_dmem_n5152, MEM_stage_inst_dmem_n5151, MEM_stage_inst_dmem_n5150, MEM_stage_inst_dmem_n5149, MEM_stage_inst_dmem_n5148, MEM_stage_inst_dmem_n5147, MEM_stage_inst_dmem_n5146, MEM_stage_inst_dmem_n5145, MEM_stage_inst_dmem_n5144, MEM_stage_inst_dmem_n5143, MEM_stage_inst_dmem_n5142, MEM_stage_inst_dmem_n5141, MEM_stage_inst_dmem_n5140, MEM_stage_inst_dmem_n5139, MEM_stage_inst_dmem_n5138, MEM_stage_inst_dmem_n5137, MEM_stage_inst_dmem_n5136, MEM_stage_inst_dmem_n5135, MEM_stage_inst_dmem_n5134, MEM_stage_inst_dmem_n5133, MEM_stage_inst_dmem_n5132, MEM_stage_inst_dmem_n5131, MEM_stage_inst_dmem_n5130, MEM_stage_inst_dmem_n5129, MEM_stage_inst_dmem_n5128, MEM_stage_inst_dmem_n5127, MEM_stage_inst_dmem_n5126, MEM_stage_inst_dmem_n5125, MEM_stage_inst_dmem_n5124, MEM_stage_inst_dmem_n5123, MEM_stage_inst_dmem_n5122, MEM_stage_inst_dmem_n5121, MEM_stage_inst_dmem_n5120, MEM_stage_inst_dmem_n5119, MEM_stage_inst_dmem_n5118, MEM_stage_inst_dmem_n5117, MEM_stage_inst_dmem_n5116, MEM_stage_inst_dmem_n5115, MEM_stage_inst_dmem_n5114, MEM_stage_inst_dmem_n5113, MEM_stage_inst_dmem_n5112, MEM_stage_inst_dmem_n5111, MEM_stage_inst_dmem_n5110, MEM_stage_inst_dmem_n5109, MEM_stage_inst_dmem_n5108, MEM_stage_inst_dmem_n5107, MEM_stage_inst_dmem_n5106, MEM_stage_inst_dmem_n5105, MEM_stage_inst_dmem_n5104, MEM_stage_inst_dmem_n5103, MEM_stage_inst_dmem_n5102, MEM_stage_inst_dmem_n5101, MEM_stage_inst_dmem_n5100, MEM_stage_inst_dmem_n5099, MEM_stage_inst_dmem_n5098, MEM_stage_inst_dmem_n5097, MEM_stage_inst_dmem_n5096, MEM_stage_inst_dmem_n5095, MEM_stage_inst_dmem_n5094, MEM_stage_inst_dmem_n5093, MEM_stage_inst_dmem_n5092, MEM_stage_inst_dmem_n5091, MEM_stage_inst_dmem_n5090, MEM_stage_inst_dmem_n5089, MEM_stage_inst_dmem_n5088, MEM_stage_inst_dmem_n5087, MEM_stage_inst_dmem_n5086, MEM_stage_inst_dmem_n5085, MEM_stage_inst_dmem_n5084, MEM_stage_inst_dmem_n5083, MEM_stage_inst_dmem_n5082, MEM_stage_inst_dmem_n5081, MEM_stage_inst_dmem_n5080, MEM_stage_inst_dmem_n5079, MEM_stage_inst_dmem_n5078, MEM_stage_inst_dmem_n5077, MEM_stage_inst_dmem_n5076, MEM_stage_inst_dmem_n5075, MEM_stage_inst_dmem_n5074, MEM_stage_inst_dmem_n5073, MEM_stage_inst_dmem_n5072, MEM_stage_inst_dmem_n5071, MEM_stage_inst_dmem_n5070, MEM_stage_inst_dmem_n5069, MEM_stage_inst_dmem_n5068, MEM_stage_inst_dmem_n5067, MEM_stage_inst_dmem_n5066, MEM_stage_inst_dmem_n5065, MEM_stage_inst_dmem_n5064, MEM_stage_inst_dmem_n5063, MEM_stage_inst_dmem_n5062, MEM_stage_inst_dmem_n5061, MEM_stage_inst_dmem_n5060, MEM_stage_inst_dmem_n5059, MEM_stage_inst_dmem_n5058, MEM_stage_inst_dmem_n5057, MEM_stage_inst_dmem_n5056, MEM_stage_inst_dmem_n5055, MEM_stage_inst_dmem_n5054, MEM_stage_inst_dmem_n5053, MEM_stage_inst_dmem_n5052, MEM_stage_inst_dmem_n5051, MEM_stage_inst_dmem_n5050, MEM_stage_inst_dmem_n5049, MEM_stage_inst_dmem_n5048, MEM_stage_inst_dmem_n5047, MEM_stage_inst_dmem_n5046, MEM_stage_inst_dmem_n5045, MEM_stage_inst_dmem_n5044, MEM_stage_inst_dmem_n5043, MEM_stage_inst_dmem_n5042, MEM_stage_inst_dmem_n5041, MEM_stage_inst_dmem_n5040, MEM_stage_inst_dmem_n5039, MEM_stage_inst_dmem_n5038, MEM_stage_inst_dmem_n5037, MEM_stage_inst_dmem_n5036, MEM_stage_inst_dmem_n5035, MEM_stage_inst_dmem_n5034, MEM_stage_inst_dmem_n5033, MEM_stage_inst_dmem_n5032, MEM_stage_inst_dmem_n5031, MEM_stage_inst_dmem_n5030, MEM_stage_inst_dmem_n5029, MEM_stage_inst_dmem_n5028, MEM_stage_inst_dmem_n5027, MEM_stage_inst_dmem_n5026, MEM_stage_inst_dmem_n5025, MEM_stage_inst_dmem_n5024, MEM_stage_inst_dmem_n5023, MEM_stage_inst_dmem_n5022, MEM_stage_inst_dmem_n5021, MEM_stage_inst_dmem_n5020, MEM_stage_inst_dmem_n5019, MEM_stage_inst_dmem_n5018, MEM_stage_inst_dmem_n5017, MEM_stage_inst_dmem_n5016, MEM_stage_inst_dmem_n5015, MEM_stage_inst_dmem_n5014, MEM_stage_inst_dmem_n5013, MEM_stage_inst_dmem_n5012, MEM_stage_inst_dmem_n5011, MEM_stage_inst_dmem_n5010, MEM_stage_inst_dmem_n5009, MEM_stage_inst_dmem_n5008, MEM_stage_inst_dmem_n5007, MEM_stage_inst_dmem_n5006, MEM_stage_inst_dmem_n5005, MEM_stage_inst_dmem_n5004, MEM_stage_inst_dmem_n5003, MEM_stage_inst_dmem_n5002, MEM_stage_inst_dmem_n5001, MEM_stage_inst_dmem_n5000, MEM_stage_inst_dmem_n4999, MEM_stage_inst_dmem_n4998, MEM_stage_inst_dmem_n4997, MEM_stage_inst_dmem_n4996, MEM_stage_inst_dmem_n4995, MEM_stage_inst_dmem_n4994, MEM_stage_inst_dmem_n4993, MEM_stage_inst_dmem_n4992, MEM_stage_inst_dmem_n4991, MEM_stage_inst_dmem_n4990, MEM_stage_inst_dmem_n4989, MEM_stage_inst_dmem_n4988, MEM_stage_inst_dmem_n4987, MEM_stage_inst_dmem_n4986, MEM_stage_inst_dmem_n4985, MEM_stage_inst_dmem_n4984, MEM_stage_inst_dmem_n4983, MEM_stage_inst_dmem_n4982, MEM_stage_inst_dmem_n4981, MEM_stage_inst_dmem_n4980, MEM_stage_inst_dmem_n4979, MEM_stage_inst_dmem_n4978, MEM_stage_inst_dmem_n4977, MEM_stage_inst_dmem_n4976, MEM_stage_inst_dmem_n4975, MEM_stage_inst_dmem_n4974, MEM_stage_inst_dmem_n4973, MEM_stage_inst_dmem_n4972, MEM_stage_inst_dmem_n4971, MEM_stage_inst_dmem_n4970, MEM_stage_inst_dmem_n4969, MEM_stage_inst_dmem_n4968, MEM_stage_inst_dmem_n4967, MEM_stage_inst_dmem_n4966, MEM_stage_inst_dmem_n4965, MEM_stage_inst_dmem_n4964, MEM_stage_inst_dmem_n4963, MEM_stage_inst_dmem_n4962, MEM_stage_inst_dmem_n4961, MEM_stage_inst_dmem_n4960, MEM_stage_inst_dmem_n4959, MEM_stage_inst_dmem_n4958, MEM_stage_inst_dmem_n4957, MEM_stage_inst_dmem_n4956, MEM_stage_inst_dmem_n4955, MEM_stage_inst_dmem_n4954, MEM_stage_inst_dmem_n4953, MEM_stage_inst_dmem_n4952, MEM_stage_inst_dmem_n4951, MEM_stage_inst_dmem_n4950, MEM_stage_inst_dmem_n4949, MEM_stage_inst_dmem_n4948, MEM_stage_inst_dmem_n4947, MEM_stage_inst_dmem_n4946, MEM_stage_inst_dmem_n4945, MEM_stage_inst_dmem_n4944, MEM_stage_inst_dmem_n4943, MEM_stage_inst_dmem_n4942, MEM_stage_inst_dmem_n4941, MEM_stage_inst_dmem_n4940, MEM_stage_inst_dmem_n4939, MEM_stage_inst_dmem_n4938, MEM_stage_inst_dmem_n4937, MEM_stage_inst_dmem_n4936, MEM_stage_inst_dmem_n4935, MEM_stage_inst_dmem_n4934, MEM_stage_inst_dmem_n4933, MEM_stage_inst_dmem_n4932, MEM_stage_inst_dmem_n4931, MEM_stage_inst_dmem_n4930, MEM_stage_inst_dmem_n4929, MEM_stage_inst_dmem_n4928, MEM_stage_inst_dmem_n4927, MEM_stage_inst_dmem_n4926, MEM_stage_inst_dmem_n4925, MEM_stage_inst_dmem_n4924, MEM_stage_inst_dmem_n4923, MEM_stage_inst_dmem_n4922, MEM_stage_inst_dmem_n4921, MEM_stage_inst_dmem_n4920, MEM_stage_inst_dmem_n4919, MEM_stage_inst_dmem_n4918, MEM_stage_inst_dmem_n4917, MEM_stage_inst_dmem_n4916, MEM_stage_inst_dmem_n4915, MEM_stage_inst_dmem_n4914, MEM_stage_inst_dmem_n4913, MEM_stage_inst_dmem_n4912, MEM_stage_inst_dmem_n4911, MEM_stage_inst_dmem_n4910, MEM_stage_inst_dmem_n4909, MEM_stage_inst_dmem_n4908, MEM_stage_inst_dmem_n4907, MEM_stage_inst_dmem_n4906, MEM_stage_inst_dmem_n4905, MEM_stage_inst_dmem_n4904, MEM_stage_inst_dmem_n4903, MEM_stage_inst_dmem_n4902, MEM_stage_inst_dmem_n4901, MEM_stage_inst_dmem_n4900, MEM_stage_inst_dmem_n4899, MEM_stage_inst_dmem_n4898, MEM_stage_inst_dmem_n4897, MEM_stage_inst_dmem_n4896, MEM_stage_inst_dmem_n4895, MEM_stage_inst_dmem_n4894, MEM_stage_inst_dmem_n4893, MEM_stage_inst_dmem_n4892, MEM_stage_inst_dmem_n4891, MEM_stage_inst_dmem_n4890, MEM_stage_inst_dmem_n4889, MEM_stage_inst_dmem_n4888, MEM_stage_inst_dmem_n4887, MEM_stage_inst_dmem_n4886, MEM_stage_inst_dmem_n4885, MEM_stage_inst_dmem_n4884, MEM_stage_inst_dmem_n4883, MEM_stage_inst_dmem_n4882, MEM_stage_inst_dmem_n4881, MEM_stage_inst_dmem_n4880, MEM_stage_inst_dmem_n4879, MEM_stage_inst_dmem_n4878, MEM_stage_inst_dmem_n4877, MEM_stage_inst_dmem_n4876, MEM_stage_inst_dmem_n4875, MEM_stage_inst_dmem_n4874, MEM_stage_inst_dmem_n4873, MEM_stage_inst_dmem_n4872, MEM_stage_inst_dmem_n4871, MEM_stage_inst_dmem_n4870, MEM_stage_inst_dmem_n4869, MEM_stage_inst_dmem_n4868, MEM_stage_inst_dmem_n4867, MEM_stage_inst_dmem_n4866, MEM_stage_inst_dmem_n4865, MEM_stage_inst_dmem_n4864, MEM_stage_inst_dmem_n4863, MEM_stage_inst_dmem_n4862, MEM_stage_inst_dmem_n4861, MEM_stage_inst_dmem_n4860, MEM_stage_inst_dmem_n4859, MEM_stage_inst_dmem_n4858, MEM_stage_inst_dmem_n4857, MEM_stage_inst_dmem_n4856, MEM_stage_inst_dmem_n4855, MEM_stage_inst_dmem_n4854, MEM_stage_inst_dmem_n4853, MEM_stage_inst_dmem_n4852, MEM_stage_inst_dmem_n4851, MEM_stage_inst_dmem_n4850, MEM_stage_inst_dmem_n4849, MEM_stage_inst_dmem_n4848, MEM_stage_inst_dmem_n4847, MEM_stage_inst_dmem_n4846, MEM_stage_inst_dmem_n4845, MEM_stage_inst_dmem_n4844, MEM_stage_inst_dmem_n4843, MEM_stage_inst_dmem_n4842, MEM_stage_inst_dmem_n4841, MEM_stage_inst_dmem_n4840, MEM_stage_inst_dmem_n4839, MEM_stage_inst_dmem_n4838, MEM_stage_inst_dmem_n4837, MEM_stage_inst_dmem_n4836, MEM_stage_inst_dmem_n4835, MEM_stage_inst_dmem_n4834, MEM_stage_inst_dmem_n4833, MEM_stage_inst_dmem_n4832, MEM_stage_inst_dmem_n4831, MEM_stage_inst_dmem_n4830, MEM_stage_inst_dmem_n4829, MEM_stage_inst_dmem_n4828, MEM_stage_inst_dmem_n4827, MEM_stage_inst_dmem_n4826, MEM_stage_inst_dmem_n4825, MEM_stage_inst_dmem_n4824, MEM_stage_inst_dmem_n4823, MEM_stage_inst_dmem_n4822, MEM_stage_inst_dmem_n4821, MEM_stage_inst_dmem_n4820, MEM_stage_inst_dmem_n4819, MEM_stage_inst_dmem_n4818, MEM_stage_inst_dmem_n4817, MEM_stage_inst_dmem_n4816, MEM_stage_inst_dmem_n4815, MEM_stage_inst_dmem_n4814, MEM_stage_inst_dmem_n4813, MEM_stage_inst_dmem_n4812, MEM_stage_inst_dmem_n4811, MEM_stage_inst_dmem_n4810, MEM_stage_inst_dmem_n4809, MEM_stage_inst_dmem_n4808, MEM_stage_inst_dmem_n4807, MEM_stage_inst_dmem_n4806, MEM_stage_inst_dmem_n4805, MEM_stage_inst_dmem_n4804, MEM_stage_inst_dmem_n4803, MEM_stage_inst_dmem_n4802, MEM_stage_inst_dmem_n4801, MEM_stage_inst_dmem_n4800, MEM_stage_inst_dmem_n4799, MEM_stage_inst_dmem_n4798, MEM_stage_inst_dmem_n4797, MEM_stage_inst_dmem_n4796, MEM_stage_inst_dmem_n4795, MEM_stage_inst_dmem_n4794, MEM_stage_inst_dmem_n4793, MEM_stage_inst_dmem_n4792, MEM_stage_inst_dmem_n4791, MEM_stage_inst_dmem_n4790, MEM_stage_inst_dmem_n4789, MEM_stage_inst_dmem_n4788, MEM_stage_inst_dmem_n4787, MEM_stage_inst_dmem_n4786, MEM_stage_inst_dmem_n4785, MEM_stage_inst_dmem_n4784, MEM_stage_inst_dmem_n4783, MEM_stage_inst_dmem_n4782, MEM_stage_inst_dmem_n4781, MEM_stage_inst_dmem_n4780, MEM_stage_inst_dmem_n4779, MEM_stage_inst_dmem_n4778, MEM_stage_inst_dmem_n4777, MEM_stage_inst_dmem_n4776, MEM_stage_inst_dmem_n4775, MEM_stage_inst_dmem_n4774, MEM_stage_inst_dmem_n4773, MEM_stage_inst_dmem_n4772, MEM_stage_inst_dmem_n4771, MEM_stage_inst_dmem_n4770, MEM_stage_inst_dmem_n4769, MEM_stage_inst_dmem_n4768, MEM_stage_inst_dmem_n4767, MEM_stage_inst_dmem_n4766, MEM_stage_inst_dmem_n4765, MEM_stage_inst_dmem_n4764, MEM_stage_inst_dmem_n4763, MEM_stage_inst_dmem_n4762, MEM_stage_inst_dmem_n4761, MEM_stage_inst_dmem_n4760, MEM_stage_inst_dmem_n4759, MEM_stage_inst_dmem_n4758, MEM_stage_inst_dmem_n4757, MEM_stage_inst_dmem_n4756, MEM_stage_inst_dmem_n4755, MEM_stage_inst_dmem_n4754, MEM_stage_inst_dmem_n4753, MEM_stage_inst_dmem_n4752, MEM_stage_inst_dmem_n4751, MEM_stage_inst_dmem_n4750, MEM_stage_inst_dmem_n4749, MEM_stage_inst_dmem_n4748, MEM_stage_inst_dmem_n4747, MEM_stage_inst_dmem_n4746, MEM_stage_inst_dmem_n4745, MEM_stage_inst_dmem_n4744, MEM_stage_inst_dmem_n4743, MEM_stage_inst_dmem_n4742, MEM_stage_inst_dmem_n4741, MEM_stage_inst_dmem_n4740, MEM_stage_inst_dmem_n4739, MEM_stage_inst_dmem_n4738, MEM_stage_inst_dmem_n4737, MEM_stage_inst_dmem_n4736, MEM_stage_inst_dmem_n4735, MEM_stage_inst_dmem_n4734, MEM_stage_inst_dmem_n4733, MEM_stage_inst_dmem_n4732, MEM_stage_inst_dmem_n4731, MEM_stage_inst_dmem_n4730, MEM_stage_inst_dmem_n4729, MEM_stage_inst_dmem_n4728, MEM_stage_inst_dmem_n4727, MEM_stage_inst_dmem_n4726, MEM_stage_inst_dmem_n4725, MEM_stage_inst_dmem_n4724, MEM_stage_inst_dmem_n4723, MEM_stage_inst_dmem_n4722, MEM_stage_inst_dmem_n4721, MEM_stage_inst_dmem_n4720, MEM_stage_inst_dmem_n4719, MEM_stage_inst_dmem_n4718, MEM_stage_inst_dmem_n4717, MEM_stage_inst_dmem_n4716, MEM_stage_inst_dmem_n4715, MEM_stage_inst_dmem_n4714, MEM_stage_inst_dmem_n4713, MEM_stage_inst_dmem_n4712, MEM_stage_inst_dmem_n4711, MEM_stage_inst_dmem_n4710, MEM_stage_inst_dmem_n4709, MEM_stage_inst_dmem_n4708, MEM_stage_inst_dmem_n4707, MEM_stage_inst_dmem_n4706, MEM_stage_inst_dmem_n4705, MEM_stage_inst_dmem_n4704, MEM_stage_inst_dmem_n4703, MEM_stage_inst_dmem_n4702, MEM_stage_inst_dmem_n4701, MEM_stage_inst_dmem_n4700, MEM_stage_inst_dmem_n4699, MEM_stage_inst_dmem_n4698, MEM_stage_inst_dmem_n4697, MEM_stage_inst_dmem_n4696, MEM_stage_inst_dmem_n4695, MEM_stage_inst_dmem_n4694, MEM_stage_inst_dmem_n4693, MEM_stage_inst_dmem_n4692, MEM_stage_inst_dmem_n4691, MEM_stage_inst_dmem_n4690, MEM_stage_inst_dmem_n4689, MEM_stage_inst_dmem_n4688, MEM_stage_inst_dmem_n4687, MEM_stage_inst_dmem_n4686, MEM_stage_inst_dmem_n4685, MEM_stage_inst_dmem_n4684, MEM_stage_inst_dmem_n4683, MEM_stage_inst_dmem_n4682, MEM_stage_inst_dmem_n4681, MEM_stage_inst_dmem_n4680, MEM_stage_inst_dmem_n4679, MEM_stage_inst_dmem_n4678, MEM_stage_inst_dmem_n4677, MEM_stage_inst_dmem_n4676, MEM_stage_inst_dmem_n4675, MEM_stage_inst_dmem_n4674, MEM_stage_inst_dmem_n4673, MEM_stage_inst_dmem_n4672, MEM_stage_inst_dmem_n4671, MEM_stage_inst_dmem_n4670, MEM_stage_inst_dmem_n4669, MEM_stage_inst_dmem_n4668, MEM_stage_inst_dmem_n4667, MEM_stage_inst_dmem_n4666, MEM_stage_inst_dmem_n4665, MEM_stage_inst_dmem_n4664, MEM_stage_inst_dmem_n4663, MEM_stage_inst_dmem_n4662, MEM_stage_inst_dmem_n4661, MEM_stage_inst_dmem_n4660, MEM_stage_inst_dmem_n4659, MEM_stage_inst_dmem_n4658, MEM_stage_inst_dmem_n4657, MEM_stage_inst_dmem_n4656, MEM_stage_inst_dmem_n4655, MEM_stage_inst_dmem_n4654, MEM_stage_inst_dmem_n4653, MEM_stage_inst_dmem_n4652, MEM_stage_inst_dmem_n4651, MEM_stage_inst_dmem_n4650, MEM_stage_inst_dmem_n4649, MEM_stage_inst_dmem_n4648, MEM_stage_inst_dmem_n4647, MEM_stage_inst_dmem_n4646, MEM_stage_inst_dmem_n4645, MEM_stage_inst_dmem_n4644, MEM_stage_inst_dmem_n4643, MEM_stage_inst_dmem_n4642, MEM_stage_inst_dmem_n4641, MEM_stage_inst_dmem_n4640, MEM_stage_inst_dmem_n4639, MEM_stage_inst_dmem_n4638, MEM_stage_inst_dmem_n4637, MEM_stage_inst_dmem_n4636, MEM_stage_inst_dmem_n4635, MEM_stage_inst_dmem_n4634, MEM_stage_inst_dmem_n4633, MEM_stage_inst_dmem_n4632, MEM_stage_inst_dmem_n4631, MEM_stage_inst_dmem_n4630, MEM_stage_inst_dmem_n4629, MEM_stage_inst_dmem_n4628, MEM_stage_inst_dmem_n4627, MEM_stage_inst_dmem_n4626, MEM_stage_inst_dmem_n4625, MEM_stage_inst_dmem_n4624, MEM_stage_inst_dmem_n4623, MEM_stage_inst_dmem_n4622, MEM_stage_inst_dmem_n4621, MEM_stage_inst_dmem_n4620, MEM_stage_inst_dmem_n4619, MEM_stage_inst_dmem_n4618, MEM_stage_inst_dmem_n4617, MEM_stage_inst_dmem_n4616, MEM_stage_inst_dmem_n4615, MEM_stage_inst_dmem_n4614, MEM_stage_inst_dmem_n4613, MEM_stage_inst_dmem_n4612, MEM_stage_inst_dmem_n4611, MEM_stage_inst_dmem_n4610, MEM_stage_inst_dmem_n4609, MEM_stage_inst_dmem_n4608, MEM_stage_inst_dmem_n4607, MEM_stage_inst_dmem_n4606, MEM_stage_inst_dmem_n4605, MEM_stage_inst_dmem_n4604, MEM_stage_inst_dmem_n4603, MEM_stage_inst_dmem_n4602, MEM_stage_inst_dmem_n4601, MEM_stage_inst_dmem_n4600, MEM_stage_inst_dmem_n4599, MEM_stage_inst_dmem_n4598, MEM_stage_inst_dmem_n4597, MEM_stage_inst_dmem_n4596, MEM_stage_inst_dmem_n4595, MEM_stage_inst_dmem_n4594, MEM_stage_inst_dmem_n4593, MEM_stage_inst_dmem_n4592, MEM_stage_inst_dmem_n4591, MEM_stage_inst_dmem_n4590, MEM_stage_inst_dmem_n4589, MEM_stage_inst_dmem_n4588, MEM_stage_inst_dmem_n4587, MEM_stage_inst_dmem_n4586, MEM_stage_inst_dmem_n4585, MEM_stage_inst_dmem_n4584, MEM_stage_inst_dmem_n4583, MEM_stage_inst_dmem_n4582, MEM_stage_inst_dmem_n4581, MEM_stage_inst_dmem_n4580, MEM_stage_inst_dmem_n4579, MEM_stage_inst_dmem_n4578, MEM_stage_inst_dmem_n4577, MEM_stage_inst_dmem_n4576, MEM_stage_inst_dmem_n4575, MEM_stage_inst_dmem_n4574, MEM_stage_inst_dmem_n4573, MEM_stage_inst_dmem_n4572, MEM_stage_inst_dmem_n4571, MEM_stage_inst_dmem_n4570, MEM_stage_inst_dmem_n4569, MEM_stage_inst_dmem_n4568, MEM_stage_inst_dmem_n4567, MEM_stage_inst_dmem_n4566, MEM_stage_inst_dmem_n4565, MEM_stage_inst_dmem_n4564, MEM_stage_inst_dmem_n4563, MEM_stage_inst_dmem_n4562, MEM_stage_inst_dmem_n4561, MEM_stage_inst_dmem_n4560, MEM_stage_inst_dmem_n4559, MEM_stage_inst_dmem_n4558, MEM_stage_inst_dmem_n4557, MEM_stage_inst_dmem_n4556, MEM_stage_inst_dmem_n4555, MEM_stage_inst_dmem_n4554, MEM_stage_inst_dmem_n4553, MEM_stage_inst_dmem_n4552, MEM_stage_inst_dmem_n4551, MEM_stage_inst_dmem_n4550, MEM_stage_inst_dmem_n4549, MEM_stage_inst_dmem_n4548, MEM_stage_inst_dmem_n4547, MEM_stage_inst_dmem_n4546, MEM_stage_inst_dmem_n4545, MEM_stage_inst_dmem_n4544, MEM_stage_inst_dmem_n4543, MEM_stage_inst_dmem_n4542, MEM_stage_inst_dmem_n4541, MEM_stage_inst_dmem_n4540, MEM_stage_inst_dmem_n4539, MEM_stage_inst_dmem_n4538, MEM_stage_inst_dmem_n4537, MEM_stage_inst_dmem_n4536, MEM_stage_inst_dmem_n4535, MEM_stage_inst_dmem_n4534, MEM_stage_inst_dmem_n4533, MEM_stage_inst_dmem_n4532, MEM_stage_inst_dmem_n4531, MEM_stage_inst_dmem_n4530, MEM_stage_inst_dmem_n4529, MEM_stage_inst_dmem_n4528, MEM_stage_inst_dmem_n4527, MEM_stage_inst_dmem_n4526, MEM_stage_inst_dmem_n4525, MEM_stage_inst_dmem_n4524, MEM_stage_inst_dmem_n4523, MEM_stage_inst_dmem_n4522, MEM_stage_inst_dmem_n4521, MEM_stage_inst_dmem_n4520, MEM_stage_inst_dmem_n4519, MEM_stage_inst_dmem_n4518, MEM_stage_inst_dmem_n4517, MEM_stage_inst_dmem_n4516, MEM_stage_inst_dmem_n4515, MEM_stage_inst_dmem_n4514, MEM_stage_inst_dmem_n4513, MEM_stage_inst_dmem_n4512, MEM_stage_inst_dmem_n4511, MEM_stage_inst_dmem_n4510, MEM_stage_inst_dmem_n4509, MEM_stage_inst_dmem_n4508, MEM_stage_inst_dmem_n4507, MEM_stage_inst_dmem_n4506, MEM_stage_inst_dmem_n4505, MEM_stage_inst_dmem_n4504, MEM_stage_inst_dmem_n4503, MEM_stage_inst_dmem_n4502, MEM_stage_inst_dmem_n4501, MEM_stage_inst_dmem_n4500, MEM_stage_inst_dmem_n4499, MEM_stage_inst_dmem_n4498, MEM_stage_inst_dmem_n4497, MEM_stage_inst_dmem_n4496, MEM_stage_inst_dmem_n4495, MEM_stage_inst_dmem_n4494, MEM_stage_inst_dmem_n4493, MEM_stage_inst_dmem_n4492, MEM_stage_inst_dmem_n4491, MEM_stage_inst_dmem_n4490, MEM_stage_inst_dmem_n4489, MEM_stage_inst_dmem_n4488, MEM_stage_inst_dmem_n4487, MEM_stage_inst_dmem_n4486, MEM_stage_inst_dmem_n4485, MEM_stage_inst_dmem_n4484, MEM_stage_inst_dmem_n4483, MEM_stage_inst_dmem_n4482, MEM_stage_inst_dmem_n4481, MEM_stage_inst_dmem_n4480, MEM_stage_inst_dmem_n4479, MEM_stage_inst_dmem_n4478, MEM_stage_inst_dmem_n4477, MEM_stage_inst_dmem_n4476, MEM_stage_inst_dmem_n4475, MEM_stage_inst_dmem_n4474, MEM_stage_inst_dmem_n4473, MEM_stage_inst_dmem_n4472, MEM_stage_inst_dmem_n4471, MEM_stage_inst_dmem_n4470, MEM_stage_inst_dmem_n4469, MEM_stage_inst_dmem_n4468, MEM_stage_inst_dmem_n4467, MEM_stage_inst_dmem_n4466, MEM_stage_inst_dmem_n4465, MEM_stage_inst_dmem_n4464, MEM_stage_inst_dmem_n4463, MEM_stage_inst_dmem_n4462, MEM_stage_inst_dmem_n4461, MEM_stage_inst_dmem_n4460, MEM_stage_inst_dmem_n4459, MEM_stage_inst_dmem_n4458, MEM_stage_inst_dmem_n4457, MEM_stage_inst_dmem_n4456, MEM_stage_inst_dmem_n4455, MEM_stage_inst_dmem_n4454, MEM_stage_inst_dmem_n4453, MEM_stage_inst_dmem_n4452, MEM_stage_inst_dmem_n4451, MEM_stage_inst_dmem_n4450, MEM_stage_inst_dmem_n4449, MEM_stage_inst_dmem_n4448, MEM_stage_inst_dmem_n4447, MEM_stage_inst_dmem_n4446, MEM_stage_inst_dmem_n4445, MEM_stage_inst_dmem_n4444, MEM_stage_inst_dmem_n4443, MEM_stage_inst_dmem_n4442, MEM_stage_inst_dmem_n4441, MEM_stage_inst_dmem_n4440, MEM_stage_inst_dmem_n4439, MEM_stage_inst_dmem_n4438, MEM_stage_inst_dmem_n4437, MEM_stage_inst_dmem_n4436, MEM_stage_inst_dmem_n4435, MEM_stage_inst_dmem_n4434, MEM_stage_inst_dmem_n4433, MEM_stage_inst_dmem_n4432, MEM_stage_inst_dmem_n4431, MEM_stage_inst_dmem_n4430, MEM_stage_inst_dmem_n4429, MEM_stage_inst_dmem_n4428, MEM_stage_inst_dmem_n4427, MEM_stage_inst_dmem_n4426, MEM_stage_inst_dmem_n4425, MEM_stage_inst_dmem_n4424, MEM_stage_inst_dmem_n4423, MEM_stage_inst_dmem_n4422, MEM_stage_inst_dmem_n4421, MEM_stage_inst_dmem_n4420, MEM_stage_inst_dmem_n4419, MEM_stage_inst_dmem_n4418, MEM_stage_inst_dmem_n4417, MEM_stage_inst_dmem_n4416, MEM_stage_inst_dmem_n4415, MEM_stage_inst_dmem_n4414, MEM_stage_inst_dmem_n4413, MEM_stage_inst_dmem_n4412, MEM_stage_inst_dmem_n4411, MEM_stage_inst_dmem_n4410, MEM_stage_inst_dmem_n4409, MEM_stage_inst_dmem_n4408, MEM_stage_inst_dmem_n4407, MEM_stage_inst_dmem_n4406, MEM_stage_inst_dmem_n4405, MEM_stage_inst_dmem_n4404, MEM_stage_inst_dmem_n4403, MEM_stage_inst_dmem_n4402, MEM_stage_inst_dmem_n4401, MEM_stage_inst_dmem_n4400, MEM_stage_inst_dmem_n4399, MEM_stage_inst_dmem_n4398, MEM_stage_inst_dmem_n4397, MEM_stage_inst_dmem_n4396, MEM_stage_inst_dmem_n4395, MEM_stage_inst_dmem_n4394, MEM_stage_inst_dmem_n4393, MEM_stage_inst_dmem_n4392, MEM_stage_inst_dmem_n4391, MEM_stage_inst_dmem_n4390, MEM_stage_inst_dmem_n4389, MEM_stage_inst_dmem_n4388, MEM_stage_inst_dmem_n4387, MEM_stage_inst_dmem_n4386, MEM_stage_inst_dmem_n4385, MEM_stage_inst_dmem_n4384, MEM_stage_inst_dmem_n4383, MEM_stage_inst_dmem_n4382, MEM_stage_inst_dmem_n4381, MEM_stage_inst_dmem_n4380, MEM_stage_inst_dmem_n4379, MEM_stage_inst_dmem_n4378, MEM_stage_inst_dmem_n4377, MEM_stage_inst_dmem_n4376, MEM_stage_inst_dmem_n4375, MEM_stage_inst_dmem_n4374, MEM_stage_inst_dmem_n4373, MEM_stage_inst_dmem_n4372, MEM_stage_inst_dmem_n4371, MEM_stage_inst_dmem_n4370, MEM_stage_inst_dmem_n4369, MEM_stage_inst_dmem_n4368, MEM_stage_inst_dmem_n4367, MEM_stage_inst_dmem_n4366, MEM_stage_inst_dmem_n4365, MEM_stage_inst_dmem_n4364, MEM_stage_inst_dmem_n4363, MEM_stage_inst_dmem_n4362, MEM_stage_inst_dmem_n4361, MEM_stage_inst_dmem_n4360, MEM_stage_inst_dmem_n4359, MEM_stage_inst_dmem_n4358, MEM_stage_inst_dmem_n4357, MEM_stage_inst_dmem_n4356, MEM_stage_inst_dmem_n4355, MEM_stage_inst_dmem_n4354, MEM_stage_inst_dmem_n4353, MEM_stage_inst_dmem_n4352, MEM_stage_inst_dmem_n4351, MEM_stage_inst_dmem_n4350, MEM_stage_inst_dmem_n4349, MEM_stage_inst_dmem_n4348, MEM_stage_inst_dmem_n4347, MEM_stage_inst_dmem_n4346, MEM_stage_inst_dmem_n4345, MEM_stage_inst_dmem_n4344, MEM_stage_inst_dmem_n4343, MEM_stage_inst_dmem_n4342, MEM_stage_inst_dmem_n4341, MEM_stage_inst_dmem_n4340, MEM_stage_inst_dmem_n4339, MEM_stage_inst_dmem_n4338, MEM_stage_inst_dmem_n4337, MEM_stage_inst_dmem_n4336, MEM_stage_inst_dmem_n4335, MEM_stage_inst_dmem_n4334, MEM_stage_inst_dmem_n4333, MEM_stage_inst_dmem_n4332, MEM_stage_inst_dmem_n4331, MEM_stage_inst_dmem_n4330, MEM_stage_inst_dmem_n4329, MEM_stage_inst_dmem_n4328, MEM_stage_inst_dmem_n4327, MEM_stage_inst_dmem_n4326, MEM_stage_inst_dmem_n4325, MEM_stage_inst_dmem_n4324, MEM_stage_inst_dmem_n4323, MEM_stage_inst_dmem_n4322, MEM_stage_inst_dmem_n4321, MEM_stage_inst_dmem_n4320, MEM_stage_inst_dmem_n4319, MEM_stage_inst_dmem_n4318, MEM_stage_inst_dmem_n4317, MEM_stage_inst_dmem_n4316, MEM_stage_inst_dmem_n4315, MEM_stage_inst_dmem_n4314, MEM_stage_inst_dmem_n4313, MEM_stage_inst_dmem_n4312, MEM_stage_inst_dmem_n4311, MEM_stage_inst_dmem_n4310, MEM_stage_inst_dmem_n4309, MEM_stage_inst_dmem_n4308, MEM_stage_inst_dmem_n4307, MEM_stage_inst_dmem_n4306, MEM_stage_inst_dmem_n4305, MEM_stage_inst_dmem_n4304, MEM_stage_inst_dmem_n4303, MEM_stage_inst_dmem_n4302, MEM_stage_inst_dmem_n4301, MEM_stage_inst_dmem_n4300, MEM_stage_inst_dmem_n4299, MEM_stage_inst_dmem_n4298, MEM_stage_inst_dmem_n4297, MEM_stage_inst_dmem_n4296, MEM_stage_inst_dmem_n4295, MEM_stage_inst_dmem_n4294, MEM_stage_inst_dmem_n4293, MEM_stage_inst_dmem_n4292, MEM_stage_inst_dmem_n4291, MEM_stage_inst_dmem_n4290, MEM_stage_inst_dmem_n4289, MEM_stage_inst_dmem_n4288, MEM_stage_inst_dmem_n4287, MEM_stage_inst_dmem_n4286, MEM_stage_inst_dmem_n4285, MEM_stage_inst_dmem_n4284, MEM_stage_inst_dmem_n4283, MEM_stage_inst_dmem_n4282, MEM_stage_inst_dmem_n4281, MEM_stage_inst_dmem_n4280, MEM_stage_inst_dmem_n4279, MEM_stage_inst_dmem_n4278, MEM_stage_inst_dmem_n4277, MEM_stage_inst_dmem_n4276, MEM_stage_inst_dmem_n4275, MEM_stage_inst_dmem_n4274, MEM_stage_inst_dmem_n4273, MEM_stage_inst_dmem_n4272, MEM_stage_inst_dmem_n4271, MEM_stage_inst_dmem_n4270, MEM_stage_inst_dmem_n4269, MEM_stage_inst_dmem_n4268, MEM_stage_inst_dmem_n4267, MEM_stage_inst_dmem_n4266, MEM_stage_inst_dmem_n4265, MEM_stage_inst_dmem_n4264, MEM_stage_inst_dmem_n4263, MEM_stage_inst_dmem_n4262, MEM_stage_inst_dmem_n4261, MEM_stage_inst_dmem_n4260, MEM_stage_inst_dmem_n4259, MEM_stage_inst_dmem_n4258, MEM_stage_inst_dmem_n4257, MEM_stage_inst_dmem_n4256, MEM_stage_inst_dmem_n4255, MEM_stage_inst_dmem_n4254, MEM_stage_inst_dmem_n4253, MEM_stage_inst_dmem_n4252, MEM_stage_inst_dmem_n4251, MEM_stage_inst_dmem_n4250, MEM_stage_inst_dmem_n4249, MEM_stage_inst_dmem_n4248, MEM_stage_inst_dmem_n4247, MEM_stage_inst_dmem_n4246, MEM_stage_inst_dmem_n4245, MEM_stage_inst_dmem_n4244, MEM_stage_inst_dmem_n4243, MEM_stage_inst_dmem_n4242, MEM_stage_inst_dmem_n4241, MEM_stage_inst_dmem_n4240, MEM_stage_inst_dmem_n4239, MEM_stage_inst_dmem_n4238, MEM_stage_inst_dmem_n4237, MEM_stage_inst_dmem_n4236, MEM_stage_inst_dmem_n4235, MEM_stage_inst_dmem_n4234, MEM_stage_inst_dmem_n4233, MEM_stage_inst_dmem_n4232, MEM_stage_inst_dmem_n4231, MEM_stage_inst_dmem_n4230, MEM_stage_inst_dmem_n4229, MEM_stage_inst_dmem_n4228, MEM_stage_inst_dmem_n4227, MEM_stage_inst_dmem_n4226, MEM_stage_inst_dmem_n4225, MEM_stage_inst_dmem_n4224, MEM_stage_inst_dmem_n4223, MEM_stage_inst_dmem_n4222, MEM_stage_inst_dmem_n4221, MEM_stage_inst_dmem_n4220, MEM_stage_inst_dmem_n4219, MEM_stage_inst_dmem_n4218, MEM_stage_inst_dmem_n4217, MEM_stage_inst_dmem_n4216, MEM_stage_inst_dmem_n4215, MEM_stage_inst_dmem_n4214, MEM_stage_inst_dmem_n4213, MEM_stage_inst_dmem_n4212, MEM_stage_inst_dmem_n4211, MEM_stage_inst_dmem_n4210, MEM_stage_inst_dmem_n4209, MEM_stage_inst_dmem_n4208, MEM_stage_inst_dmem_n4207, MEM_stage_inst_dmem_n4206, MEM_stage_inst_dmem_n4205, MEM_stage_inst_dmem_n4204, MEM_stage_inst_dmem_n4203, MEM_stage_inst_dmem_n4202, MEM_stage_inst_dmem_n4201, MEM_stage_inst_dmem_n4200, MEM_stage_inst_dmem_n4199, MEM_stage_inst_dmem_n4198, MEM_stage_inst_dmem_n4197, MEM_stage_inst_dmem_n4196, MEM_stage_inst_dmem_n4195, MEM_stage_inst_dmem_n4194, MEM_stage_inst_dmem_n4193, MEM_stage_inst_dmem_n4192, MEM_stage_inst_dmem_n4191, MEM_stage_inst_dmem_n4190, MEM_stage_inst_dmem_n4189, MEM_stage_inst_dmem_n4188, MEM_stage_inst_dmem_n4187, MEM_stage_inst_dmem_n4186, MEM_stage_inst_dmem_n4185, MEM_stage_inst_dmem_n4184, MEM_stage_inst_dmem_n4183, MEM_stage_inst_dmem_n4182, MEM_stage_inst_dmem_n4181, MEM_stage_inst_dmem_n4180, MEM_stage_inst_dmem_n4179, MEM_stage_inst_dmem_n4178, MEM_stage_inst_dmem_n4177, MEM_stage_inst_dmem_n4176, MEM_stage_inst_dmem_n4175, MEM_stage_inst_dmem_n4174, MEM_stage_inst_dmem_n4173, MEM_stage_inst_dmem_n4172, MEM_stage_inst_dmem_n4171, MEM_stage_inst_dmem_n4170, MEM_stage_inst_dmem_n4169, MEM_stage_inst_dmem_n4168, MEM_stage_inst_dmem_n4167, MEM_stage_inst_dmem_n4166, MEM_stage_inst_dmem_n4165, MEM_stage_inst_dmem_n4164, MEM_stage_inst_dmem_n4163, MEM_stage_inst_dmem_n4162, MEM_stage_inst_dmem_n4161, MEM_stage_inst_dmem_n4160, MEM_stage_inst_dmem_n4159, MEM_stage_inst_dmem_n4158, MEM_stage_inst_dmem_n4157, MEM_stage_inst_dmem_n4156, MEM_stage_inst_dmem_n4155, MEM_stage_inst_dmem_n4154, MEM_stage_inst_dmem_n4153, MEM_stage_inst_dmem_n4152, MEM_stage_inst_dmem_n4151, MEM_stage_inst_dmem_n4150, MEM_stage_inst_dmem_n4149, MEM_stage_inst_dmem_n4148, MEM_stage_inst_dmem_n4147, MEM_stage_inst_dmem_n4146, MEM_stage_inst_dmem_n4145, MEM_stage_inst_dmem_n4144, MEM_stage_inst_dmem_n4143, MEM_stage_inst_dmem_n4142, MEM_stage_inst_dmem_n4141, MEM_stage_inst_dmem_n4140, MEM_stage_inst_dmem_n4139, MEM_stage_inst_dmem_n4138, MEM_stage_inst_dmem_n4137, MEM_stage_inst_dmem_n4136, MEM_stage_inst_dmem_n4135, MEM_stage_inst_dmem_n4134, MEM_stage_inst_dmem_n4133, MEM_stage_inst_dmem_n4132, MEM_stage_inst_dmem_n4131, MEM_stage_inst_dmem_n4130, MEM_stage_inst_dmem_n4129, MEM_stage_inst_dmem_n4128, MEM_stage_inst_dmem_n4127, MEM_stage_inst_dmem_n4126, MEM_stage_inst_dmem_n4125, MEM_stage_inst_dmem_n4124, MEM_stage_inst_dmem_n4123, MEM_stage_inst_dmem_n4122, MEM_stage_inst_dmem_n4121, MEM_stage_inst_dmem_n4120, MEM_stage_inst_dmem_n4119, MEM_stage_inst_dmem_n4118, MEM_stage_inst_dmem_n4117, MEM_stage_inst_dmem_n4116, MEM_stage_inst_dmem_n4115, MEM_stage_inst_dmem_n4114, MEM_stage_inst_dmem_n4113, MEM_stage_inst_dmem_n4112, MEM_stage_inst_dmem_n4111, MEM_stage_inst_dmem_n4110, MEM_stage_inst_dmem_n4109, MEM_stage_inst_dmem_n4108, MEM_stage_inst_dmem_n4107, MEM_stage_inst_dmem_n4106, MEM_stage_inst_dmem_n4105, MEM_stage_inst_dmem_n4104, MEM_stage_inst_dmem_n4103, MEM_stage_inst_dmem_n4102, MEM_stage_inst_dmem_n4101, MEM_stage_inst_dmem_n4100, MEM_stage_inst_dmem_n4099, MEM_stage_inst_dmem_n4098, MEM_stage_inst_dmem_n4097, MEM_stage_inst_dmem_n4096, MEM_stage_inst_dmem_n4095, MEM_stage_inst_dmem_n4094, MEM_stage_inst_dmem_n4093, MEM_stage_inst_dmem_n4092, MEM_stage_inst_dmem_n4091, MEM_stage_inst_dmem_n4090, MEM_stage_inst_dmem_n4089, MEM_stage_inst_dmem_n4088, MEM_stage_inst_dmem_n4087, MEM_stage_inst_dmem_n4086, MEM_stage_inst_dmem_n4085, MEM_stage_inst_dmem_n4084, MEM_stage_inst_dmem_n4083, MEM_stage_inst_dmem_n4082, MEM_stage_inst_dmem_n4081, MEM_stage_inst_dmem_n4080, MEM_stage_inst_dmem_n4079, MEM_stage_inst_dmem_n4078, MEM_stage_inst_dmem_n4077, MEM_stage_inst_dmem_n4076, MEM_stage_inst_dmem_n4075, MEM_stage_inst_dmem_n4074, MEM_stage_inst_dmem_n4073, MEM_stage_inst_dmem_n4072, MEM_stage_inst_dmem_n4071, MEM_stage_inst_dmem_n4070, MEM_stage_inst_dmem_n4069, MEM_stage_inst_dmem_n4068, MEM_stage_inst_dmem_n4067, MEM_stage_inst_dmem_n4066, MEM_stage_inst_dmem_n4065, MEM_stage_inst_dmem_n4064, MEM_stage_inst_dmem_n4063, MEM_stage_inst_dmem_n4062, MEM_stage_inst_dmem_n4061, MEM_stage_inst_dmem_n4060, MEM_stage_inst_dmem_n4059, MEM_stage_inst_dmem_n4058, MEM_stage_inst_dmem_n4057, MEM_stage_inst_dmem_n4056, MEM_stage_inst_dmem_n4055, MEM_stage_inst_dmem_n4054, MEM_stage_inst_dmem_n4053, MEM_stage_inst_dmem_n4052, MEM_stage_inst_dmem_n4051, MEM_stage_inst_dmem_n4050, MEM_stage_inst_dmem_n4049, MEM_stage_inst_dmem_n4048, MEM_stage_inst_dmem_n4047, MEM_stage_inst_dmem_n4046, MEM_stage_inst_dmem_n4045, MEM_stage_inst_dmem_n4044, MEM_stage_inst_dmem_n4043, MEM_stage_inst_dmem_n4042, MEM_stage_inst_dmem_n4041, MEM_stage_inst_dmem_n4040, MEM_stage_inst_dmem_n4039, MEM_stage_inst_dmem_n4038, MEM_stage_inst_dmem_n4037, MEM_stage_inst_dmem_n4036, MEM_stage_inst_dmem_n4035, MEM_stage_inst_dmem_n4034, MEM_stage_inst_dmem_n4033, MEM_stage_inst_dmem_n4032, MEM_stage_inst_dmem_n4031, MEM_stage_inst_dmem_n4030, MEM_stage_inst_dmem_n4029, MEM_stage_inst_dmem_n4028, MEM_stage_inst_dmem_n4027, MEM_stage_inst_dmem_n4026, MEM_stage_inst_dmem_n4025, MEM_stage_inst_dmem_n4024, MEM_stage_inst_dmem_n4023, MEM_stage_inst_dmem_n4022, MEM_stage_inst_dmem_n4021, MEM_stage_inst_dmem_n4020, MEM_stage_inst_dmem_n4019, MEM_stage_inst_dmem_n4018, MEM_stage_inst_dmem_n4017, MEM_stage_inst_dmem_n4016, MEM_stage_inst_dmem_n4015, MEM_stage_inst_dmem_n4014, MEM_stage_inst_dmem_n4013, MEM_stage_inst_dmem_n4012, MEM_stage_inst_dmem_n4011, MEM_stage_inst_dmem_n4010, MEM_stage_inst_dmem_n4009, MEM_stage_inst_dmem_n4008, MEM_stage_inst_dmem_n4007, MEM_stage_inst_dmem_n4006, MEM_stage_inst_dmem_n4005, MEM_stage_inst_dmem_n4004, MEM_stage_inst_dmem_n4003, MEM_stage_inst_dmem_n4002, MEM_stage_inst_dmem_n4001, MEM_stage_inst_dmem_n4000, MEM_stage_inst_dmem_n3999, MEM_stage_inst_dmem_n3998, MEM_stage_inst_dmem_n3997, MEM_stage_inst_dmem_n3996, MEM_stage_inst_dmem_n3995, MEM_stage_inst_dmem_n3994, MEM_stage_inst_dmem_n3993, MEM_stage_inst_dmem_n3992, MEM_stage_inst_dmem_n3991, MEM_stage_inst_dmem_n3990, MEM_stage_inst_dmem_n3989, MEM_stage_inst_dmem_n3988, MEM_stage_inst_dmem_n3987, MEM_stage_inst_dmem_n3986, MEM_stage_inst_dmem_n3985, MEM_stage_inst_dmem_n3984, MEM_stage_inst_dmem_n3983, MEM_stage_inst_dmem_n3982, MEM_stage_inst_dmem_n3981, MEM_stage_inst_dmem_n3980, MEM_stage_inst_dmem_n3979, MEM_stage_inst_dmem_n3978, MEM_stage_inst_dmem_n3977, MEM_stage_inst_dmem_n3976, MEM_stage_inst_dmem_n3975, MEM_stage_inst_dmem_n3974, MEM_stage_inst_dmem_n3973, MEM_stage_inst_dmem_n3972, MEM_stage_inst_dmem_n3971, MEM_stage_inst_dmem_n3970, MEM_stage_inst_dmem_n3969, MEM_stage_inst_dmem_n3968, MEM_stage_inst_dmem_n3967, MEM_stage_inst_dmem_n3966, MEM_stage_inst_dmem_n3965, MEM_stage_inst_dmem_n3964, MEM_stage_inst_dmem_n3963, MEM_stage_inst_dmem_n3962, MEM_stage_inst_dmem_n3961, MEM_stage_inst_dmem_n3960, MEM_stage_inst_dmem_n3959, MEM_stage_inst_dmem_n3958, MEM_stage_inst_dmem_n3957, MEM_stage_inst_dmem_n3956, MEM_stage_inst_dmem_n3955, MEM_stage_inst_dmem_n3954, MEM_stage_inst_dmem_n3953, MEM_stage_inst_dmem_n3952, MEM_stage_inst_dmem_n3951, MEM_stage_inst_dmem_n3950, MEM_stage_inst_dmem_n3949, MEM_stage_inst_dmem_n3948, MEM_stage_inst_dmem_n3947, MEM_stage_inst_dmem_n3946, MEM_stage_inst_dmem_n3945, MEM_stage_inst_dmem_n3944, MEM_stage_inst_dmem_n3943, MEM_stage_inst_dmem_n3942, MEM_stage_inst_dmem_n3941, MEM_stage_inst_dmem_n3940, MEM_stage_inst_dmem_n3939, MEM_stage_inst_dmem_n3938, MEM_stage_inst_dmem_n3937, MEM_stage_inst_dmem_n3936, MEM_stage_inst_dmem_n3935, MEM_stage_inst_dmem_n3934, MEM_stage_inst_dmem_n3933, MEM_stage_inst_dmem_n3932, MEM_stage_inst_dmem_n3931, MEM_stage_inst_dmem_n3930, MEM_stage_inst_dmem_n3929, MEM_stage_inst_dmem_n3928, MEM_stage_inst_dmem_n3927, MEM_stage_inst_dmem_n3926, MEM_stage_inst_dmem_n3925, MEM_stage_inst_dmem_n3924, MEM_stage_inst_dmem_n3923, MEM_stage_inst_dmem_n3922, MEM_stage_inst_dmem_n3921, MEM_stage_inst_dmem_n3920, MEM_stage_inst_dmem_n3919, MEM_stage_inst_dmem_n3918, MEM_stage_inst_dmem_n3917, MEM_stage_inst_dmem_n3916, MEM_stage_inst_dmem_n3915, MEM_stage_inst_dmem_n3914, MEM_stage_inst_dmem_n3913, MEM_stage_inst_dmem_n3912, MEM_stage_inst_dmem_n3911, MEM_stage_inst_dmem_n3910, MEM_stage_inst_dmem_n3909, MEM_stage_inst_dmem_n3908, MEM_stage_inst_dmem_n3907, MEM_stage_inst_dmem_n3906, MEM_stage_inst_dmem_n3905, MEM_stage_inst_dmem_n3904, MEM_stage_inst_dmem_n3903, MEM_stage_inst_dmem_n3902, MEM_stage_inst_dmem_n3901, MEM_stage_inst_dmem_n3900, MEM_stage_inst_dmem_n3899, MEM_stage_inst_dmem_n3898, MEM_stage_inst_dmem_n3897, MEM_stage_inst_dmem_n3896, MEM_stage_inst_dmem_n3895, MEM_stage_inst_dmem_n3894, MEM_stage_inst_dmem_n3893, MEM_stage_inst_dmem_n3892, MEM_stage_inst_dmem_n3891, MEM_stage_inst_dmem_n3890, MEM_stage_inst_dmem_n3889, MEM_stage_inst_dmem_n3888, MEM_stage_inst_dmem_n3887, MEM_stage_inst_dmem_n3886, MEM_stage_inst_dmem_n3885, MEM_stage_inst_dmem_n3884, MEM_stage_inst_dmem_n3883, MEM_stage_inst_dmem_n3882, MEM_stage_inst_dmem_n3881, MEM_stage_inst_dmem_n3880, MEM_stage_inst_dmem_n3879, MEM_stage_inst_dmem_n3878, MEM_stage_inst_dmem_n3877, MEM_stage_inst_dmem_n3876, MEM_stage_inst_dmem_n3875, MEM_stage_inst_dmem_n3874, MEM_stage_inst_dmem_n3873, MEM_stage_inst_dmem_n3872, MEM_stage_inst_dmem_n3871, MEM_stage_inst_dmem_n3870, MEM_stage_inst_dmem_n3869, MEM_stage_inst_dmem_n3868, MEM_stage_inst_dmem_n3867, MEM_stage_inst_dmem_n3866, MEM_stage_inst_dmem_n3865, MEM_stage_inst_dmem_n3864, MEM_stage_inst_dmem_n3863, MEM_stage_inst_dmem_n3862, MEM_stage_inst_dmem_n3861, MEM_stage_inst_dmem_n3860, MEM_stage_inst_dmem_n3859, MEM_stage_inst_dmem_n3858, MEM_stage_inst_dmem_n3857, MEM_stage_inst_dmem_n3856, MEM_stage_inst_dmem_n3855, MEM_stage_inst_dmem_n3854, MEM_stage_inst_dmem_n3853, MEM_stage_inst_dmem_n3852, MEM_stage_inst_dmem_n3851, MEM_stage_inst_dmem_n3850, MEM_stage_inst_dmem_n3849, MEM_stage_inst_dmem_n3848, MEM_stage_inst_dmem_n3847, MEM_stage_inst_dmem_n3846, MEM_stage_inst_dmem_n3845, MEM_stage_inst_dmem_n3844, MEM_stage_inst_dmem_n3843, MEM_stage_inst_dmem_n3842, MEM_stage_inst_dmem_n3841, MEM_stage_inst_dmem_n3840, MEM_stage_inst_dmem_n3839, MEM_stage_inst_dmem_n3838, MEM_stage_inst_dmem_n3837, MEM_stage_inst_dmem_n3836, MEM_stage_inst_dmem_n3835, MEM_stage_inst_dmem_n3834, MEM_stage_inst_dmem_n3833, MEM_stage_inst_dmem_n3832, MEM_stage_inst_dmem_n3831, MEM_stage_inst_dmem_n3830, MEM_stage_inst_dmem_n3829, MEM_stage_inst_dmem_n3828, MEM_stage_inst_dmem_n3827, MEM_stage_inst_dmem_n3826, MEM_stage_inst_dmem_n3825, MEM_stage_inst_dmem_n3824, MEM_stage_inst_dmem_n3823, MEM_stage_inst_dmem_n3822, MEM_stage_inst_dmem_n3821, MEM_stage_inst_dmem_n3820, MEM_stage_inst_dmem_n3819, MEM_stage_inst_dmem_n3818, MEM_stage_inst_dmem_n3817, MEM_stage_inst_dmem_n3816, MEM_stage_inst_dmem_n3815, MEM_stage_inst_dmem_n3814, MEM_stage_inst_dmem_n3813, MEM_stage_inst_dmem_n3812, MEM_stage_inst_dmem_n3811, MEM_stage_inst_dmem_n3810, MEM_stage_inst_dmem_n3809, MEM_stage_inst_dmem_n3808, MEM_stage_inst_dmem_n3807, MEM_stage_inst_dmem_n3806, MEM_stage_inst_dmem_n3805, MEM_stage_inst_dmem_n3804, MEM_stage_inst_dmem_n3803, MEM_stage_inst_dmem_n3802, MEM_stage_inst_dmem_n3801, MEM_stage_inst_dmem_n3800, MEM_stage_inst_dmem_n3799, MEM_stage_inst_dmem_n3798, MEM_stage_inst_dmem_n3797, MEM_stage_inst_dmem_n3796, MEM_stage_inst_dmem_n3795, MEM_stage_inst_dmem_n3794, MEM_stage_inst_dmem_n3793, MEM_stage_inst_dmem_n3792, MEM_stage_inst_dmem_n3791, MEM_stage_inst_dmem_n3790, MEM_stage_inst_dmem_n3789, MEM_stage_inst_dmem_n3788, MEM_stage_inst_dmem_n3787, MEM_stage_inst_dmem_n3786, MEM_stage_inst_dmem_n3785, MEM_stage_inst_dmem_n3784, MEM_stage_inst_dmem_n3783, MEM_stage_inst_dmem_n3782, MEM_stage_inst_dmem_n3781, MEM_stage_inst_dmem_n3780, MEM_stage_inst_dmem_n3779, MEM_stage_inst_dmem_n3778, MEM_stage_inst_dmem_n3777, MEM_stage_inst_dmem_n3776, MEM_stage_inst_dmem_n3775, MEM_stage_inst_dmem_n3774, MEM_stage_inst_dmem_n3773, MEM_stage_inst_dmem_n3772, MEM_stage_inst_dmem_n3771, MEM_stage_inst_dmem_n3770, MEM_stage_inst_dmem_n3769, MEM_stage_inst_dmem_n3768, MEM_stage_inst_dmem_n3767, MEM_stage_inst_dmem_n3766, MEM_stage_inst_dmem_n3765, MEM_stage_inst_dmem_n3764, MEM_stage_inst_dmem_n3763, MEM_stage_inst_dmem_n3762, MEM_stage_inst_dmem_n3761, MEM_stage_inst_dmem_n3760, MEM_stage_inst_dmem_n3759, MEM_stage_inst_dmem_n3758, MEM_stage_inst_dmem_n3757, MEM_stage_inst_dmem_n3756, MEM_stage_inst_dmem_n3755, MEM_stage_inst_dmem_n3754, MEM_stage_inst_dmem_n3753, MEM_stage_inst_dmem_n3752, MEM_stage_inst_dmem_n3751, MEM_stage_inst_dmem_n3750, MEM_stage_inst_dmem_n3749, MEM_stage_inst_dmem_n3748, MEM_stage_inst_dmem_n3747, MEM_stage_inst_dmem_n3746, MEM_stage_inst_dmem_n3745, MEM_stage_inst_dmem_n3744, MEM_stage_inst_dmem_n3743, MEM_stage_inst_dmem_n3742, MEM_stage_inst_dmem_n3741, MEM_stage_inst_dmem_n3740, MEM_stage_inst_dmem_n3739, MEM_stage_inst_dmem_n3738, MEM_stage_inst_dmem_n3737, MEM_stage_inst_dmem_n3736, MEM_stage_inst_dmem_n3735, MEM_stage_inst_dmem_n3734, MEM_stage_inst_dmem_n3733, MEM_stage_inst_dmem_n3732, MEM_stage_inst_dmem_n3731, MEM_stage_inst_dmem_n3730, MEM_stage_inst_dmem_n3729, MEM_stage_inst_dmem_n3728, MEM_stage_inst_dmem_n3727, MEM_stage_inst_dmem_n3726, MEM_stage_inst_dmem_n3725, MEM_stage_inst_dmem_n3724, MEM_stage_inst_dmem_n3723, MEM_stage_inst_dmem_n3722, MEM_stage_inst_dmem_n3721, MEM_stage_inst_dmem_n3720, MEM_stage_inst_dmem_n3719, MEM_stage_inst_dmem_n3718, MEM_stage_inst_dmem_n3717, MEM_stage_inst_dmem_n3716, MEM_stage_inst_dmem_n3715, MEM_stage_inst_dmem_n3714, MEM_stage_inst_dmem_n3713, MEM_stage_inst_dmem_n3712, MEM_stage_inst_dmem_n3711, MEM_stage_inst_dmem_n3710, MEM_stage_inst_dmem_n3709, MEM_stage_inst_dmem_n3708, MEM_stage_inst_dmem_n3707, MEM_stage_inst_dmem_n3706, MEM_stage_inst_dmem_n3705, MEM_stage_inst_dmem_n3704, MEM_stage_inst_dmem_n3703, MEM_stage_inst_dmem_n3702, MEM_stage_inst_dmem_n3701, MEM_stage_inst_dmem_n3700, MEM_stage_inst_dmem_n3699, MEM_stage_inst_dmem_n3698, MEM_stage_inst_dmem_n3697, MEM_stage_inst_dmem_n3696, MEM_stage_inst_dmem_n3695, MEM_stage_inst_dmem_n3694, MEM_stage_inst_dmem_n3693, MEM_stage_inst_dmem_n3692, MEM_stage_inst_dmem_n3691, MEM_stage_inst_dmem_n3690, MEM_stage_inst_dmem_n3689, MEM_stage_inst_dmem_n3688, MEM_stage_inst_dmem_n3687, MEM_stage_inst_dmem_n3686, MEM_stage_inst_dmem_n3685, MEM_stage_inst_dmem_n3684, MEM_stage_inst_dmem_n3683, MEM_stage_inst_dmem_n3682, MEM_stage_inst_dmem_n3681, MEM_stage_inst_dmem_n3680, MEM_stage_inst_dmem_n3679, MEM_stage_inst_dmem_n3678, MEM_stage_inst_dmem_n3677, MEM_stage_inst_dmem_n3676, MEM_stage_inst_dmem_n3675, MEM_stage_inst_dmem_n3674, MEM_stage_inst_dmem_n3673, MEM_stage_inst_dmem_n3672, MEM_stage_inst_dmem_n3671, MEM_stage_inst_dmem_n3670, MEM_stage_inst_dmem_n3669, MEM_stage_inst_dmem_n3668, MEM_stage_inst_dmem_n3667, MEM_stage_inst_dmem_n3666, MEM_stage_inst_dmem_n3665, MEM_stage_inst_dmem_n3664, MEM_stage_inst_dmem_n3663, MEM_stage_inst_dmem_n3662, MEM_stage_inst_dmem_n3661, MEM_stage_inst_dmem_n3660, MEM_stage_inst_dmem_n3659, MEM_stage_inst_dmem_n3658, MEM_stage_inst_dmem_n3657, MEM_stage_inst_dmem_n3656, MEM_stage_inst_dmem_n3655, MEM_stage_inst_dmem_n3654, MEM_stage_inst_dmem_n3653, MEM_stage_inst_dmem_n3652, MEM_stage_inst_dmem_n3651, MEM_stage_inst_dmem_n3650, MEM_stage_inst_dmem_n3649, MEM_stage_inst_dmem_n3648, MEM_stage_inst_dmem_n3647, MEM_stage_inst_dmem_n3646, MEM_stage_inst_dmem_n3645, MEM_stage_inst_dmem_n3644, MEM_stage_inst_dmem_n3643, MEM_stage_inst_dmem_n3642, MEM_stage_inst_dmem_n3641, MEM_stage_inst_dmem_n3640, MEM_stage_inst_dmem_n3639, MEM_stage_inst_dmem_n3638, MEM_stage_inst_dmem_n3637, MEM_stage_inst_dmem_n3636, MEM_stage_inst_dmem_n3635, MEM_stage_inst_dmem_n3634, MEM_stage_inst_dmem_n3633, MEM_stage_inst_dmem_n3632, MEM_stage_inst_dmem_n3631, MEM_stage_inst_dmem_n3630, MEM_stage_inst_dmem_n3629, MEM_stage_inst_dmem_n3628, MEM_stage_inst_dmem_n3627, MEM_stage_inst_dmem_n3626, MEM_stage_inst_dmem_n3625, MEM_stage_inst_dmem_n3624, MEM_stage_inst_dmem_n3623, MEM_stage_inst_dmem_n3622, MEM_stage_inst_dmem_n3621, MEM_stage_inst_dmem_n3620, MEM_stage_inst_dmem_n3619, MEM_stage_inst_dmem_n3618, MEM_stage_inst_dmem_n3617, MEM_stage_inst_dmem_n3616, MEM_stage_inst_dmem_n3615, MEM_stage_inst_dmem_n3614, MEM_stage_inst_dmem_n3613, MEM_stage_inst_dmem_n3612, MEM_stage_inst_dmem_n3611, MEM_stage_inst_dmem_n3610, MEM_stage_inst_dmem_n3609, MEM_stage_inst_dmem_n3608, MEM_stage_inst_dmem_n3607, MEM_stage_inst_dmem_n3606, MEM_stage_inst_dmem_n3605, MEM_stage_inst_dmem_n3604, MEM_stage_inst_dmem_n3603, MEM_stage_inst_dmem_n3602, MEM_stage_inst_dmem_n3601, MEM_stage_inst_dmem_n3600, MEM_stage_inst_dmem_n3599, MEM_stage_inst_dmem_n3598, MEM_stage_inst_dmem_n3597, MEM_stage_inst_dmem_n3596, MEM_stage_inst_dmem_n3595, MEM_stage_inst_dmem_n3594, MEM_stage_inst_dmem_n3593, MEM_stage_inst_dmem_n3592, MEM_stage_inst_dmem_n3591, MEM_stage_inst_dmem_n3590, MEM_stage_inst_dmem_n3589, MEM_stage_inst_dmem_n3588, MEM_stage_inst_dmem_n3587, MEM_stage_inst_dmem_n3586, MEM_stage_inst_dmem_n3585, MEM_stage_inst_dmem_n3584, MEM_stage_inst_dmem_n3583, MEM_stage_inst_dmem_n3582, MEM_stage_inst_dmem_n3581, MEM_stage_inst_dmem_n3580, MEM_stage_inst_dmem_n3579, MEM_stage_inst_dmem_n3578, MEM_stage_inst_dmem_n3577, MEM_stage_inst_dmem_n3576, MEM_stage_inst_dmem_n3575, MEM_stage_inst_dmem_n3574, MEM_stage_inst_dmem_n3573, MEM_stage_inst_dmem_n3572, MEM_stage_inst_dmem_n3571, MEM_stage_inst_dmem_n3570, MEM_stage_inst_dmem_n3569, MEM_stage_inst_dmem_n3568, MEM_stage_inst_dmem_n3567, MEM_stage_inst_dmem_n3566, MEM_stage_inst_dmem_n3565, MEM_stage_inst_dmem_n3564, MEM_stage_inst_dmem_n3563, MEM_stage_inst_dmem_n3562, MEM_stage_inst_dmem_n3561, MEM_stage_inst_dmem_n3560, MEM_stage_inst_dmem_n3559, MEM_stage_inst_dmem_n3558, MEM_stage_inst_dmem_n3557, MEM_stage_inst_dmem_n3556, MEM_stage_inst_dmem_n3555, MEM_stage_inst_dmem_n3554, MEM_stage_inst_dmem_n3553, MEM_stage_inst_dmem_n3552, MEM_stage_inst_dmem_n3551, MEM_stage_inst_dmem_n3550, MEM_stage_inst_dmem_n3549, MEM_stage_inst_dmem_n3548, MEM_stage_inst_dmem_n3547, MEM_stage_inst_dmem_n3546, MEM_stage_inst_dmem_n3545, MEM_stage_inst_dmem_n3544, MEM_stage_inst_dmem_n3543, MEM_stage_inst_dmem_n3542, MEM_stage_inst_dmem_n3541, MEM_stage_inst_dmem_n3540, MEM_stage_inst_dmem_n3539, MEM_stage_inst_dmem_n3538, MEM_stage_inst_dmem_n3537, MEM_stage_inst_dmem_n3536, MEM_stage_inst_dmem_n3535, MEM_stage_inst_dmem_n3534, MEM_stage_inst_dmem_n3533, MEM_stage_inst_dmem_n3532, MEM_stage_inst_dmem_n3531, MEM_stage_inst_dmem_n3530, MEM_stage_inst_dmem_n3529, MEM_stage_inst_dmem_n3528, MEM_stage_inst_dmem_n3527, MEM_stage_inst_dmem_n3526, MEM_stage_inst_dmem_n3525, MEM_stage_inst_dmem_n3524, MEM_stage_inst_dmem_n3523, MEM_stage_inst_dmem_n3522, MEM_stage_inst_dmem_n3521, MEM_stage_inst_dmem_n3520, MEM_stage_inst_dmem_n3519, MEM_stage_inst_dmem_n3518, MEM_stage_inst_dmem_n3517, MEM_stage_inst_dmem_n3516, MEM_stage_inst_dmem_n3515, MEM_stage_inst_dmem_n3514, MEM_stage_inst_dmem_n3513, MEM_stage_inst_dmem_n3512, MEM_stage_inst_dmem_n3511, MEM_stage_inst_dmem_n3510, MEM_stage_inst_dmem_n3509, MEM_stage_inst_dmem_n3508, MEM_stage_inst_dmem_n3507, MEM_stage_inst_dmem_n3506, MEM_stage_inst_dmem_n3505, MEM_stage_inst_dmem_n3504, MEM_stage_inst_dmem_n3503, MEM_stage_inst_dmem_n3502, MEM_stage_inst_dmem_n3501, MEM_stage_inst_dmem_n3500, MEM_stage_inst_dmem_n3499, MEM_stage_inst_dmem_n3498, MEM_stage_inst_dmem_n3497, MEM_stage_inst_dmem_n3496, MEM_stage_inst_dmem_n3495, MEM_stage_inst_dmem_n3494, MEM_stage_inst_dmem_n3493, MEM_stage_inst_dmem_n3492, MEM_stage_inst_dmem_n3491, MEM_stage_inst_dmem_n3490, MEM_stage_inst_dmem_n3489, MEM_stage_inst_dmem_n3488, MEM_stage_inst_dmem_n3487, MEM_stage_inst_dmem_n3486, MEM_stage_inst_dmem_n3485, MEM_stage_inst_dmem_n3484, MEM_stage_inst_dmem_n3483, MEM_stage_inst_dmem_n3482, MEM_stage_inst_dmem_n3481, MEM_stage_inst_dmem_n3480, MEM_stage_inst_dmem_n3479, MEM_stage_inst_dmem_n3478, MEM_stage_inst_dmem_n3477, MEM_stage_inst_dmem_n3476, MEM_stage_inst_dmem_n3475, MEM_stage_inst_dmem_n3474, MEM_stage_inst_dmem_n3473, MEM_stage_inst_dmem_n3472, MEM_stage_inst_dmem_n3471, MEM_stage_inst_dmem_n3470, MEM_stage_inst_dmem_n3469, MEM_stage_inst_dmem_n3468, MEM_stage_inst_dmem_n3467, MEM_stage_inst_dmem_n3466, MEM_stage_inst_dmem_n3465, MEM_stage_inst_dmem_n3464, MEM_stage_inst_dmem_n3463, MEM_stage_inst_dmem_n3462, MEM_stage_inst_dmem_n3461, MEM_stage_inst_dmem_n3460, MEM_stage_inst_dmem_n3459, MEM_stage_inst_dmem_n3458, MEM_stage_inst_dmem_n3457, MEM_stage_inst_dmem_n3456, MEM_stage_inst_dmem_n3455, MEM_stage_inst_dmem_n3454, MEM_stage_inst_dmem_n3453, MEM_stage_inst_dmem_n3452, MEM_stage_inst_dmem_n3451, MEM_stage_inst_dmem_n3450, MEM_stage_inst_dmem_n3449, MEM_stage_inst_dmem_n3448, MEM_stage_inst_dmem_n3447, MEM_stage_inst_dmem_n3446, MEM_stage_inst_dmem_n3445, MEM_stage_inst_dmem_n3444, MEM_stage_inst_dmem_n3443, MEM_stage_inst_dmem_n3442, MEM_stage_inst_dmem_n3441, MEM_stage_inst_dmem_n3440, MEM_stage_inst_dmem_n3439, MEM_stage_inst_dmem_n3438, MEM_stage_inst_dmem_n3437, MEM_stage_inst_dmem_n3436, MEM_stage_inst_dmem_n3435, MEM_stage_inst_dmem_n3434, MEM_stage_inst_dmem_n3433, MEM_stage_inst_dmem_n3432, MEM_stage_inst_dmem_n3431, MEM_stage_inst_dmem_n3430, MEM_stage_inst_dmem_n3429, MEM_stage_inst_dmem_n3428, MEM_stage_inst_dmem_n3427, MEM_stage_inst_dmem_n3426, MEM_stage_inst_dmem_n3425, MEM_stage_inst_dmem_n3424, MEM_stage_inst_dmem_n3423, MEM_stage_inst_dmem_n3422, MEM_stage_inst_dmem_n3421, MEM_stage_inst_dmem_n3420, MEM_stage_inst_dmem_n3419, MEM_stage_inst_dmem_n3418, MEM_stage_inst_dmem_n3417, MEM_stage_inst_dmem_n3416, MEM_stage_inst_dmem_n3415, MEM_stage_inst_dmem_n3414, MEM_stage_inst_dmem_n3413, MEM_stage_inst_dmem_n3412, MEM_stage_inst_dmem_n3411, MEM_stage_inst_dmem_n3410, MEM_stage_inst_dmem_n3409, MEM_stage_inst_dmem_n3408, MEM_stage_inst_dmem_n3407, MEM_stage_inst_dmem_n3406, MEM_stage_inst_dmem_n3405, MEM_stage_inst_dmem_n3404, MEM_stage_inst_dmem_n3403, MEM_stage_inst_dmem_n3402, MEM_stage_inst_dmem_n3401, MEM_stage_inst_dmem_n3400, MEM_stage_inst_dmem_n3399, MEM_stage_inst_dmem_n3398, MEM_stage_inst_dmem_n3397, MEM_stage_inst_dmem_n3396, MEM_stage_inst_dmem_n3395, MEM_stage_inst_dmem_n3394, MEM_stage_inst_dmem_n3393, MEM_stage_inst_dmem_n3392, MEM_stage_inst_dmem_n3391, MEM_stage_inst_dmem_n3390, MEM_stage_inst_dmem_n3389, MEM_stage_inst_dmem_n3388, MEM_stage_inst_dmem_n3387, MEM_stage_inst_dmem_n3386, MEM_stage_inst_dmem_n3385, MEM_stage_inst_dmem_n3384, MEM_stage_inst_dmem_n3383, MEM_stage_inst_dmem_n3382, MEM_stage_inst_dmem_n3381, MEM_stage_inst_dmem_n3380, MEM_stage_inst_dmem_n3379, MEM_stage_inst_dmem_n3378, MEM_stage_inst_dmem_n3377, MEM_stage_inst_dmem_n3376, MEM_stage_inst_dmem_n3375, MEM_stage_inst_dmem_n3374, MEM_stage_inst_dmem_n3373, MEM_stage_inst_dmem_n3372, MEM_stage_inst_dmem_n3371, MEM_stage_inst_dmem_n3370, MEM_stage_inst_dmem_n3369, MEM_stage_inst_dmem_n3368, MEM_stage_inst_dmem_n3367, MEM_stage_inst_dmem_n3366, MEM_stage_inst_dmem_n3365, MEM_stage_inst_dmem_n3364, MEM_stage_inst_dmem_n3363, MEM_stage_inst_dmem_n3362, MEM_stage_inst_dmem_n3361, MEM_stage_inst_dmem_n3360, MEM_stage_inst_dmem_n3359, MEM_stage_inst_dmem_n3358, MEM_stage_inst_dmem_n3357, MEM_stage_inst_dmem_n3356, MEM_stage_inst_dmem_n3355, MEM_stage_inst_dmem_n3354, MEM_stage_inst_dmem_n3353, MEM_stage_inst_dmem_n3352, MEM_stage_inst_dmem_n3351, MEM_stage_inst_dmem_n3350, MEM_stage_inst_dmem_n3349, MEM_stage_inst_dmem_n3348, MEM_stage_inst_dmem_n3347, MEM_stage_inst_dmem_n3346, MEM_stage_inst_dmem_n3345, MEM_stage_inst_dmem_n3344, MEM_stage_inst_dmem_n3343, MEM_stage_inst_dmem_n3342, MEM_stage_inst_dmem_n3341, MEM_stage_inst_dmem_n3340, MEM_stage_inst_dmem_n3339, MEM_stage_inst_dmem_n3338, MEM_stage_inst_dmem_n3337, MEM_stage_inst_dmem_n3336, MEM_stage_inst_dmem_n3335, MEM_stage_inst_dmem_n3334, MEM_stage_inst_dmem_n3333, MEM_stage_inst_dmem_n3332, MEM_stage_inst_dmem_n3331, MEM_stage_inst_dmem_n3330, MEM_stage_inst_dmem_n3329, MEM_stage_inst_dmem_n3328, MEM_stage_inst_dmem_n3327, MEM_stage_inst_dmem_n3326, MEM_stage_inst_dmem_n3325, MEM_stage_inst_dmem_n3324, MEM_stage_inst_dmem_n3323, MEM_stage_inst_dmem_n3322, MEM_stage_inst_dmem_n3321, MEM_stage_inst_dmem_n3320, MEM_stage_inst_dmem_n3319, MEM_stage_inst_dmem_n3318, MEM_stage_inst_dmem_n3317, MEM_stage_inst_dmem_n3316, MEM_stage_inst_dmem_n3315, MEM_stage_inst_dmem_n3314, MEM_stage_inst_dmem_n3313, MEM_stage_inst_dmem_n3312, MEM_stage_inst_dmem_n3311, MEM_stage_inst_dmem_n3310, MEM_stage_inst_dmem_n3309, MEM_stage_inst_dmem_n3308, MEM_stage_inst_dmem_n3307, MEM_stage_inst_dmem_n3306, MEM_stage_inst_dmem_n3305, MEM_stage_inst_dmem_n3304, MEM_stage_inst_dmem_n3303, MEM_stage_inst_dmem_n3302, MEM_stage_inst_dmem_n3301, MEM_stage_inst_dmem_n3300, MEM_stage_inst_dmem_n3299, MEM_stage_inst_dmem_n3298, MEM_stage_inst_dmem_n3297, MEM_stage_inst_dmem_n3296, MEM_stage_inst_dmem_n3295, MEM_stage_inst_dmem_n3294, MEM_stage_inst_dmem_n3293, MEM_stage_inst_dmem_n3292, MEM_stage_inst_dmem_n3291, MEM_stage_inst_dmem_n3290, MEM_stage_inst_dmem_n3289, MEM_stage_inst_dmem_n3288, MEM_stage_inst_dmem_n3287, MEM_stage_inst_dmem_n3286, MEM_stage_inst_dmem_n3285, MEM_stage_inst_dmem_n3284, MEM_stage_inst_dmem_n3283, MEM_stage_inst_dmem_n3282, MEM_stage_inst_dmem_n3281, MEM_stage_inst_dmem_n3280, MEM_stage_inst_dmem_n3279, MEM_stage_inst_dmem_n3278, MEM_stage_inst_dmem_n3277, MEM_stage_inst_dmem_n3276, MEM_stage_inst_dmem_n3275, MEM_stage_inst_dmem_n3274, MEM_stage_inst_dmem_n3273, MEM_stage_inst_dmem_n3272, MEM_stage_inst_dmem_n3271, MEM_stage_inst_dmem_n3270, MEM_stage_inst_dmem_n3269, MEM_stage_inst_dmem_n3268, MEM_stage_inst_dmem_n3267, MEM_stage_inst_dmem_n3266, MEM_stage_inst_dmem_n3265, MEM_stage_inst_dmem_n3264, MEM_stage_inst_dmem_n3263, MEM_stage_inst_dmem_n3262, MEM_stage_inst_dmem_n3261, MEM_stage_inst_dmem_n3260, MEM_stage_inst_dmem_n3259, MEM_stage_inst_dmem_n3258, MEM_stage_inst_dmem_n3257, MEM_stage_inst_dmem_n3256, MEM_stage_inst_dmem_n3255, MEM_stage_inst_dmem_n3254, MEM_stage_inst_dmem_n3253, MEM_stage_inst_dmem_n3252, MEM_stage_inst_dmem_n3251, MEM_stage_inst_dmem_n3250, MEM_stage_inst_dmem_n3249, MEM_stage_inst_dmem_n3248, MEM_stage_inst_dmem_n3247, MEM_stage_inst_dmem_n3246, MEM_stage_inst_dmem_n3245, MEM_stage_inst_dmem_n3244, MEM_stage_inst_dmem_n3243, MEM_stage_inst_dmem_n3242, MEM_stage_inst_dmem_n3241, MEM_stage_inst_dmem_n3240, MEM_stage_inst_dmem_n3239, MEM_stage_inst_dmem_n3238, MEM_stage_inst_dmem_n3237, MEM_stage_inst_dmem_n3236, MEM_stage_inst_dmem_n3235, MEM_stage_inst_dmem_n3234, MEM_stage_inst_dmem_n3233, MEM_stage_inst_dmem_n3232, MEM_stage_inst_dmem_n3231, MEM_stage_inst_dmem_n3230, MEM_stage_inst_dmem_n3229, MEM_stage_inst_dmem_n3228, MEM_stage_inst_dmem_n3227, MEM_stage_inst_dmem_n3226, MEM_stage_inst_dmem_n3225, MEM_stage_inst_dmem_n3224, MEM_stage_inst_dmem_n3223, MEM_stage_inst_dmem_n3222, MEM_stage_inst_dmem_n3221, MEM_stage_inst_dmem_n3220, MEM_stage_inst_dmem_n3219, MEM_stage_inst_dmem_n3218, MEM_stage_inst_dmem_n3217, MEM_stage_inst_dmem_n3216, MEM_stage_inst_dmem_n3215, MEM_stage_inst_dmem_n3214, MEM_stage_inst_dmem_n3213, MEM_stage_inst_dmem_n3212, MEM_stage_inst_dmem_n3211, MEM_stage_inst_dmem_n3210, MEM_stage_inst_dmem_n3209, MEM_stage_inst_dmem_n3208, MEM_stage_inst_dmem_n3207, MEM_stage_inst_dmem_n3206, MEM_stage_inst_dmem_n3205, MEM_stage_inst_dmem_n3204, MEM_stage_inst_dmem_n3203, MEM_stage_inst_dmem_n3202, MEM_stage_inst_dmem_n3201, MEM_stage_inst_dmem_n3200, MEM_stage_inst_dmem_n3199, MEM_stage_inst_dmem_n3198, MEM_stage_inst_dmem_n3197, MEM_stage_inst_dmem_n3196, MEM_stage_inst_dmem_n3195, MEM_stage_inst_dmem_n3194, MEM_stage_inst_dmem_n3193, MEM_stage_inst_dmem_n3192, MEM_stage_inst_dmem_n3191, MEM_stage_inst_dmem_n3190, MEM_stage_inst_dmem_n3189, MEM_stage_inst_dmem_n3188, MEM_stage_inst_dmem_n3187, MEM_stage_inst_dmem_n3186, MEM_stage_inst_dmem_n3185, MEM_stage_inst_dmem_n3184, MEM_stage_inst_dmem_n3183, MEM_stage_inst_dmem_n3182, MEM_stage_inst_dmem_n3181, MEM_stage_inst_dmem_n3180, MEM_stage_inst_dmem_n3179, MEM_stage_inst_dmem_n3178, MEM_stage_inst_dmem_n3177, MEM_stage_inst_dmem_n3176, MEM_stage_inst_dmem_n3175, MEM_stage_inst_dmem_n3174, MEM_stage_inst_dmem_n3173, MEM_stage_inst_dmem_n3172, MEM_stage_inst_dmem_n3171, MEM_stage_inst_dmem_n3170, MEM_stage_inst_dmem_n3169, MEM_stage_inst_dmem_n3168, MEM_stage_inst_dmem_n3167, MEM_stage_inst_dmem_n3166, MEM_stage_inst_dmem_n3165, MEM_stage_inst_dmem_n3164, MEM_stage_inst_dmem_n3163, MEM_stage_inst_dmem_n3162, MEM_stage_inst_dmem_n3161, MEM_stage_inst_dmem_n3160, MEM_stage_inst_dmem_n3159, MEM_stage_inst_dmem_n3158, MEM_stage_inst_dmem_n3157, MEM_stage_inst_dmem_n3156, MEM_stage_inst_dmem_n3155, MEM_stage_inst_dmem_n3154, MEM_stage_inst_dmem_n3153, MEM_stage_inst_dmem_n3152, MEM_stage_inst_dmem_n3151, MEM_stage_inst_dmem_n3150, MEM_stage_inst_dmem_n3149, MEM_stage_inst_dmem_n3148, MEM_stage_inst_dmem_n3147, MEM_stage_inst_dmem_n3146, MEM_stage_inst_dmem_n3145, MEM_stage_inst_dmem_n3144, MEM_stage_inst_dmem_n3143, MEM_stage_inst_dmem_n3142, MEM_stage_inst_dmem_n3141, MEM_stage_inst_dmem_n3140, MEM_stage_inst_dmem_n3139, MEM_stage_inst_dmem_n3138, MEM_stage_inst_dmem_n3137, MEM_stage_inst_dmem_n3136, MEM_stage_inst_dmem_n3135, MEM_stage_inst_dmem_n3134, MEM_stage_inst_dmem_n3133, MEM_stage_inst_dmem_n3132, MEM_stage_inst_dmem_n3131, MEM_stage_inst_dmem_n3130, MEM_stage_inst_dmem_n3129, MEM_stage_inst_dmem_n3128, MEM_stage_inst_dmem_n3127, MEM_stage_inst_dmem_n3126, MEM_stage_inst_dmem_n3125, MEM_stage_inst_dmem_n3124, MEM_stage_inst_dmem_n3123, MEM_stage_inst_dmem_n3122, MEM_stage_inst_dmem_n3121, MEM_stage_inst_dmem_n3120, MEM_stage_inst_dmem_n3119, MEM_stage_inst_dmem_n3118, MEM_stage_inst_dmem_n3117, MEM_stage_inst_dmem_n3116, MEM_stage_inst_dmem_n3115, MEM_stage_inst_dmem_n3114, MEM_stage_inst_dmem_n3113, MEM_stage_inst_dmem_n3112, MEM_stage_inst_dmem_n3111, MEM_stage_inst_dmem_n3110, MEM_stage_inst_dmem_n3109, MEM_stage_inst_dmem_n3108, MEM_stage_inst_dmem_n3107, MEM_stage_inst_dmem_n3106, MEM_stage_inst_dmem_n3105, MEM_stage_inst_dmem_n3104, MEM_stage_inst_dmem_n3103, MEM_stage_inst_dmem_n3102, MEM_stage_inst_dmem_n3101, MEM_stage_inst_dmem_n3100, MEM_stage_inst_dmem_n3099, MEM_stage_inst_dmem_n3098, MEM_stage_inst_dmem_n3097, MEM_stage_inst_dmem_n3096, MEM_stage_inst_dmem_n3095, MEM_stage_inst_dmem_n3094, MEM_stage_inst_dmem_n3093, MEM_stage_inst_dmem_n3092, MEM_stage_inst_dmem_n3091, MEM_stage_inst_dmem_n3090, MEM_stage_inst_dmem_n3089, MEM_stage_inst_dmem_n3088, MEM_stage_inst_dmem_n3087, MEM_stage_inst_dmem_n3086, MEM_stage_inst_dmem_n3085, MEM_stage_inst_dmem_n3084, MEM_stage_inst_dmem_n3083, MEM_stage_inst_dmem_n3082, MEM_stage_inst_dmem_n3081, MEM_stage_inst_dmem_n3080, MEM_stage_inst_dmem_n3079, MEM_stage_inst_dmem_n3078, MEM_stage_inst_dmem_n3077, MEM_stage_inst_dmem_n3076, MEM_stage_inst_dmem_n3075, MEM_stage_inst_dmem_n3074, MEM_stage_inst_dmem_n3073, MEM_stage_inst_dmem_n3072, MEM_stage_inst_dmem_n3071, MEM_stage_inst_dmem_n3070, MEM_stage_inst_dmem_n3069, MEM_stage_inst_dmem_n3068, MEM_stage_inst_dmem_n3067, MEM_stage_inst_dmem_n3066, MEM_stage_inst_dmem_n3065, MEM_stage_inst_dmem_n3064, MEM_stage_inst_dmem_n3063, MEM_stage_inst_dmem_n3062, MEM_stage_inst_dmem_n3061, MEM_stage_inst_dmem_n3060, MEM_stage_inst_dmem_n3059, MEM_stage_inst_dmem_n3058, MEM_stage_inst_dmem_n3057, MEM_stage_inst_dmem_n3056, MEM_stage_inst_dmem_n3055, MEM_stage_inst_dmem_n3054, MEM_stage_inst_dmem_n3053, MEM_stage_inst_dmem_n3052, MEM_stage_inst_dmem_n3051, MEM_stage_inst_dmem_n3050, MEM_stage_inst_dmem_n3049, MEM_stage_inst_dmem_n3048, MEM_stage_inst_dmem_n3047, MEM_stage_inst_dmem_n3046, MEM_stage_inst_dmem_n3045, MEM_stage_inst_dmem_n3044, MEM_stage_inst_dmem_n3043, MEM_stage_inst_dmem_n3042, MEM_stage_inst_dmem_n3041, MEM_stage_inst_dmem_n3040, MEM_stage_inst_dmem_n3039, MEM_stage_inst_dmem_n3038, MEM_stage_inst_dmem_n3037, MEM_stage_inst_dmem_n3036, MEM_stage_inst_dmem_n3035, MEM_stage_inst_dmem_n3034, MEM_stage_inst_dmem_n3033, MEM_stage_inst_dmem_n3032, MEM_stage_inst_dmem_n3031, MEM_stage_inst_dmem_n3030, MEM_stage_inst_dmem_n3029, MEM_stage_inst_dmem_n3028, MEM_stage_inst_dmem_n3027, MEM_stage_inst_dmem_n3026, MEM_stage_inst_dmem_n3025, MEM_stage_inst_dmem_n3024, MEM_stage_inst_dmem_n3023, MEM_stage_inst_dmem_n3022, MEM_stage_inst_dmem_n3021, MEM_stage_inst_dmem_n3020, MEM_stage_inst_dmem_n3019, MEM_stage_inst_dmem_n3018, MEM_stage_inst_dmem_n3017, MEM_stage_inst_dmem_n3016, MEM_stage_inst_dmem_n3015, MEM_stage_inst_dmem_n3014, MEM_stage_inst_dmem_n3013, MEM_stage_inst_dmem_n3012, MEM_stage_inst_dmem_n3011, MEM_stage_inst_dmem_n3010, MEM_stage_inst_dmem_n3009, MEM_stage_inst_dmem_n3008, MEM_stage_inst_dmem_n3007, MEM_stage_inst_dmem_n3006, MEM_stage_inst_dmem_n3005, MEM_stage_inst_dmem_n3004, MEM_stage_inst_dmem_n3003, MEM_stage_inst_dmem_n3002, MEM_stage_inst_dmem_n3001, MEM_stage_inst_dmem_n3000, MEM_stage_inst_dmem_n2999, MEM_stage_inst_dmem_n2998, MEM_stage_inst_dmem_n2997, MEM_stage_inst_dmem_n2996, MEM_stage_inst_dmem_n2995, MEM_stage_inst_dmem_n2994, MEM_stage_inst_dmem_n2993, MEM_stage_inst_dmem_n2992, MEM_stage_inst_dmem_n2991, MEM_stage_inst_dmem_n2990, MEM_stage_inst_dmem_n2989, MEM_stage_inst_dmem_n2988, MEM_stage_inst_dmem_n2987, MEM_stage_inst_dmem_n2986, MEM_stage_inst_dmem_n2985, MEM_stage_inst_dmem_n2984, MEM_stage_inst_dmem_n2983, MEM_stage_inst_dmem_n2982, MEM_stage_inst_dmem_n2981, MEM_stage_inst_dmem_n2980, MEM_stage_inst_dmem_n2979, MEM_stage_inst_dmem_n2978, MEM_stage_inst_dmem_n2977, MEM_stage_inst_dmem_n2976, MEM_stage_inst_dmem_n2975, MEM_stage_inst_dmem_n2974, MEM_stage_inst_dmem_n2973, MEM_stage_inst_dmem_n2972, MEM_stage_inst_dmem_n2971, MEM_stage_inst_dmem_n2970, MEM_stage_inst_dmem_n2969, MEM_stage_inst_dmem_n2968, MEM_stage_inst_dmem_n2967, MEM_stage_inst_dmem_n2966, MEM_stage_inst_dmem_n2965, MEM_stage_inst_dmem_n2964, MEM_stage_inst_dmem_n2963, MEM_stage_inst_dmem_n2962, MEM_stage_inst_dmem_n2961, MEM_stage_inst_dmem_n2960, MEM_stage_inst_dmem_n2959, MEM_stage_inst_dmem_n2958, MEM_stage_inst_dmem_n2957, MEM_stage_inst_dmem_n2956, MEM_stage_inst_dmem_n2955, MEM_stage_inst_dmem_n2954, MEM_stage_inst_dmem_n2953, MEM_stage_inst_dmem_n2952, MEM_stage_inst_dmem_n2951, MEM_stage_inst_dmem_n2950, MEM_stage_inst_dmem_n2949, MEM_stage_inst_dmem_n2948, MEM_stage_inst_dmem_n2947, MEM_stage_inst_dmem_n2946, MEM_stage_inst_dmem_n2945, MEM_stage_inst_dmem_n2944, MEM_stage_inst_dmem_n2943, MEM_stage_inst_dmem_n2942, MEM_stage_inst_dmem_n2941, MEM_stage_inst_dmem_n2940, MEM_stage_inst_dmem_n2939, MEM_stage_inst_dmem_n2938, MEM_stage_inst_dmem_n2937, MEM_stage_inst_dmem_n2936, MEM_stage_inst_dmem_n2935, MEM_stage_inst_dmem_n2934, MEM_stage_inst_dmem_n2933, MEM_stage_inst_dmem_n2932, MEM_stage_inst_dmem_n2931, MEM_stage_inst_dmem_n2930, MEM_stage_inst_dmem_n2929, MEM_stage_inst_dmem_n2928, MEM_stage_inst_dmem_n2927, MEM_stage_inst_dmem_n2926, MEM_stage_inst_dmem_n2925, MEM_stage_inst_dmem_n2924, MEM_stage_inst_dmem_n2923, MEM_stage_inst_dmem_n2922, MEM_stage_inst_dmem_n2921, MEM_stage_inst_dmem_n2920, MEM_stage_inst_dmem_n2919, MEM_stage_inst_dmem_n2918, MEM_stage_inst_dmem_n2917, MEM_stage_inst_dmem_n2916, MEM_stage_inst_dmem_n2915, MEM_stage_inst_dmem_n2914, MEM_stage_inst_dmem_n2913, MEM_stage_inst_dmem_n2912, MEM_stage_inst_dmem_n2911, MEM_stage_inst_dmem_n2910, MEM_stage_inst_dmem_n2909, MEM_stage_inst_dmem_n2908, MEM_stage_inst_dmem_n2907, MEM_stage_inst_dmem_n2906, MEM_stage_inst_dmem_n2905, MEM_stage_inst_dmem_n2904, MEM_stage_inst_dmem_n2903, MEM_stage_inst_dmem_n2902, MEM_stage_inst_dmem_n2901, MEM_stage_inst_dmem_n2900, MEM_stage_inst_dmem_n2899, MEM_stage_inst_dmem_n2898, MEM_stage_inst_dmem_n2897, MEM_stage_inst_dmem_n2896, MEM_stage_inst_dmem_n2895, MEM_stage_inst_dmem_n2894, MEM_stage_inst_dmem_n2893, MEM_stage_inst_dmem_n2892, MEM_stage_inst_dmem_n2891, MEM_stage_inst_dmem_n2890, MEM_stage_inst_dmem_n2889, MEM_stage_inst_dmem_n2888, MEM_stage_inst_dmem_n2887, MEM_stage_inst_dmem_n2886, MEM_stage_inst_dmem_n2885, MEM_stage_inst_dmem_n2884, MEM_stage_inst_dmem_n2883, MEM_stage_inst_dmem_n2882, MEM_stage_inst_dmem_n2881, MEM_stage_inst_dmem_n2880, MEM_stage_inst_dmem_n2879, MEM_stage_inst_dmem_n2878, MEM_stage_inst_dmem_n2877, MEM_stage_inst_dmem_n2876, MEM_stage_inst_dmem_n2875, MEM_stage_inst_dmem_n2874, MEM_stage_inst_dmem_n2873, MEM_stage_inst_dmem_n2872, MEM_stage_inst_dmem_n2871, MEM_stage_inst_dmem_n2870, MEM_stage_inst_dmem_n2869, MEM_stage_inst_dmem_n2868, MEM_stage_inst_dmem_n2867, MEM_stage_inst_dmem_n2866, MEM_stage_inst_dmem_n2865, MEM_stage_inst_dmem_n2864, MEM_stage_inst_dmem_n2863, MEM_stage_inst_dmem_n2862, MEM_stage_inst_dmem_n2861, MEM_stage_inst_dmem_n2860, MEM_stage_inst_dmem_n2859, MEM_stage_inst_dmem_n2858, MEM_stage_inst_dmem_n2857, MEM_stage_inst_dmem_n2856, MEM_stage_inst_dmem_n2855, MEM_stage_inst_dmem_n2854, MEM_stage_inst_dmem_n2853, MEM_stage_inst_dmem_n2852, MEM_stage_inst_dmem_n2851, MEM_stage_inst_dmem_n2850, MEM_stage_inst_dmem_n2849, MEM_stage_inst_dmem_n2848, MEM_stage_inst_dmem_n2847, MEM_stage_inst_dmem_n2846, MEM_stage_inst_dmem_n2845, MEM_stage_inst_dmem_n2844, MEM_stage_inst_dmem_n2843, MEM_stage_inst_dmem_n2842, MEM_stage_inst_dmem_n2841, MEM_stage_inst_dmem_n2840, MEM_stage_inst_dmem_n2839, MEM_stage_inst_dmem_n2838, MEM_stage_inst_dmem_n2837, MEM_stage_inst_dmem_n2836, MEM_stage_inst_dmem_n2835, MEM_stage_inst_dmem_n2834, MEM_stage_inst_dmem_n2833, MEM_stage_inst_dmem_n2832, MEM_stage_inst_dmem_n2831, MEM_stage_inst_dmem_n2830, MEM_stage_inst_dmem_n2829, MEM_stage_inst_dmem_n2828, MEM_stage_inst_dmem_n2827, MEM_stage_inst_dmem_n2826, MEM_stage_inst_dmem_n2825, MEM_stage_inst_dmem_n2824, MEM_stage_inst_dmem_n2823, MEM_stage_inst_dmem_n2822, MEM_stage_inst_dmem_n2821, MEM_stage_inst_dmem_n2820, MEM_stage_inst_dmem_n2819, MEM_stage_inst_dmem_n2818, MEM_stage_inst_dmem_n2817, MEM_stage_inst_dmem_n2816, MEM_stage_inst_dmem_n2815, MEM_stage_inst_dmem_n2814, MEM_stage_inst_dmem_n2813, MEM_stage_inst_dmem_n2812, MEM_stage_inst_dmem_n2811, MEM_stage_inst_dmem_n2810, MEM_stage_inst_dmem_n2809, MEM_stage_inst_dmem_n2808, MEM_stage_inst_dmem_n2807, MEM_stage_inst_dmem_n2806, MEM_stage_inst_dmem_n2805, MEM_stage_inst_dmem_n2804, MEM_stage_inst_dmem_n2803, MEM_stage_inst_dmem_n2802, MEM_stage_inst_dmem_n2801, MEM_stage_inst_dmem_n2800, MEM_stage_inst_dmem_n2799, MEM_stage_inst_dmem_n2798, MEM_stage_inst_dmem_n2797, MEM_stage_inst_dmem_n2796, MEM_stage_inst_dmem_n2795, MEM_stage_inst_dmem_n2794, MEM_stage_inst_dmem_n2793, MEM_stage_inst_dmem_n2792, MEM_stage_inst_dmem_n2791, MEM_stage_inst_dmem_n2790, MEM_stage_inst_dmem_n2789, MEM_stage_inst_dmem_n2788, MEM_stage_inst_dmem_n2787, MEM_stage_inst_dmem_n2786, MEM_stage_inst_dmem_n2785, MEM_stage_inst_dmem_n2784, MEM_stage_inst_dmem_n2783, MEM_stage_inst_dmem_n2782, MEM_stage_inst_dmem_n2781, MEM_stage_inst_dmem_n2780, MEM_stage_inst_dmem_n2779, MEM_stage_inst_dmem_n2778, MEM_stage_inst_dmem_n2777, MEM_stage_inst_dmem_n2776, MEM_stage_inst_dmem_n2775, MEM_stage_inst_dmem_n2774, MEM_stage_inst_dmem_n2773, MEM_stage_inst_dmem_n2772, MEM_stage_inst_dmem_n2771, MEM_stage_inst_dmem_n2770, MEM_stage_inst_dmem_n2769, MEM_stage_inst_dmem_n2768, MEM_stage_inst_dmem_n2767, MEM_stage_inst_dmem_n2766, MEM_stage_inst_dmem_n2765, MEM_stage_inst_dmem_n2764, MEM_stage_inst_dmem_n2763, MEM_stage_inst_dmem_n2762, MEM_stage_inst_dmem_n2761, MEM_stage_inst_dmem_n2760, MEM_stage_inst_dmem_n2759, MEM_stage_inst_dmem_n2758, MEM_stage_inst_dmem_n2757, MEM_stage_inst_dmem_n2756, MEM_stage_inst_dmem_n2755, MEM_stage_inst_dmem_n2754, MEM_stage_inst_dmem_n2753, MEM_stage_inst_dmem_n2752, MEM_stage_inst_dmem_n2751, MEM_stage_inst_dmem_n2750, MEM_stage_inst_dmem_n2749, MEM_stage_inst_dmem_n2748, MEM_stage_inst_dmem_n2747, MEM_stage_inst_dmem_n2746, MEM_stage_inst_dmem_n2745, MEM_stage_inst_dmem_n2744, MEM_stage_inst_dmem_n2743, MEM_stage_inst_dmem_n2742, MEM_stage_inst_dmem_n2741, MEM_stage_inst_dmem_n2740, MEM_stage_inst_dmem_n2739, MEM_stage_inst_dmem_n2738, MEM_stage_inst_dmem_n2737, MEM_stage_inst_dmem_n2736, MEM_stage_inst_dmem_n2735, MEM_stage_inst_dmem_n2734, MEM_stage_inst_dmem_n2733, MEM_stage_inst_dmem_n2732, MEM_stage_inst_dmem_n2731, MEM_stage_inst_dmem_n2730, MEM_stage_inst_dmem_n2729, MEM_stage_inst_dmem_n2728, MEM_stage_inst_dmem_n2727, MEM_stage_inst_dmem_n2726, MEM_stage_inst_dmem_n2725, MEM_stage_inst_dmem_n2724, MEM_stage_inst_dmem_n2723, MEM_stage_inst_dmem_n2722, MEM_stage_inst_dmem_n2721, MEM_stage_inst_dmem_n2720, MEM_stage_inst_dmem_n2719, MEM_stage_inst_dmem_n2718, MEM_stage_inst_dmem_n2717, MEM_stage_inst_dmem_n2716, MEM_stage_inst_dmem_n2715, MEM_stage_inst_dmem_n2714, MEM_stage_inst_dmem_n2713, MEM_stage_inst_dmem_n2712, MEM_stage_inst_dmem_n2711, MEM_stage_inst_dmem_n2710, MEM_stage_inst_dmem_n2709, MEM_stage_inst_dmem_n2708, MEM_stage_inst_dmem_n2707, MEM_stage_inst_dmem_n2706, MEM_stage_inst_dmem_n2705, MEM_stage_inst_dmem_n2704, MEM_stage_inst_dmem_n2703, MEM_stage_inst_dmem_n2702, MEM_stage_inst_dmem_n2701, MEM_stage_inst_dmem_n2700, MEM_stage_inst_dmem_n2699, MEM_stage_inst_dmem_n2698, MEM_stage_inst_dmem_n2697, MEM_stage_inst_dmem_n2696, MEM_stage_inst_dmem_n2695, MEM_stage_inst_dmem_n2694, MEM_stage_inst_dmem_n2693, MEM_stage_inst_dmem_n2692, MEM_stage_inst_dmem_n2691, MEM_stage_inst_dmem_n2690, MEM_stage_inst_dmem_n2689, MEM_stage_inst_dmem_n2688, MEM_stage_inst_dmem_n2687, MEM_stage_inst_dmem_n2686, MEM_stage_inst_dmem_n2685, MEM_stage_inst_dmem_n2684, MEM_stage_inst_dmem_n2683, MEM_stage_inst_dmem_n2682, MEM_stage_inst_dmem_n2681, MEM_stage_inst_dmem_n2680, MEM_stage_inst_dmem_n2679, MEM_stage_inst_dmem_n2678, MEM_stage_inst_dmem_n2677, MEM_stage_inst_dmem_n2676, MEM_stage_inst_dmem_n2675, MEM_stage_inst_dmem_n2674, MEM_stage_inst_dmem_n2673, MEM_stage_inst_dmem_n2672, MEM_stage_inst_dmem_n2671, MEM_stage_inst_dmem_n2670, MEM_stage_inst_dmem_n2669, MEM_stage_inst_dmem_n2668, MEM_stage_inst_dmem_n2667, MEM_stage_inst_dmem_n2666, MEM_stage_inst_dmem_n2665, MEM_stage_inst_dmem_n2664, MEM_stage_inst_dmem_n2663, MEM_stage_inst_dmem_n2662, MEM_stage_inst_dmem_n2661, MEM_stage_inst_dmem_n2660, MEM_stage_inst_dmem_n2659, MEM_stage_inst_dmem_n2658, MEM_stage_inst_dmem_n2657, MEM_stage_inst_dmem_n2656, MEM_stage_inst_dmem_n2655, MEM_stage_inst_dmem_n2654, MEM_stage_inst_dmem_n2653, MEM_stage_inst_dmem_n2652, MEM_stage_inst_dmem_n2651, MEM_stage_inst_dmem_n2650, MEM_stage_inst_dmem_n2649, MEM_stage_inst_dmem_n2648, MEM_stage_inst_dmem_n2647, MEM_stage_inst_dmem_n2646, MEM_stage_inst_dmem_n2645, MEM_stage_inst_dmem_n2644, MEM_stage_inst_dmem_n2643, MEM_stage_inst_dmem_n2642, MEM_stage_inst_dmem_n2641, MEM_stage_inst_dmem_n2640, MEM_stage_inst_dmem_n2639, MEM_stage_inst_dmem_n2638, MEM_stage_inst_dmem_n2637, MEM_stage_inst_dmem_n2636, MEM_stage_inst_dmem_n2635, MEM_stage_inst_dmem_n2634, MEM_stage_inst_dmem_n2633, MEM_stage_inst_dmem_n2632, MEM_stage_inst_dmem_n2631, MEM_stage_inst_dmem_n2630, MEM_stage_inst_dmem_n2629, MEM_stage_inst_dmem_n2628, MEM_stage_inst_dmem_n2627, MEM_stage_inst_dmem_n2626, MEM_stage_inst_dmem_n2625, MEM_stage_inst_dmem_n2624, MEM_stage_inst_dmem_n2623, MEM_stage_inst_dmem_n2622, MEM_stage_inst_dmem_n2621, MEM_stage_inst_dmem_n2620, MEM_stage_inst_dmem_n2619, MEM_stage_inst_dmem_n2618, MEM_stage_inst_dmem_n2617, MEM_stage_inst_dmem_n2616, MEM_stage_inst_dmem_n2615, MEM_stage_inst_dmem_n2614, MEM_stage_inst_dmem_n2613, MEM_stage_inst_dmem_n2612, MEM_stage_inst_dmem_n2611, MEM_stage_inst_dmem_n2610, MEM_stage_inst_dmem_n2609, MEM_stage_inst_dmem_n2608, MEM_stage_inst_dmem_n2607, MEM_stage_inst_dmem_n2606, MEM_stage_inst_dmem_n2605, MEM_stage_inst_dmem_n2604, MEM_stage_inst_dmem_n2603, MEM_stage_inst_dmem_n2602, MEM_stage_inst_dmem_n2601, MEM_stage_inst_dmem_n2600, MEM_stage_inst_dmem_n2599, MEM_stage_inst_dmem_n2598, MEM_stage_inst_dmem_n2597, MEM_stage_inst_dmem_n2596, MEM_stage_inst_dmem_n2595, MEM_stage_inst_dmem_n2594, MEM_stage_inst_dmem_n2593, MEM_stage_inst_dmem_n2592, MEM_stage_inst_dmem_n2591, MEM_stage_inst_dmem_n2590, MEM_stage_inst_dmem_n2589, MEM_stage_inst_dmem_n2588, MEM_stage_inst_dmem_n2587, MEM_stage_inst_dmem_n2586, MEM_stage_inst_dmem_n2585, MEM_stage_inst_dmem_n2584, MEM_stage_inst_dmem_n2583, MEM_stage_inst_dmem_n2582, MEM_stage_inst_dmem_n2581, MEM_stage_inst_dmem_n2580, MEM_stage_inst_dmem_n2579, MEM_stage_inst_dmem_n2578, MEM_stage_inst_dmem_n2577, MEM_stage_inst_dmem_n2576, MEM_stage_inst_dmem_n2575, MEM_stage_inst_dmem_n2574, MEM_stage_inst_dmem_n2573, MEM_stage_inst_dmem_n2572, MEM_stage_inst_dmem_n2571, MEM_stage_inst_dmem_n2570, MEM_stage_inst_dmem_n2569, MEM_stage_inst_dmem_n2568, MEM_stage_inst_dmem_n2567, MEM_stage_inst_dmem_n2566, MEM_stage_inst_dmem_n2565, MEM_stage_inst_dmem_n2564, MEM_stage_inst_dmem_n2563, MEM_stage_inst_dmem_n2562, MEM_stage_inst_dmem_n2561, MEM_stage_inst_dmem_n2560, MEM_stage_inst_dmem_n2559, MEM_stage_inst_dmem_n2558, MEM_stage_inst_dmem_n2557, MEM_stage_inst_dmem_n2556, MEM_stage_inst_dmem_n2555, MEM_stage_inst_dmem_n2554, MEM_stage_inst_dmem_n2553, MEM_stage_inst_dmem_n2552, MEM_stage_inst_dmem_n2551, MEM_stage_inst_dmem_n2550, MEM_stage_inst_dmem_n2549, MEM_stage_inst_dmem_n2548, MEM_stage_inst_dmem_n2547, MEM_stage_inst_dmem_n2546, MEM_stage_inst_dmem_n2545, MEM_stage_inst_dmem_n2544, MEM_stage_inst_dmem_n2543, MEM_stage_inst_dmem_n2542, MEM_stage_inst_dmem_n2541, MEM_stage_inst_dmem_n2540, MEM_stage_inst_dmem_n2539, MEM_stage_inst_dmem_n2538, MEM_stage_inst_dmem_n2537, MEM_stage_inst_dmem_n2536, MEM_stage_inst_dmem_n2535, MEM_stage_inst_dmem_n2534, MEM_stage_inst_dmem_n2533, MEM_stage_inst_dmem_n2532, MEM_stage_inst_dmem_n2531, MEM_stage_inst_dmem_n2530, MEM_stage_inst_dmem_n2529, MEM_stage_inst_dmem_n2528, MEM_stage_inst_dmem_n2527, MEM_stage_inst_dmem_n2526, MEM_stage_inst_dmem_n2525, MEM_stage_inst_dmem_n2524, MEM_stage_inst_dmem_n2523, MEM_stage_inst_dmem_n2522, MEM_stage_inst_dmem_n2521, MEM_stage_inst_dmem_n2520, MEM_stage_inst_dmem_n2519, MEM_stage_inst_dmem_n2518, MEM_stage_inst_dmem_n2517, MEM_stage_inst_dmem_n2516, MEM_stage_inst_dmem_n2515, MEM_stage_inst_dmem_n2514, MEM_stage_inst_dmem_n2513, MEM_stage_inst_dmem_n2512, MEM_stage_inst_dmem_n2511, MEM_stage_inst_dmem_n2510, MEM_stage_inst_dmem_n2509, MEM_stage_inst_dmem_n2508, MEM_stage_inst_dmem_n2507, MEM_stage_inst_dmem_n2506, MEM_stage_inst_dmem_n2505, MEM_stage_inst_dmem_n2504, MEM_stage_inst_dmem_n2503, MEM_stage_inst_dmem_n2502, MEM_stage_inst_dmem_n2501, MEM_stage_inst_dmem_n2500, MEM_stage_inst_dmem_n2499, MEM_stage_inst_dmem_n2498, MEM_stage_inst_dmem_n2497, MEM_stage_inst_dmem_n2496, MEM_stage_inst_dmem_n2495, MEM_stage_inst_dmem_n2494, MEM_stage_inst_dmem_n2493, MEM_stage_inst_dmem_n2492, MEM_stage_inst_dmem_n2491, MEM_stage_inst_dmem_n2490, MEM_stage_inst_dmem_n2489, MEM_stage_inst_dmem_n2488, MEM_stage_inst_dmem_n2487, MEM_stage_inst_dmem_n2486, MEM_stage_inst_dmem_n2485, MEM_stage_inst_dmem_n2484, MEM_stage_inst_dmem_n2483, MEM_stage_inst_dmem_n2482, MEM_stage_inst_dmem_n2481, MEM_stage_inst_dmem_n2480, MEM_stage_inst_dmem_n2479, MEM_stage_inst_dmem_n2478, MEM_stage_inst_dmem_n2477, MEM_stage_inst_dmem_n2476, MEM_stage_inst_dmem_n2475, MEM_stage_inst_dmem_n2474, MEM_stage_inst_dmem_n2473, MEM_stage_inst_dmem_n2472, MEM_stage_inst_dmem_n2471, MEM_stage_inst_dmem_n2470, MEM_stage_inst_dmem_n2469, MEM_stage_inst_dmem_n2468, MEM_stage_inst_dmem_n2467, MEM_stage_inst_dmem_n2466, MEM_stage_inst_dmem_n2465, MEM_stage_inst_dmem_n2464, MEM_stage_inst_dmem_n2463, MEM_stage_inst_dmem_n2462, MEM_stage_inst_dmem_n2461, MEM_stage_inst_dmem_n2460, MEM_stage_inst_dmem_n2459, MEM_stage_inst_dmem_n2458, MEM_stage_inst_dmem_n2457, MEM_stage_inst_dmem_n2456, MEM_stage_inst_dmem_n2455, MEM_stage_inst_dmem_n2454, MEM_stage_inst_dmem_n2453, MEM_stage_inst_dmem_n2452, MEM_stage_inst_dmem_n2451, MEM_stage_inst_dmem_n2450, MEM_stage_inst_dmem_n2449, MEM_stage_inst_dmem_n2448, MEM_stage_inst_dmem_n2447, MEM_stage_inst_dmem_n2446, MEM_stage_inst_dmem_n2445, MEM_stage_inst_dmem_n2444, MEM_stage_inst_dmem_n2443, MEM_stage_inst_dmem_n2442, MEM_stage_inst_dmem_n2441, MEM_stage_inst_dmem_n2440, MEM_stage_inst_dmem_n2439, MEM_stage_inst_dmem_n2438, MEM_stage_inst_dmem_n2437, MEM_stage_inst_dmem_n2436, MEM_stage_inst_dmem_n2435, MEM_stage_inst_dmem_n2434, MEM_stage_inst_dmem_n2433, MEM_stage_inst_dmem_n2432, MEM_stage_inst_dmem_n2431, MEM_stage_inst_dmem_n2430, MEM_stage_inst_dmem_n2429, MEM_stage_inst_dmem_n2428, MEM_stage_inst_dmem_n2427, MEM_stage_inst_dmem_n2426, MEM_stage_inst_dmem_n2425, MEM_stage_inst_dmem_n2424, MEM_stage_inst_dmem_n2423, MEM_stage_inst_dmem_n2422, MEM_stage_inst_dmem_n2421, MEM_stage_inst_dmem_n2420, MEM_stage_inst_dmem_n2419, MEM_stage_inst_dmem_n2418, MEM_stage_inst_dmem_n2417, MEM_stage_inst_dmem_n2416, MEM_stage_inst_dmem_n2415, MEM_stage_inst_dmem_n2414, MEM_stage_inst_dmem_n2413, MEM_stage_inst_dmem_n2412, MEM_stage_inst_dmem_n2411, MEM_stage_inst_dmem_n2410, MEM_stage_inst_dmem_n2409, MEM_stage_inst_dmem_n2408, MEM_stage_inst_dmem_n2407, MEM_stage_inst_dmem_n2406, MEM_stage_inst_dmem_n2405, MEM_stage_inst_dmem_n2404, MEM_stage_inst_dmem_n2403, MEM_stage_inst_dmem_n2402, MEM_stage_inst_dmem_n2401, MEM_stage_inst_dmem_n2400, MEM_stage_inst_dmem_n2399, MEM_stage_inst_dmem_n2398, MEM_stage_inst_dmem_n2397, MEM_stage_inst_dmem_n2396, MEM_stage_inst_dmem_n2395, MEM_stage_inst_dmem_n2394, MEM_stage_inst_dmem_n2393, MEM_stage_inst_dmem_n2392, MEM_stage_inst_dmem_n2391, MEM_stage_inst_dmem_n2390, MEM_stage_inst_dmem_n2389, MEM_stage_inst_dmem_n2388, MEM_stage_inst_dmem_n2387, MEM_stage_inst_dmem_n2386, MEM_stage_inst_dmem_n2385, MEM_stage_inst_dmem_n2384, MEM_stage_inst_dmem_n2383, MEM_stage_inst_dmem_n2382, MEM_stage_inst_dmem_n2381, MEM_stage_inst_dmem_n2380, MEM_stage_inst_dmem_n2379, MEM_stage_inst_dmem_n2378, MEM_stage_inst_dmem_n2377, MEM_stage_inst_dmem_n2376, MEM_stage_inst_dmem_n2375, MEM_stage_inst_dmem_n2374, MEM_stage_inst_dmem_n2373, MEM_stage_inst_dmem_n2372, MEM_stage_inst_dmem_n2371, MEM_stage_inst_dmem_n2370, MEM_stage_inst_dmem_n2369, MEM_stage_inst_dmem_n2368, MEM_stage_inst_dmem_n2367, MEM_stage_inst_dmem_n2366, MEM_stage_inst_dmem_n2365, MEM_stage_inst_dmem_n2364, MEM_stage_inst_dmem_n2363, MEM_stage_inst_dmem_n2362, MEM_stage_inst_dmem_n2361, MEM_stage_inst_dmem_n2360, MEM_stage_inst_dmem_n2359, MEM_stage_inst_dmem_n2358, MEM_stage_inst_dmem_n2357, MEM_stage_inst_dmem_n2356, MEM_stage_inst_dmem_n2355, MEM_stage_inst_dmem_n2354, MEM_stage_inst_dmem_n2353, MEM_stage_inst_dmem_n2352, MEM_stage_inst_dmem_n2351, MEM_stage_inst_dmem_n2350, MEM_stage_inst_dmem_n2349, MEM_stage_inst_dmem_n2348, MEM_stage_inst_dmem_n2347, MEM_stage_inst_dmem_n2346, MEM_stage_inst_dmem_n2345, MEM_stage_inst_dmem_n2344, MEM_stage_inst_dmem_n2343, MEM_stage_inst_dmem_n2342, MEM_stage_inst_dmem_n2341, MEM_stage_inst_dmem_n2340, MEM_stage_inst_dmem_n2339, MEM_stage_inst_dmem_n2338, MEM_stage_inst_dmem_n2337, MEM_stage_inst_dmem_n2336, MEM_stage_inst_dmem_n2335, MEM_stage_inst_dmem_n2334, MEM_stage_inst_dmem_n2333, MEM_stage_inst_dmem_n2332, MEM_stage_inst_dmem_n2331, MEM_stage_inst_dmem_n2330, MEM_stage_inst_dmem_n2329, MEM_stage_inst_dmem_n2328, MEM_stage_inst_dmem_n2327, MEM_stage_inst_dmem_n2326, MEM_stage_inst_dmem_n2325, MEM_stage_inst_dmem_n2324, MEM_stage_inst_dmem_n2323, MEM_stage_inst_dmem_n2322, MEM_stage_inst_dmem_n2321, MEM_stage_inst_dmem_n2320, MEM_stage_inst_dmem_n2319, MEM_stage_inst_dmem_n2318, MEM_stage_inst_dmem_n2317, MEM_stage_inst_dmem_n2316, MEM_stage_inst_dmem_n2315, MEM_stage_inst_dmem_n2314, MEM_stage_inst_dmem_n2313, MEM_stage_inst_dmem_n2312, MEM_stage_inst_dmem_n2311, MEM_stage_inst_dmem_n2310, MEM_stage_inst_dmem_n2309, MEM_stage_inst_dmem_n2308, MEM_stage_inst_dmem_n2307, MEM_stage_inst_dmem_n2306, MEM_stage_inst_dmem_n2305, MEM_stage_inst_dmem_n2304, MEM_stage_inst_dmem_n2303, MEM_stage_inst_dmem_n2302, MEM_stage_inst_dmem_n2301, MEM_stage_inst_dmem_n2300, MEM_stage_inst_dmem_n2299, MEM_stage_inst_dmem_n2298, MEM_stage_inst_dmem_n2297, MEM_stage_inst_dmem_n2296, MEM_stage_inst_dmem_n2295, MEM_stage_inst_dmem_n2294, MEM_stage_inst_dmem_n2293, MEM_stage_inst_dmem_n2292, MEM_stage_inst_dmem_n2291, MEM_stage_inst_dmem_n2290, MEM_stage_inst_dmem_n2289, MEM_stage_inst_dmem_n2288, MEM_stage_inst_dmem_n2287, MEM_stage_inst_dmem_n2286, MEM_stage_inst_dmem_n2285, MEM_stage_inst_dmem_n2284, MEM_stage_inst_dmem_n2283, MEM_stage_inst_dmem_n2282, MEM_stage_inst_dmem_n2281, MEM_stage_inst_dmem_n2280, MEM_stage_inst_dmem_n2279, MEM_stage_inst_dmem_n2278, MEM_stage_inst_dmem_n2277, MEM_stage_inst_dmem_n2276, MEM_stage_inst_dmem_n2275, MEM_stage_inst_dmem_n2274, MEM_stage_inst_dmem_n2273, MEM_stage_inst_dmem_n2272, MEM_stage_inst_dmem_n2271, MEM_stage_inst_dmem_n2270, MEM_stage_inst_dmem_n2269, MEM_stage_inst_dmem_n2268, MEM_stage_inst_dmem_n2267, MEM_stage_inst_dmem_n2266, MEM_stage_inst_dmem_n2265, MEM_stage_inst_dmem_n2264, MEM_stage_inst_dmem_n2263, MEM_stage_inst_dmem_n2262, MEM_stage_inst_dmem_n2261, MEM_stage_inst_dmem_n2260, MEM_stage_inst_dmem_n2259, MEM_stage_inst_dmem_n2258, MEM_stage_inst_dmem_n2257, MEM_stage_inst_dmem_n2256, MEM_stage_inst_dmem_n2255, MEM_stage_inst_dmem_n2254, MEM_stage_inst_dmem_n2253, MEM_stage_inst_dmem_n2252, MEM_stage_inst_dmem_n2251, MEM_stage_inst_dmem_n2250, MEM_stage_inst_dmem_n2249, MEM_stage_inst_dmem_n2248, MEM_stage_inst_dmem_n2247, MEM_stage_inst_dmem_n2246, MEM_stage_inst_dmem_n2245, MEM_stage_inst_dmem_n2244, MEM_stage_inst_dmem_n2243, MEM_stage_inst_dmem_n2242, MEM_stage_inst_dmem_n2241, MEM_stage_inst_dmem_n2240, MEM_stage_inst_dmem_n2239, MEM_stage_inst_dmem_n2238, MEM_stage_inst_dmem_n2237, MEM_stage_inst_dmem_n2236, MEM_stage_inst_dmem_n2235, MEM_stage_inst_dmem_n2234, MEM_stage_inst_dmem_n2233, MEM_stage_inst_dmem_n2232, MEM_stage_inst_dmem_n2231, MEM_stage_inst_dmem_n2230, MEM_stage_inst_dmem_n2229, MEM_stage_inst_dmem_n2228, MEM_stage_inst_dmem_n2227, MEM_stage_inst_dmem_n2226, MEM_stage_inst_dmem_n2225, MEM_stage_inst_dmem_n2224, MEM_stage_inst_dmem_n2223, MEM_stage_inst_dmem_n2222, MEM_stage_inst_dmem_n2221, MEM_stage_inst_dmem_n2220, MEM_stage_inst_dmem_n2219, MEM_stage_inst_dmem_n2218, MEM_stage_inst_dmem_n2217, MEM_stage_inst_dmem_n2216, MEM_stage_inst_dmem_n2215, MEM_stage_inst_dmem_n2214, MEM_stage_inst_dmem_n2213, MEM_stage_inst_dmem_n2212, MEM_stage_inst_dmem_n2211, MEM_stage_inst_dmem_n2210, MEM_stage_inst_dmem_n2209, MEM_stage_inst_dmem_n2208, MEM_stage_inst_dmem_n2207, MEM_stage_inst_dmem_n2206, MEM_stage_inst_dmem_n2205, MEM_stage_inst_dmem_n2204, MEM_stage_inst_dmem_n2203, MEM_stage_inst_dmem_n2202, MEM_stage_inst_dmem_n2201, MEM_stage_inst_dmem_n2200, MEM_stage_inst_dmem_n2199, MEM_stage_inst_dmem_n2198, MEM_stage_inst_dmem_n2197, MEM_stage_inst_dmem_n2196, MEM_stage_inst_dmem_n2195, MEM_stage_inst_dmem_n2194, MEM_stage_inst_dmem_n2193, MEM_stage_inst_dmem_n2192, MEM_stage_inst_dmem_n2191, MEM_stage_inst_dmem_n2190, MEM_stage_inst_dmem_n2189, MEM_stage_inst_dmem_n2188, MEM_stage_inst_dmem_n2187, MEM_stage_inst_dmem_n2186, MEM_stage_inst_dmem_n2185, MEM_stage_inst_dmem_n2184, MEM_stage_inst_dmem_n2183, MEM_stage_inst_dmem_n2182, MEM_stage_inst_dmem_n2181, MEM_stage_inst_dmem_n2180, MEM_stage_inst_dmem_n2179, MEM_stage_inst_dmem_n2178, MEM_stage_inst_dmem_n2177, MEM_stage_inst_dmem_n2176, MEM_stage_inst_dmem_n2175, MEM_stage_inst_dmem_n2174, MEM_stage_inst_dmem_n2173, MEM_stage_inst_dmem_n2172, MEM_stage_inst_dmem_n2171, MEM_stage_inst_dmem_n2170, MEM_stage_inst_dmem_n2169, MEM_stage_inst_dmem_n2168, MEM_stage_inst_dmem_n2167, MEM_stage_inst_dmem_n2166, MEM_stage_inst_dmem_n2165, MEM_stage_inst_dmem_n2164, MEM_stage_inst_dmem_n2163, MEM_stage_inst_dmem_n2162, MEM_stage_inst_dmem_n2161, MEM_stage_inst_dmem_n2160, MEM_stage_inst_dmem_n2159, MEM_stage_inst_dmem_n2158, MEM_stage_inst_dmem_n2157, MEM_stage_inst_dmem_n2156, MEM_stage_inst_dmem_n2155, MEM_stage_inst_dmem_n2154, MEM_stage_inst_dmem_n2153, MEM_stage_inst_dmem_n2152, MEM_stage_inst_dmem_n2151, MEM_stage_inst_dmem_n2150, MEM_stage_inst_dmem_n2149, MEM_stage_inst_dmem_n2148, MEM_stage_inst_dmem_n2147, MEM_stage_inst_dmem_n2146, MEM_stage_inst_dmem_n2145, MEM_stage_inst_dmem_n2144, MEM_stage_inst_dmem_n2143, MEM_stage_inst_dmem_n2142, MEM_stage_inst_dmem_n2141, MEM_stage_inst_dmem_n2140, MEM_stage_inst_dmem_n2139, MEM_stage_inst_dmem_n2138, MEM_stage_inst_dmem_n2137, MEM_stage_inst_dmem_n2136, MEM_stage_inst_dmem_n2135, MEM_stage_inst_dmem_n2134, MEM_stage_inst_dmem_n2133, MEM_stage_inst_dmem_n2132, MEM_stage_inst_dmem_n2131, MEM_stage_inst_dmem_n2130, MEM_stage_inst_dmem_n2129, MEM_stage_inst_dmem_n2128, MEM_stage_inst_dmem_n2127, MEM_stage_inst_dmem_n2126, MEM_stage_inst_dmem_n2125, MEM_stage_inst_dmem_n2124, MEM_stage_inst_dmem_n2123, MEM_stage_inst_dmem_n2122, MEM_stage_inst_dmem_n2121, MEM_stage_inst_dmem_n2120, MEM_stage_inst_dmem_n2119, MEM_stage_inst_dmem_n2118, MEM_stage_inst_dmem_n2117, MEM_stage_inst_dmem_n2116, MEM_stage_inst_dmem_n2115, MEM_stage_inst_dmem_n2114, MEM_stage_inst_dmem_n2113, MEM_stage_inst_dmem_n2112, MEM_stage_inst_dmem_n2111, MEM_stage_inst_dmem_n2110, MEM_stage_inst_dmem_n2109, MEM_stage_inst_dmem_n2108, MEM_stage_inst_dmem_n2107, MEM_stage_inst_dmem_n2106, MEM_stage_inst_dmem_n2105, MEM_stage_inst_dmem_n2104, MEM_stage_inst_dmem_n2103, MEM_stage_inst_dmem_n2102, MEM_stage_inst_dmem_n2101, MEM_stage_inst_dmem_n2100, MEM_stage_inst_dmem_n2099, MEM_stage_inst_dmem_n2098, MEM_stage_inst_dmem_n2097, MEM_stage_inst_dmem_n2096, MEM_stage_inst_dmem_n2095, MEM_stage_inst_dmem_n2094, MEM_stage_inst_dmem_n2093, MEM_stage_inst_dmem_n2092, MEM_stage_inst_dmem_n2091, MEM_stage_inst_dmem_n2090, MEM_stage_inst_dmem_n2089, MEM_stage_inst_dmem_n2088, MEM_stage_inst_dmem_n2087, MEM_stage_inst_dmem_n2086, MEM_stage_inst_dmem_n2085, MEM_stage_inst_dmem_n2084, MEM_stage_inst_dmem_n2083, MEM_stage_inst_dmem_n2082, MEM_stage_inst_dmem_n2081, MEM_stage_inst_dmem_n2080, MEM_stage_inst_dmem_n2079, MEM_stage_inst_dmem_n2078, MEM_stage_inst_dmem_n2077, MEM_stage_inst_dmem_n2076, MEM_stage_inst_dmem_n2075, MEM_stage_inst_dmem_n2074, MEM_stage_inst_dmem_n2073, MEM_stage_inst_dmem_n2072, MEM_stage_inst_dmem_n2071, MEM_stage_inst_dmem_n2070, MEM_stage_inst_dmem_n2069, MEM_stage_inst_dmem_n2068, MEM_stage_inst_dmem_n2067, MEM_stage_inst_dmem_n2066, MEM_stage_inst_dmem_n2065, MEM_stage_inst_dmem_n2064, MEM_stage_inst_dmem_n2063, MEM_stage_inst_dmem_n2062, MEM_stage_inst_dmem_n2061, MEM_stage_inst_dmem_n2060, MEM_stage_inst_dmem_n2059, MEM_stage_inst_dmem_n2058, MEM_stage_inst_dmem_n2057, MEM_stage_inst_dmem_n2056, MEM_stage_inst_dmem_n2055, MEM_stage_inst_dmem_n2054, MEM_stage_inst_dmem_n2053, MEM_stage_inst_dmem_n2052, MEM_stage_inst_dmem_n2051, MEM_stage_inst_dmem_n2050, MEM_stage_inst_dmem_n2049, MEM_stage_inst_dmem_n2048, MEM_stage_inst_dmem_n2047, MEM_stage_inst_dmem_n2046, MEM_stage_inst_dmem_n2045, MEM_stage_inst_dmem_n2044, MEM_stage_inst_dmem_n2043, MEM_stage_inst_dmem_n2042, MEM_stage_inst_dmem_n2041, MEM_stage_inst_dmem_n2040, MEM_stage_inst_dmem_n2039, MEM_stage_inst_dmem_n2038, MEM_stage_inst_dmem_n2037, MEM_stage_inst_dmem_n2036, MEM_stage_inst_dmem_n2035, MEM_stage_inst_dmem_n2034, MEM_stage_inst_dmem_n2033, MEM_stage_inst_dmem_n2032, MEM_stage_inst_dmem_n2031, MEM_stage_inst_dmem_n2030, MEM_stage_inst_dmem_n2029, MEM_stage_inst_dmem_n2028, MEM_stage_inst_dmem_n2027, MEM_stage_inst_dmem_n2026, MEM_stage_inst_dmem_n2025, MEM_stage_inst_dmem_n2024, MEM_stage_inst_dmem_n2023, MEM_stage_inst_dmem_n2022, MEM_stage_inst_dmem_n2021, MEM_stage_inst_dmem_n2020, MEM_stage_inst_dmem_n2019, MEM_stage_inst_dmem_n2018, MEM_stage_inst_dmem_n2017, MEM_stage_inst_dmem_n2016, MEM_stage_inst_dmem_n2015, MEM_stage_inst_dmem_n2014, MEM_stage_inst_dmem_n2013, MEM_stage_inst_dmem_n2012, MEM_stage_inst_dmem_n2011, MEM_stage_inst_dmem_n2010, MEM_stage_inst_dmem_n2009, MEM_stage_inst_dmem_n2008, MEM_stage_inst_dmem_n2007, MEM_stage_inst_dmem_n2006, MEM_stage_inst_dmem_n2005, MEM_stage_inst_dmem_n2004, MEM_stage_inst_dmem_n2003, MEM_stage_inst_dmem_n2002, MEM_stage_inst_dmem_n2001, MEM_stage_inst_dmem_n2000, MEM_stage_inst_dmem_n1999, MEM_stage_inst_dmem_n1998, MEM_stage_inst_dmem_n1997, MEM_stage_inst_dmem_n1996, MEM_stage_inst_dmem_n1995, MEM_stage_inst_dmem_n1994, MEM_stage_inst_dmem_n1993, MEM_stage_inst_dmem_n1992, MEM_stage_inst_dmem_n1991, MEM_stage_inst_dmem_n1990, MEM_stage_inst_dmem_n1989, MEM_stage_inst_dmem_n1988, MEM_stage_inst_dmem_n1987, MEM_stage_inst_dmem_n1986, MEM_stage_inst_dmem_n1985, MEM_stage_inst_dmem_n1984, MEM_stage_inst_dmem_n1983, MEM_stage_inst_dmem_n1982, MEM_stage_inst_dmem_n1981, MEM_stage_inst_dmem_n1980, MEM_stage_inst_dmem_n1979, MEM_stage_inst_dmem_n1978, MEM_stage_inst_dmem_n1977, MEM_stage_inst_dmem_n1976, MEM_stage_inst_dmem_n1975, MEM_stage_inst_dmem_n1974, MEM_stage_inst_dmem_n1973, MEM_stage_inst_dmem_n1972, MEM_stage_inst_dmem_n1971, MEM_stage_inst_dmem_n1970, MEM_stage_inst_dmem_n1969, MEM_stage_inst_dmem_n1968, MEM_stage_inst_dmem_n1967, MEM_stage_inst_dmem_n1966, MEM_stage_inst_dmem_n1965, MEM_stage_inst_dmem_n1964, MEM_stage_inst_dmem_n1963, MEM_stage_inst_dmem_n1962, MEM_stage_inst_dmem_n1961, MEM_stage_inst_dmem_n1960, MEM_stage_inst_dmem_n1959, MEM_stage_inst_dmem_n1958, MEM_stage_inst_dmem_n1957, MEM_stage_inst_dmem_n1956, MEM_stage_inst_dmem_n1955, MEM_stage_inst_dmem_n1954, MEM_stage_inst_dmem_n1953, MEM_stage_inst_dmem_n1952, MEM_stage_inst_dmem_n1951, MEM_stage_inst_dmem_n1950, MEM_stage_inst_dmem_n1949, MEM_stage_inst_dmem_n1948, MEM_stage_inst_dmem_n1947, MEM_stage_inst_dmem_n1946, MEM_stage_inst_dmem_n1945, MEM_stage_inst_dmem_n1944, MEM_stage_inst_dmem_n1943, MEM_stage_inst_dmem_n1942, MEM_stage_inst_dmem_n1941, MEM_stage_inst_dmem_n1940, MEM_stage_inst_dmem_n1939, MEM_stage_inst_dmem_n1938, MEM_stage_inst_dmem_n1937, MEM_stage_inst_dmem_n1936, MEM_stage_inst_dmem_n1935, MEM_stage_inst_dmem_n1934, MEM_stage_inst_dmem_n1933, MEM_stage_inst_dmem_n1932, MEM_stage_inst_dmem_n1931, MEM_stage_inst_dmem_n1930, MEM_stage_inst_dmem_n1929, MEM_stage_inst_dmem_n1928, MEM_stage_inst_dmem_n1927, MEM_stage_inst_dmem_n1926, MEM_stage_inst_dmem_n1925, MEM_stage_inst_dmem_n1924, MEM_stage_inst_dmem_n1923, MEM_stage_inst_dmem_n1922, MEM_stage_inst_dmem_n1921, MEM_stage_inst_dmem_n1920, MEM_stage_inst_dmem_n1919, MEM_stage_inst_dmem_n1918, MEM_stage_inst_dmem_n1917, MEM_stage_inst_dmem_n1916, MEM_stage_inst_dmem_n1915, MEM_stage_inst_dmem_n1914, MEM_stage_inst_dmem_n1913, MEM_stage_inst_dmem_n1912, MEM_stage_inst_dmem_n1911, MEM_stage_inst_dmem_n1910, MEM_stage_inst_dmem_n1909, MEM_stage_inst_dmem_n1908, MEM_stage_inst_dmem_n1907, MEM_stage_inst_dmem_n1906, MEM_stage_inst_dmem_n1905, MEM_stage_inst_dmem_n1904, MEM_stage_inst_dmem_n1903, MEM_stage_inst_dmem_n1902, MEM_stage_inst_dmem_n1901, MEM_stage_inst_dmem_n1900, MEM_stage_inst_dmem_n1899, MEM_stage_inst_dmem_n1898, MEM_stage_inst_dmem_n1897, MEM_stage_inst_dmem_n1896, MEM_stage_inst_dmem_n1895, MEM_stage_inst_dmem_n1894, MEM_stage_inst_dmem_n1893, MEM_stage_inst_dmem_n1892, MEM_stage_inst_dmem_n1891, MEM_stage_inst_dmem_n1890, MEM_stage_inst_dmem_n1889, MEM_stage_inst_dmem_n1888, MEM_stage_inst_dmem_n1887, MEM_stage_inst_dmem_n1886, MEM_stage_inst_dmem_n1885, MEM_stage_inst_dmem_n1884, MEM_stage_inst_dmem_n1883, MEM_stage_inst_dmem_n1882, MEM_stage_inst_dmem_n1881, MEM_stage_inst_dmem_n1880, MEM_stage_inst_dmem_n1879, MEM_stage_inst_dmem_n1878, MEM_stage_inst_dmem_n1877, MEM_stage_inst_dmem_n1876, MEM_stage_inst_dmem_n1875, MEM_stage_inst_dmem_n1874, MEM_stage_inst_dmem_n1873, MEM_stage_inst_dmem_n1872, MEM_stage_inst_dmem_n1871, MEM_stage_inst_dmem_n1870, MEM_stage_inst_dmem_n1869, MEM_stage_inst_dmem_n1868, MEM_stage_inst_dmem_n1867, MEM_stage_inst_dmem_n1866, MEM_stage_inst_dmem_n1865, MEM_stage_inst_dmem_n1864, MEM_stage_inst_dmem_n1863, MEM_stage_inst_dmem_n1862, MEM_stage_inst_dmem_n1861, MEM_stage_inst_dmem_n1860, MEM_stage_inst_dmem_n1859, MEM_stage_inst_dmem_n1858, MEM_stage_inst_dmem_n1857, MEM_stage_inst_dmem_n1856, MEM_stage_inst_dmem_n1855, MEM_stage_inst_dmem_n1854, MEM_stage_inst_dmem_n1853, MEM_stage_inst_dmem_n1852, MEM_stage_inst_dmem_n1851, MEM_stage_inst_dmem_n1850, MEM_stage_inst_dmem_n1849, MEM_stage_inst_dmem_n1848, MEM_stage_inst_dmem_n1847, MEM_stage_inst_dmem_n1846, MEM_stage_inst_dmem_n1845, MEM_stage_inst_dmem_n1844, MEM_stage_inst_dmem_n1843, MEM_stage_inst_dmem_n1842, MEM_stage_inst_dmem_n1841, MEM_stage_inst_dmem_n1840, MEM_stage_inst_dmem_n1839, MEM_stage_inst_dmem_n1838, MEM_stage_inst_dmem_n1837, MEM_stage_inst_dmem_n1836, MEM_stage_inst_dmem_n1835, MEM_stage_inst_dmem_n1834, MEM_stage_inst_dmem_n1833, MEM_stage_inst_dmem_n1832, MEM_stage_inst_dmem_n1831, MEM_stage_inst_dmem_n1830, MEM_stage_inst_dmem_n1829, MEM_stage_inst_dmem_n1828, MEM_stage_inst_dmem_n1827, MEM_stage_inst_dmem_n1826, MEM_stage_inst_dmem_n1825, MEM_stage_inst_dmem_n1824, MEM_stage_inst_dmem_n1823, MEM_stage_inst_dmem_n1822, MEM_stage_inst_dmem_n1821, MEM_stage_inst_dmem_n1820, MEM_stage_inst_dmem_n1819, MEM_stage_inst_dmem_n1818, MEM_stage_inst_dmem_n1817, MEM_stage_inst_dmem_n1816, MEM_stage_inst_dmem_n1815, MEM_stage_inst_dmem_n1814, MEM_stage_inst_dmem_n1813, MEM_stage_inst_dmem_n1812, MEM_stage_inst_dmem_n1811, MEM_stage_inst_dmem_n1810, MEM_stage_inst_dmem_n1809, MEM_stage_inst_dmem_n1808, MEM_stage_inst_dmem_n1807, MEM_stage_inst_dmem_n1806, MEM_stage_inst_dmem_n1805, MEM_stage_inst_dmem_n1804, MEM_stage_inst_dmem_n1803, MEM_stage_inst_dmem_n1802, MEM_stage_inst_dmem_n1801, MEM_stage_inst_dmem_n1800, MEM_stage_inst_dmem_n1799, MEM_stage_inst_dmem_n1798, MEM_stage_inst_dmem_n1797, MEM_stage_inst_dmem_n1796, MEM_stage_inst_dmem_n1795, MEM_stage_inst_dmem_n1794, MEM_stage_inst_dmem_n1793, MEM_stage_inst_dmem_n1792, MEM_stage_inst_dmem_n1791, MEM_stage_inst_dmem_n1790, MEM_stage_inst_dmem_n1789, MEM_stage_inst_dmem_n1788, MEM_stage_inst_dmem_n1787, MEM_stage_inst_dmem_n1786, MEM_stage_inst_dmem_n1785, MEM_stage_inst_dmem_n1784, MEM_stage_inst_dmem_n1783, MEM_stage_inst_dmem_n1782, MEM_stage_inst_dmem_n1781, MEM_stage_inst_dmem_n1780, MEM_stage_inst_dmem_n1779, MEM_stage_inst_dmem_n1778, MEM_stage_inst_dmem_n1777, MEM_stage_inst_dmem_n1776, MEM_stage_inst_dmem_n1775, MEM_stage_inst_dmem_n1774, MEM_stage_inst_dmem_n1773, MEM_stage_inst_dmem_n1772, MEM_stage_inst_dmem_n1771, MEM_stage_inst_dmem_n1770, MEM_stage_inst_dmem_n1769, MEM_stage_inst_dmem_n1768, MEM_stage_inst_dmem_n1767, MEM_stage_inst_dmem_n1766, MEM_stage_inst_dmem_n1765, MEM_stage_inst_dmem_n1764, MEM_stage_inst_dmem_n1763, MEM_stage_inst_dmem_n1762, MEM_stage_inst_dmem_n1761, MEM_stage_inst_dmem_n1760, MEM_stage_inst_dmem_n1759, MEM_stage_inst_dmem_n1758, MEM_stage_inst_dmem_n1757, MEM_stage_inst_dmem_n1756, MEM_stage_inst_dmem_n1755, MEM_stage_inst_dmem_n1754, MEM_stage_inst_dmem_n1753, MEM_stage_inst_dmem_n1752, MEM_stage_inst_dmem_n1751, MEM_stage_inst_dmem_n1750, MEM_stage_inst_dmem_n1749, MEM_stage_inst_dmem_n1748, MEM_stage_inst_dmem_n1747, MEM_stage_inst_dmem_n1746, MEM_stage_inst_dmem_n1745, MEM_stage_inst_dmem_n1744, MEM_stage_inst_dmem_n1743, MEM_stage_inst_dmem_n1742, MEM_stage_inst_dmem_n1741, MEM_stage_inst_dmem_n1740, MEM_stage_inst_dmem_n1739, MEM_stage_inst_dmem_n1738, MEM_stage_inst_dmem_n1737, MEM_stage_inst_dmem_n1736, MEM_stage_inst_dmem_n1735, MEM_stage_inst_dmem_n1734, MEM_stage_inst_dmem_n1733, MEM_stage_inst_dmem_n1732, MEM_stage_inst_dmem_n1731, MEM_stage_inst_dmem_n1730, MEM_stage_inst_dmem_n1729, MEM_stage_inst_dmem_n1728, MEM_stage_inst_dmem_n1727, MEM_stage_inst_dmem_n1726, MEM_stage_inst_dmem_n1725, MEM_stage_inst_dmem_n1724, MEM_stage_inst_dmem_n1723, MEM_stage_inst_dmem_n1722, MEM_stage_inst_dmem_n1721, MEM_stage_inst_dmem_n1720, MEM_stage_inst_dmem_n1719, MEM_stage_inst_dmem_n1718, MEM_stage_inst_dmem_n1717, MEM_stage_inst_dmem_n1716, MEM_stage_inst_dmem_n1715, MEM_stage_inst_dmem_n1714, MEM_stage_inst_dmem_n1713, MEM_stage_inst_dmem_n1712, MEM_stage_inst_dmem_n1711, MEM_stage_inst_dmem_n1710, MEM_stage_inst_dmem_n1709, MEM_stage_inst_dmem_n1708, MEM_stage_inst_dmem_n1707, MEM_stage_inst_dmem_n1706, MEM_stage_inst_dmem_n1705, MEM_stage_inst_dmem_n1704, MEM_stage_inst_dmem_n1703, MEM_stage_inst_dmem_n1702, MEM_stage_inst_dmem_n1701, MEM_stage_inst_dmem_n1700, MEM_stage_inst_dmem_n1699, MEM_stage_inst_dmem_n1698, MEM_stage_inst_dmem_n1697, MEM_stage_inst_dmem_n1696, MEM_stage_inst_dmem_n1695, MEM_stage_inst_dmem_n1694, MEM_stage_inst_dmem_n1693, MEM_stage_inst_dmem_n1692, MEM_stage_inst_dmem_n1691, MEM_stage_inst_dmem_n1690, MEM_stage_inst_dmem_n1689, MEM_stage_inst_dmem_n1688, MEM_stage_inst_dmem_n1687, MEM_stage_inst_dmem_n1686, MEM_stage_inst_dmem_n1685, MEM_stage_inst_dmem_n1684, MEM_stage_inst_dmem_n1683, MEM_stage_inst_dmem_n1682, MEM_stage_inst_dmem_n1681, MEM_stage_inst_dmem_n1680, MEM_stage_inst_dmem_n1679, MEM_stage_inst_dmem_n1678, MEM_stage_inst_dmem_n1677, MEM_stage_inst_dmem_n1676, MEM_stage_inst_dmem_n1675, MEM_stage_inst_dmem_n1674, MEM_stage_inst_dmem_n1673, MEM_stage_inst_dmem_n1672, MEM_stage_inst_dmem_n1671, MEM_stage_inst_dmem_n1670, MEM_stage_inst_dmem_n1669, MEM_stage_inst_dmem_n1668, MEM_stage_inst_dmem_n1667, MEM_stage_inst_dmem_n1666, MEM_stage_inst_dmem_n1665, MEM_stage_inst_dmem_n1664, MEM_stage_inst_dmem_n1663, MEM_stage_inst_dmem_n1662, MEM_stage_inst_dmem_n1661, MEM_stage_inst_dmem_n1660, MEM_stage_inst_dmem_n1659, MEM_stage_inst_dmem_n1658, MEM_stage_inst_dmem_n1657, MEM_stage_inst_dmem_n1656, MEM_stage_inst_dmem_n1655, MEM_stage_inst_dmem_n1654, MEM_stage_inst_dmem_n1653, MEM_stage_inst_dmem_n1652, MEM_stage_inst_dmem_n1651, MEM_stage_inst_dmem_n1650, MEM_stage_inst_dmem_n1649, MEM_stage_inst_dmem_n1648, MEM_stage_inst_dmem_n1647, MEM_stage_inst_dmem_n1646, MEM_stage_inst_dmem_n1645, MEM_stage_inst_dmem_n1644, MEM_stage_inst_dmem_n1643, MEM_stage_inst_dmem_n1642, MEM_stage_inst_dmem_n1641, MEM_stage_inst_dmem_n1640, MEM_stage_inst_dmem_n1639, MEM_stage_inst_dmem_n1638, MEM_stage_inst_dmem_n1637, MEM_stage_inst_dmem_n1636, MEM_stage_inst_dmem_n1635, MEM_stage_inst_dmem_n1634, MEM_stage_inst_dmem_n1633, MEM_stage_inst_dmem_n1632, MEM_stage_inst_dmem_n1631, MEM_stage_inst_dmem_n1630, MEM_stage_inst_dmem_n1629, MEM_stage_inst_dmem_n1628, MEM_stage_inst_dmem_n1627, MEM_stage_inst_dmem_n1626, MEM_stage_inst_dmem_n1625, MEM_stage_inst_dmem_n1624, MEM_stage_inst_dmem_n1623, MEM_stage_inst_dmem_n1622, MEM_stage_inst_dmem_n1621, MEM_stage_inst_dmem_n1620, MEM_stage_inst_dmem_n1619, MEM_stage_inst_dmem_n1618, MEM_stage_inst_dmem_n1617, MEM_stage_inst_dmem_n1616, MEM_stage_inst_dmem_n1615, MEM_stage_inst_dmem_n1614, MEM_stage_inst_dmem_n1613, MEM_stage_inst_dmem_n1612, MEM_stage_inst_dmem_n1611, MEM_stage_inst_dmem_n1610, MEM_stage_inst_dmem_n1609, MEM_stage_inst_dmem_n1608, MEM_stage_inst_dmem_n1607, MEM_stage_inst_dmem_n1606, MEM_stage_inst_dmem_n1605, MEM_stage_inst_dmem_n1604, MEM_stage_inst_dmem_n1603, MEM_stage_inst_dmem_n1602, MEM_stage_inst_dmem_n1601, MEM_stage_inst_dmem_n1600, MEM_stage_inst_dmem_n1599, MEM_stage_inst_dmem_n1598, MEM_stage_inst_dmem_n1597, MEM_stage_inst_dmem_n1596, MEM_stage_inst_dmem_n1595, MEM_stage_inst_dmem_n1594, MEM_stage_inst_dmem_n1593, MEM_stage_inst_dmem_n1592, MEM_stage_inst_dmem_n1591, MEM_stage_inst_dmem_n1590, MEM_stage_inst_dmem_n1589, MEM_stage_inst_dmem_n1588, MEM_stage_inst_dmem_n1587, MEM_stage_inst_dmem_n1586, MEM_stage_inst_dmem_n1585, MEM_stage_inst_dmem_n1584, MEM_stage_inst_dmem_n1583, MEM_stage_inst_dmem_n1582, MEM_stage_inst_dmem_n1581, MEM_stage_inst_dmem_n1580, MEM_stage_inst_dmem_n1579, MEM_stage_inst_dmem_n1578, MEM_stage_inst_dmem_n1577, MEM_stage_inst_dmem_n1576, MEM_stage_inst_dmem_n1575, MEM_stage_inst_dmem_n1574, MEM_stage_inst_dmem_n1573, MEM_stage_inst_dmem_n1572, MEM_stage_inst_dmem_n1571, MEM_stage_inst_dmem_n1570, MEM_stage_inst_dmem_n1569, MEM_stage_inst_dmem_n1568, MEM_stage_inst_dmem_n1567, MEM_stage_inst_dmem_n1566, MEM_stage_inst_dmem_n1565, MEM_stage_inst_dmem_n1564, MEM_stage_inst_dmem_n1563, MEM_stage_inst_dmem_n1562, MEM_stage_inst_dmem_n1561, MEM_stage_inst_dmem_n1560, MEM_stage_inst_dmem_n1559, MEM_stage_inst_dmem_n1558, MEM_stage_inst_dmem_n1557, MEM_stage_inst_dmem_n1556, MEM_stage_inst_dmem_n1555, MEM_stage_inst_dmem_n1554, MEM_stage_inst_dmem_n1553, MEM_stage_inst_dmem_n1552, MEM_stage_inst_dmem_n1551, MEM_stage_inst_dmem_n1550, MEM_stage_inst_dmem_n1549, MEM_stage_inst_dmem_n1548, MEM_stage_inst_dmem_n1547, MEM_stage_inst_dmem_n1546, MEM_stage_inst_dmem_n1545, MEM_stage_inst_dmem_n1544, MEM_stage_inst_dmem_n1543, MEM_stage_inst_dmem_n1542, MEM_stage_inst_dmem_n1541, MEM_stage_inst_dmem_n1540, MEM_stage_inst_dmem_n1539, MEM_stage_inst_dmem_n1538, MEM_stage_inst_dmem_n1537, MEM_stage_inst_dmem_n1536, MEM_stage_inst_dmem_n1535, MEM_stage_inst_dmem_n1534, MEM_stage_inst_dmem_n1533, MEM_stage_inst_dmem_n1532, MEM_stage_inst_dmem_n1531, MEM_stage_inst_dmem_n1530, MEM_stage_inst_dmem_n1529, MEM_stage_inst_dmem_n1528, MEM_stage_inst_dmem_n1527, MEM_stage_inst_dmem_n1526, MEM_stage_inst_dmem_n1525, MEM_stage_inst_dmem_n1524, MEM_stage_inst_dmem_n1523, MEM_stage_inst_dmem_n1522, MEM_stage_inst_dmem_n1521, MEM_stage_inst_dmem_n1520, MEM_stage_inst_dmem_n1519, MEM_stage_inst_dmem_n1518, MEM_stage_inst_dmem_n1517, MEM_stage_inst_dmem_n1516, MEM_stage_inst_dmem_n1515, MEM_stage_inst_dmem_n1514, MEM_stage_inst_dmem_n1513, MEM_stage_inst_dmem_n1512, MEM_stage_inst_dmem_n1511, MEM_stage_inst_dmem_n1510, MEM_stage_inst_dmem_n1509, MEM_stage_inst_dmem_n1508, MEM_stage_inst_dmem_n1507, MEM_stage_inst_dmem_n1506, MEM_stage_inst_dmem_n1505, MEM_stage_inst_dmem_n1504, MEM_stage_inst_dmem_n1503, MEM_stage_inst_dmem_n1502, MEM_stage_inst_dmem_n1501, MEM_stage_inst_dmem_n1500, MEM_stage_inst_dmem_n1499, MEM_stage_inst_dmem_n1498, MEM_stage_inst_dmem_n1497, MEM_stage_inst_dmem_n1496, MEM_stage_inst_dmem_n1495, MEM_stage_inst_dmem_n1494, MEM_stage_inst_dmem_n1493, MEM_stage_inst_dmem_n1492, MEM_stage_inst_dmem_n1491, MEM_stage_inst_dmem_n1490, MEM_stage_inst_dmem_n1489, MEM_stage_inst_dmem_n1488, MEM_stage_inst_dmem_n1487, MEM_stage_inst_dmem_n1486, MEM_stage_inst_dmem_n1485, MEM_stage_inst_dmem_n1484, MEM_stage_inst_dmem_n1483, MEM_stage_inst_dmem_n1482, MEM_stage_inst_dmem_n1481, MEM_stage_inst_dmem_n1480, MEM_stage_inst_dmem_n1479, MEM_stage_inst_dmem_n1478, MEM_stage_inst_dmem_n1477, MEM_stage_inst_dmem_n1476, MEM_stage_inst_dmem_n1475, MEM_stage_inst_dmem_n1474, MEM_stage_inst_dmem_n1473, MEM_stage_inst_dmem_n1472, MEM_stage_inst_dmem_n1471, MEM_stage_inst_dmem_n1470, MEM_stage_inst_dmem_n1469, MEM_stage_inst_dmem_n1468, MEM_stage_inst_dmem_n1467, MEM_stage_inst_dmem_n1466, MEM_stage_inst_dmem_n1465, MEM_stage_inst_dmem_n1464, MEM_stage_inst_dmem_n1463, MEM_stage_inst_dmem_n1462, MEM_stage_inst_dmem_n1461, MEM_stage_inst_dmem_n1460, MEM_stage_inst_dmem_n1459, MEM_stage_inst_dmem_n1458, MEM_stage_inst_dmem_n1457, MEM_stage_inst_dmem_n1456, MEM_stage_inst_dmem_n1455, MEM_stage_inst_dmem_n1454, MEM_stage_inst_dmem_n1453, MEM_stage_inst_dmem_n1452, MEM_stage_inst_dmem_n1451, MEM_stage_inst_dmem_n1450, MEM_stage_inst_dmem_n1449, MEM_stage_inst_dmem_n1448, MEM_stage_inst_dmem_n1447, MEM_stage_inst_dmem_n1446, MEM_stage_inst_dmem_n1445, MEM_stage_inst_dmem_n1444, MEM_stage_inst_dmem_n1443, MEM_stage_inst_dmem_n1442, MEM_stage_inst_dmem_n1441, MEM_stage_inst_dmem_n1440, MEM_stage_inst_dmem_n1439, MEM_stage_inst_dmem_n1438, MEM_stage_inst_dmem_n1437, MEM_stage_inst_dmem_n1436, MEM_stage_inst_dmem_n1435, MEM_stage_inst_dmem_n1434, MEM_stage_inst_dmem_n1433, MEM_stage_inst_dmem_n1432, MEM_stage_inst_dmem_n1431, MEM_stage_inst_dmem_n1430, MEM_stage_inst_dmem_n1429, MEM_stage_inst_dmem_n1428, MEM_stage_inst_dmem_n1427, MEM_stage_inst_dmem_n1426, MEM_stage_inst_dmem_n1425, MEM_stage_inst_dmem_n1424, MEM_stage_inst_dmem_n1423, MEM_stage_inst_dmem_n1422, MEM_stage_inst_dmem_n1421, MEM_stage_inst_dmem_n1420, MEM_stage_inst_dmem_n1419, MEM_stage_inst_dmem_n1418, MEM_stage_inst_dmem_n1417, MEM_stage_inst_dmem_n1416, MEM_stage_inst_dmem_n1415, MEM_stage_inst_dmem_n1414, MEM_stage_inst_dmem_n1413, MEM_stage_inst_dmem_n1412, MEM_stage_inst_dmem_n1411, MEM_stage_inst_dmem_n1410, MEM_stage_inst_dmem_n1409, MEM_stage_inst_dmem_n1408, MEM_stage_inst_dmem_n1407, MEM_stage_inst_dmem_n1406, MEM_stage_inst_dmem_n1405, MEM_stage_inst_dmem_n1404, MEM_stage_inst_dmem_n1403, MEM_stage_inst_dmem_n1402, MEM_stage_inst_dmem_n1401, MEM_stage_inst_dmem_n1400, MEM_stage_inst_dmem_n1399, MEM_stage_inst_dmem_n1398, MEM_stage_inst_dmem_n1397, MEM_stage_inst_dmem_n1396, MEM_stage_inst_dmem_n1395, MEM_stage_inst_dmem_n1394, MEM_stage_inst_dmem_n1393, MEM_stage_inst_dmem_n1392, MEM_stage_inst_dmem_n1391, MEM_stage_inst_dmem_n1390, MEM_stage_inst_dmem_n1389, MEM_stage_inst_dmem_n1388, MEM_stage_inst_dmem_n1387, MEM_stage_inst_dmem_n1386, MEM_stage_inst_dmem_n1385, MEM_stage_inst_dmem_n1384, MEM_stage_inst_dmem_n1383, MEM_stage_inst_dmem_n1382, MEM_stage_inst_dmem_n1381, MEM_stage_inst_dmem_n1380, MEM_stage_inst_dmem_n1379, MEM_stage_inst_dmem_n1378, MEM_stage_inst_dmem_n1377, MEM_stage_inst_dmem_n1376, MEM_stage_inst_dmem_n1375, MEM_stage_inst_dmem_n1374, MEM_stage_inst_dmem_n1373, MEM_stage_inst_dmem_n1372, MEM_stage_inst_dmem_n1371, MEM_stage_inst_dmem_n1370, MEM_stage_inst_dmem_n1369, MEM_stage_inst_dmem_n1368, MEM_stage_inst_dmem_n1367, MEM_stage_inst_dmem_n1366, MEM_stage_inst_dmem_n1365, MEM_stage_inst_dmem_n1364, MEM_stage_inst_dmem_n1363, MEM_stage_inst_dmem_n1362, MEM_stage_inst_dmem_n1361, MEM_stage_inst_dmem_n1360, MEM_stage_inst_dmem_n1359, MEM_stage_inst_dmem_n1358, MEM_stage_inst_dmem_n1357, MEM_stage_inst_dmem_n1356, MEM_stage_inst_dmem_n1355, MEM_stage_inst_dmem_n1354, MEM_stage_inst_dmem_n1353, MEM_stage_inst_dmem_n1352, MEM_stage_inst_dmem_n1351, MEM_stage_inst_dmem_n1350, MEM_stage_inst_dmem_n1349, MEM_stage_inst_dmem_n1348, MEM_stage_inst_dmem_n1347, MEM_stage_inst_dmem_n1346, MEM_stage_inst_dmem_n1345, MEM_stage_inst_dmem_n1344, MEM_stage_inst_dmem_n1343, MEM_stage_inst_dmem_n1342, MEM_stage_inst_dmem_n1341, MEM_stage_inst_dmem_n1340, MEM_stage_inst_dmem_n1339, MEM_stage_inst_dmem_n1338, MEM_stage_inst_dmem_n1337, MEM_stage_inst_dmem_n1336, MEM_stage_inst_dmem_n1335, MEM_stage_inst_dmem_n1334, MEM_stage_inst_dmem_n1333, MEM_stage_inst_dmem_n1332, MEM_stage_inst_dmem_n1331, MEM_stage_inst_dmem_n1330, MEM_stage_inst_dmem_n1329, MEM_stage_inst_dmem_n1328, MEM_stage_inst_dmem_n1327, MEM_stage_inst_dmem_n1326, MEM_stage_inst_dmem_n1325, MEM_stage_inst_dmem_n1324, MEM_stage_inst_dmem_n1323, MEM_stage_inst_dmem_n1322, MEM_stage_inst_dmem_n1321, MEM_stage_inst_dmem_n1320, MEM_stage_inst_dmem_n1319, MEM_stage_inst_dmem_n1318, MEM_stage_inst_dmem_n1317, MEM_stage_inst_dmem_n1316, MEM_stage_inst_dmem_n1315, MEM_stage_inst_dmem_n1314, MEM_stage_inst_dmem_n1313, MEM_stage_inst_dmem_n1312, MEM_stage_inst_dmem_n1311, MEM_stage_inst_dmem_n1310, MEM_stage_inst_dmem_n1309, MEM_stage_inst_dmem_n1308, MEM_stage_inst_dmem_n1307, MEM_stage_inst_dmem_n1306, MEM_stage_inst_dmem_n1305, MEM_stage_inst_dmem_n1304, MEM_stage_inst_dmem_n1303, MEM_stage_inst_dmem_n1302, MEM_stage_inst_dmem_n1301, MEM_stage_inst_dmem_n1300, MEM_stage_inst_dmem_n1299, MEM_stage_inst_dmem_n1298, MEM_stage_inst_dmem_n1297, MEM_stage_inst_dmem_n1296, MEM_stage_inst_dmem_n1295, MEM_stage_inst_dmem_n1294, MEM_stage_inst_dmem_n1293, MEM_stage_inst_dmem_n1292, MEM_stage_inst_dmem_n1291, MEM_stage_inst_dmem_n1290, MEM_stage_inst_dmem_n1289, MEM_stage_inst_dmem_n1288, MEM_stage_inst_dmem_n1287, MEM_stage_inst_dmem_n1286, MEM_stage_inst_dmem_n1285, MEM_stage_inst_dmem_n1284, MEM_stage_inst_dmem_n1283, MEM_stage_inst_dmem_n1282, MEM_stage_inst_dmem_n1281, MEM_stage_inst_dmem_n1280, MEM_stage_inst_dmem_n1279, MEM_stage_inst_dmem_n1278, MEM_stage_inst_dmem_n1277, MEM_stage_inst_dmem_n1276, MEM_stage_inst_dmem_n1275, MEM_stage_inst_dmem_n1274, MEM_stage_inst_dmem_n1273, MEM_stage_inst_dmem_n1272, MEM_stage_inst_dmem_n1271, MEM_stage_inst_dmem_n1270, MEM_stage_inst_dmem_n1269, MEM_stage_inst_dmem_n1268, MEM_stage_inst_dmem_n1267, MEM_stage_inst_dmem_n1266, MEM_stage_inst_dmem_n1265, MEM_stage_inst_dmem_n1264, MEM_stage_inst_dmem_n1263, MEM_stage_inst_dmem_n1262, MEM_stage_inst_dmem_n1261, MEM_stage_inst_dmem_n1260, MEM_stage_inst_dmem_n1259, MEM_stage_inst_dmem_n1258, MEM_stage_inst_dmem_n1257, MEM_stage_inst_dmem_n1256, MEM_stage_inst_dmem_n1255, MEM_stage_inst_dmem_n1254, MEM_stage_inst_dmem_n1253, MEM_stage_inst_dmem_n1252, MEM_stage_inst_dmem_n1251, MEM_stage_inst_dmem_n1250, MEM_stage_inst_dmem_n1249, MEM_stage_inst_dmem_n1248, MEM_stage_inst_dmem_n1247, MEM_stage_inst_dmem_n1246, MEM_stage_inst_dmem_n1245, MEM_stage_inst_dmem_n1244, MEM_stage_inst_dmem_n1243, MEM_stage_inst_dmem_n1242, MEM_stage_inst_dmem_n1241, MEM_stage_inst_dmem_n1240, MEM_stage_inst_dmem_n1239, MEM_stage_inst_dmem_n1238, MEM_stage_inst_dmem_n1237, MEM_stage_inst_dmem_n1236, MEM_stage_inst_dmem_n1235, MEM_stage_inst_dmem_n1234, MEM_stage_inst_dmem_n1233, MEM_stage_inst_dmem_n1232, MEM_stage_inst_dmem_n1231, MEM_stage_inst_dmem_n1230, MEM_stage_inst_dmem_n1229, MEM_stage_inst_dmem_n1228, MEM_stage_inst_dmem_n1227, MEM_stage_inst_dmem_n1226, MEM_stage_inst_dmem_n1225, MEM_stage_inst_dmem_n1224, MEM_stage_inst_dmem_n1223, MEM_stage_inst_dmem_n1222, MEM_stage_inst_dmem_n1221, MEM_stage_inst_dmem_n1220, MEM_stage_inst_dmem_n1219, MEM_stage_inst_dmem_n1218, MEM_stage_inst_dmem_n1217, MEM_stage_inst_dmem_n1216, MEM_stage_inst_dmem_n1215, MEM_stage_inst_dmem_n1214, MEM_stage_inst_dmem_n1213, MEM_stage_inst_dmem_n1212, MEM_stage_inst_dmem_n1211, MEM_stage_inst_dmem_n1210, MEM_stage_inst_dmem_n1209, MEM_stage_inst_dmem_n1208, MEM_stage_inst_dmem_n1207, MEM_stage_inst_dmem_n1206, MEM_stage_inst_dmem_n1205, MEM_stage_inst_dmem_n1204, MEM_stage_inst_dmem_n1203, MEM_stage_inst_dmem_n1202, MEM_stage_inst_dmem_n1201, MEM_stage_inst_dmem_n1200, MEM_stage_inst_dmem_n1199, MEM_stage_inst_dmem_n1198, MEM_stage_inst_dmem_n1197, MEM_stage_inst_dmem_n1196, MEM_stage_inst_dmem_n1195, MEM_stage_inst_dmem_n1194, MEM_stage_inst_dmem_n1193, MEM_stage_inst_dmem_n1192, MEM_stage_inst_dmem_n1191, MEM_stage_inst_dmem_n1190, MEM_stage_inst_dmem_n1189, MEM_stage_inst_dmem_n1188, MEM_stage_inst_dmem_n1187, MEM_stage_inst_dmem_n1186, MEM_stage_inst_dmem_n1185, MEM_stage_inst_dmem_n1184, MEM_stage_inst_dmem_n1183, MEM_stage_inst_dmem_n1182, MEM_stage_inst_dmem_n1181, MEM_stage_inst_dmem_n1180, MEM_stage_inst_dmem_n1179, MEM_stage_inst_dmem_n1178, MEM_stage_inst_dmem_n1177, MEM_stage_inst_dmem_n1176, MEM_stage_inst_dmem_n1175, MEM_stage_inst_dmem_n1174, MEM_stage_inst_dmem_n1173, MEM_stage_inst_dmem_n1172, MEM_stage_inst_dmem_n1171, MEM_stage_inst_dmem_n1170, MEM_stage_inst_dmem_n1169, MEM_stage_inst_dmem_n1168, MEM_stage_inst_dmem_n1167, MEM_stage_inst_dmem_n1166, MEM_stage_inst_dmem_n1165, MEM_stage_inst_dmem_n1164, MEM_stage_inst_dmem_n1163, MEM_stage_inst_dmem_n1162, MEM_stage_inst_dmem_n1161, MEM_stage_inst_dmem_n1160, MEM_stage_inst_dmem_n1159, MEM_stage_inst_dmem_n1158, MEM_stage_inst_dmem_n1157, MEM_stage_inst_dmem_n1156, MEM_stage_inst_dmem_n1155, MEM_stage_inst_dmem_n1154, MEM_stage_inst_dmem_n1153, MEM_stage_inst_dmem_n1152, MEM_stage_inst_dmem_n1151, MEM_stage_inst_dmem_n1150, MEM_stage_inst_dmem_n1149, MEM_stage_inst_dmem_n1148, MEM_stage_inst_dmem_n1147, MEM_stage_inst_dmem_n1146, MEM_stage_inst_dmem_n1145, MEM_stage_inst_dmem_n1144, MEM_stage_inst_dmem_n1143, MEM_stage_inst_dmem_n1142, MEM_stage_inst_dmem_n1141, MEM_stage_inst_dmem_n1140, MEM_stage_inst_dmem_n1139, MEM_stage_inst_dmem_n1138, MEM_stage_inst_dmem_n1137, MEM_stage_inst_dmem_n1136, MEM_stage_inst_dmem_n1135, MEM_stage_inst_dmem_n1134, MEM_stage_inst_dmem_n1133, MEM_stage_inst_dmem_n1132, MEM_stage_inst_dmem_n1131, MEM_stage_inst_dmem_n1130, MEM_stage_inst_dmem_n1129, MEM_stage_inst_dmem_n1128, MEM_stage_inst_dmem_n1127, MEM_stage_inst_dmem_n1126, MEM_stage_inst_dmem_n1125, MEM_stage_inst_dmem_n1124, MEM_stage_inst_dmem_n1123, MEM_stage_inst_dmem_n1122, MEM_stage_inst_dmem_n1121, MEM_stage_inst_dmem_n1120, MEM_stage_inst_dmem_n1119, MEM_stage_inst_dmem_n1118, MEM_stage_inst_dmem_n1117, MEM_stage_inst_dmem_n1116, MEM_stage_inst_dmem_n1115, MEM_stage_inst_dmem_n1114, MEM_stage_inst_dmem_n1113, MEM_stage_inst_dmem_n1112, MEM_stage_inst_dmem_n1111, MEM_stage_inst_dmem_n1110, MEM_stage_inst_dmem_n1109, MEM_stage_inst_dmem_n1108, MEM_stage_inst_dmem_n1107, MEM_stage_inst_dmem_n1106, MEM_stage_inst_dmem_n1105, MEM_stage_inst_dmem_n1104, MEM_stage_inst_dmem_n1103, MEM_stage_inst_dmem_n1102, MEM_stage_inst_dmem_n1101, MEM_stage_inst_dmem_n1100, MEM_stage_inst_dmem_n1099, MEM_stage_inst_dmem_n1098, MEM_stage_inst_dmem_n1097, MEM_stage_inst_dmem_n1096, MEM_stage_inst_dmem_n1095, MEM_stage_inst_dmem_n1094, MEM_stage_inst_dmem_n1093, MEM_stage_inst_dmem_n1092, MEM_stage_inst_dmem_n1091, MEM_stage_inst_dmem_n1090, MEM_stage_inst_dmem_n1089, MEM_stage_inst_dmem_n1088, MEM_stage_inst_dmem_n1087, MEM_stage_inst_dmem_n1086, MEM_stage_inst_dmem_n1085, MEM_stage_inst_dmem_n1084, MEM_stage_inst_dmem_n1083, MEM_stage_inst_dmem_n1082, MEM_stage_inst_dmem_n1081, MEM_stage_inst_dmem_n1080, MEM_stage_inst_dmem_n1079, MEM_stage_inst_dmem_n1078, MEM_stage_inst_dmem_n1077, MEM_stage_inst_dmem_n1076, MEM_stage_inst_dmem_n1075, MEM_stage_inst_dmem_n1074, MEM_stage_inst_dmem_n1073, MEM_stage_inst_dmem_n1072, MEM_stage_inst_dmem_n1071, MEM_stage_inst_dmem_n1070, MEM_stage_inst_dmem_n1069, MEM_stage_inst_dmem_n1068, MEM_stage_inst_dmem_n1067, MEM_stage_inst_dmem_n1066, MEM_stage_inst_dmem_n1065, MEM_stage_inst_dmem_n1064, MEM_stage_inst_dmem_n1063, MEM_stage_inst_dmem_n1062, MEM_stage_inst_dmem_n1061, MEM_stage_inst_dmem_n1060, MEM_stage_inst_dmem_n1059, MEM_stage_inst_dmem_n1058, MEM_stage_inst_dmem_n1057, MEM_stage_inst_dmem_n1056, MEM_stage_inst_dmem_n1055, MEM_stage_inst_dmem_n1054, MEM_stage_inst_dmem_n1053, MEM_stage_inst_dmem_n1052, MEM_stage_inst_dmem_n1051, MEM_stage_inst_dmem_n1050, MEM_stage_inst_dmem_n1049, MEM_stage_inst_dmem_n1048, MEM_stage_inst_dmem_n1047, MEM_stage_inst_dmem_n1046, MEM_stage_inst_dmem_n1045, MEM_stage_inst_dmem_n1044, MEM_stage_inst_dmem_n1043, MEM_stage_inst_dmem_n1042, MEM_stage_inst_dmem_n1041, MEM_stage_inst_dmem_n1040, MEM_stage_inst_dmem_n1039, MEM_stage_inst_dmem_n1038, MEM_stage_inst_dmem_n1037, MEM_stage_inst_dmem_n1036, MEM_stage_inst_dmem_n1035, MEM_stage_inst_dmem_n1034, MEM_stage_inst_dmem_n1033, MEM_stage_inst_dmem_n1032, MEM_stage_inst_dmem_n1031, MEM_stage_inst_dmem_n1030, MEM_stage_inst_dmem_n1029, MEM_stage_inst_dmem_n1028, MEM_stage_inst_dmem_n1027, MEM_stage_inst_dmem_n1026, MEM_stage_inst_dmem_n1025, MEM_stage_inst_dmem_n1024, MEM_stage_inst_dmem_n1023, MEM_stage_inst_dmem_n1022, MEM_stage_inst_dmem_n1021, MEM_stage_inst_dmem_n1020, MEM_stage_inst_dmem_n1019, MEM_stage_inst_dmem_n1018, MEM_stage_inst_dmem_n1017, MEM_stage_inst_dmem_n1016, MEM_stage_inst_dmem_n1015, MEM_stage_inst_dmem_n1014, MEM_stage_inst_dmem_n1013, MEM_stage_inst_dmem_n1012, MEM_stage_inst_dmem_n1011, MEM_stage_inst_dmem_n1010, MEM_stage_inst_dmem_n1009, MEM_stage_inst_dmem_n1008, MEM_stage_inst_dmem_n1007, MEM_stage_inst_dmem_n1006, MEM_stage_inst_dmem_n1005, MEM_stage_inst_dmem_n1004, MEM_stage_inst_dmem_n1003, MEM_stage_inst_dmem_n1002, MEM_stage_inst_dmem_n1001, MEM_stage_inst_dmem_n1000, MEM_stage_inst_dmem_n999, MEM_stage_inst_dmem_n998, MEM_stage_inst_dmem_n997, MEM_stage_inst_dmem_n996, MEM_stage_inst_dmem_n995, MEM_stage_inst_dmem_n994, MEM_stage_inst_dmem_n993, MEM_stage_inst_dmem_n992, MEM_stage_inst_dmem_n991, MEM_stage_inst_dmem_n990, MEM_stage_inst_dmem_n989, MEM_stage_inst_dmem_n988, MEM_stage_inst_dmem_n987, MEM_stage_inst_dmem_n986, MEM_stage_inst_dmem_n985, MEM_stage_inst_dmem_n984, MEM_stage_inst_dmem_n983, MEM_stage_inst_dmem_n982, MEM_stage_inst_dmem_n981, MEM_stage_inst_dmem_n980, MEM_stage_inst_dmem_n979, MEM_stage_inst_dmem_n978, MEM_stage_inst_dmem_n977, MEM_stage_inst_dmem_n976, MEM_stage_inst_dmem_n975, MEM_stage_inst_dmem_n974, MEM_stage_inst_dmem_n973, MEM_stage_inst_dmem_n972, MEM_stage_inst_dmem_n971, MEM_stage_inst_dmem_n970, MEM_stage_inst_dmem_n969, MEM_stage_inst_dmem_n968, MEM_stage_inst_dmem_n967, MEM_stage_inst_dmem_n966, MEM_stage_inst_dmem_n965, MEM_stage_inst_dmem_n964, MEM_stage_inst_dmem_n963, MEM_stage_inst_dmem_n962, MEM_stage_inst_dmem_n961, MEM_stage_inst_dmem_n960, MEM_stage_inst_dmem_n959, MEM_stage_inst_dmem_n958, MEM_stage_inst_dmem_n957, MEM_stage_inst_dmem_n956, MEM_stage_inst_dmem_n955, MEM_stage_inst_dmem_n954, MEM_stage_inst_dmem_n953, MEM_stage_inst_dmem_n952, MEM_stage_inst_dmem_n951, MEM_stage_inst_dmem_n950, MEM_stage_inst_dmem_n949, MEM_stage_inst_dmem_n948, MEM_stage_inst_dmem_n947, MEM_stage_inst_dmem_n946, MEM_stage_inst_dmem_n945, MEM_stage_inst_dmem_n944, MEM_stage_inst_dmem_n943, MEM_stage_inst_dmem_n942, MEM_stage_inst_dmem_n941, MEM_stage_inst_dmem_n940, MEM_stage_inst_dmem_n939, MEM_stage_inst_dmem_n938, MEM_stage_inst_dmem_n937, MEM_stage_inst_dmem_n936, MEM_stage_inst_dmem_n935, MEM_stage_inst_dmem_n934, MEM_stage_inst_dmem_n933, MEM_stage_inst_dmem_n932, MEM_stage_inst_dmem_n931, MEM_stage_inst_dmem_n930, MEM_stage_inst_dmem_n929, MEM_stage_inst_dmem_n928, MEM_stage_inst_dmem_n927, MEM_stage_inst_dmem_n926, MEM_stage_inst_dmem_n925, MEM_stage_inst_dmem_n924, MEM_stage_inst_dmem_n923, MEM_stage_inst_dmem_n922, MEM_stage_inst_dmem_n921, MEM_stage_inst_dmem_n920, MEM_stage_inst_dmem_n919, MEM_stage_inst_dmem_n918, MEM_stage_inst_dmem_n917, MEM_stage_inst_dmem_n916, MEM_stage_inst_dmem_n915, MEM_stage_inst_dmem_n914, MEM_stage_inst_dmem_n913, MEM_stage_inst_dmem_n912, MEM_stage_inst_dmem_n911, MEM_stage_inst_dmem_n910, MEM_stage_inst_dmem_n909, MEM_stage_inst_dmem_n908, MEM_stage_inst_dmem_n907, MEM_stage_inst_dmem_n906, MEM_stage_inst_dmem_n905, MEM_stage_inst_dmem_n904, MEM_stage_inst_dmem_n903, MEM_stage_inst_dmem_n902, MEM_stage_inst_dmem_n901, MEM_stage_inst_dmem_n900, MEM_stage_inst_dmem_n899, MEM_stage_inst_dmem_n898, MEM_stage_inst_dmem_n897, MEM_stage_inst_dmem_n896, MEM_stage_inst_dmem_n895, MEM_stage_inst_dmem_n894, MEM_stage_inst_dmem_n893, MEM_stage_inst_dmem_n892, MEM_stage_inst_dmem_n891, MEM_stage_inst_dmem_n890, MEM_stage_inst_dmem_n889, MEM_stage_inst_dmem_n888, MEM_stage_inst_dmem_n887, MEM_stage_inst_dmem_n886, MEM_stage_inst_dmem_n885, MEM_stage_inst_dmem_n884, MEM_stage_inst_dmem_n883, MEM_stage_inst_dmem_n882, MEM_stage_inst_dmem_n881, MEM_stage_inst_dmem_n880, MEM_stage_inst_dmem_n879, MEM_stage_inst_dmem_n878, MEM_stage_inst_dmem_n877, MEM_stage_inst_dmem_n876, MEM_stage_inst_dmem_n875, MEM_stage_inst_dmem_n874, MEM_stage_inst_dmem_n873, MEM_stage_inst_dmem_n872, MEM_stage_inst_dmem_n871, MEM_stage_inst_dmem_n870, MEM_stage_inst_dmem_n869, MEM_stage_inst_dmem_n868, MEM_stage_inst_dmem_n867, MEM_stage_inst_dmem_n866, MEM_stage_inst_dmem_n865, MEM_stage_inst_dmem_n864, MEM_stage_inst_dmem_n863, MEM_stage_inst_dmem_n862, MEM_stage_inst_dmem_n861, MEM_stage_inst_dmem_n860, MEM_stage_inst_dmem_n859, MEM_stage_inst_dmem_n858, MEM_stage_inst_dmem_n857, MEM_stage_inst_dmem_n856, MEM_stage_inst_dmem_n855, MEM_stage_inst_dmem_n854, MEM_stage_inst_dmem_n853, MEM_stage_inst_dmem_n852, MEM_stage_inst_dmem_n851, MEM_stage_inst_dmem_n850, MEM_stage_inst_dmem_n849, MEM_stage_inst_dmem_n848, MEM_stage_inst_dmem_n847, MEM_stage_inst_dmem_n846, MEM_stage_inst_dmem_n845, MEM_stage_inst_dmem_n844, MEM_stage_inst_dmem_n843, MEM_stage_inst_dmem_n842, MEM_stage_inst_dmem_n841, MEM_stage_inst_dmem_n840, MEM_stage_inst_dmem_n839, MEM_stage_inst_dmem_n838, MEM_stage_inst_dmem_n837, MEM_stage_inst_dmem_n836, MEM_stage_inst_dmem_n835, MEM_stage_inst_dmem_n834, MEM_stage_inst_dmem_n833, MEM_stage_inst_dmem_n832, MEM_stage_inst_dmem_n831, MEM_stage_inst_dmem_n830, MEM_stage_inst_dmem_n829, MEM_stage_inst_dmem_n828, MEM_stage_inst_dmem_n827, MEM_stage_inst_dmem_n826, MEM_stage_inst_dmem_n825, MEM_stage_inst_dmem_n824, MEM_stage_inst_dmem_n823, MEM_stage_inst_dmem_n822, MEM_stage_inst_dmem_n821, MEM_stage_inst_dmem_n820, MEM_stage_inst_dmem_n819, MEM_stage_inst_dmem_n818, MEM_stage_inst_dmem_n817, MEM_stage_inst_dmem_n816, MEM_stage_inst_dmem_n815, MEM_stage_inst_dmem_n814, MEM_stage_inst_dmem_n813, MEM_stage_inst_dmem_n812, MEM_stage_inst_dmem_n811, MEM_stage_inst_dmem_n810, MEM_stage_inst_dmem_n809, MEM_stage_inst_dmem_n808, MEM_stage_inst_dmem_n807, MEM_stage_inst_dmem_n806, MEM_stage_inst_dmem_n805, MEM_stage_inst_dmem_n804, MEM_stage_inst_dmem_n803, MEM_stage_inst_dmem_n802, MEM_stage_inst_dmem_n801, MEM_stage_inst_dmem_n800, MEM_stage_inst_dmem_n799, MEM_stage_inst_dmem_n798, MEM_stage_inst_dmem_n797, MEM_stage_inst_dmem_n796, MEM_stage_inst_dmem_n795, MEM_stage_inst_dmem_n794, MEM_stage_inst_dmem_n793, MEM_stage_inst_dmem_n792, MEM_stage_inst_dmem_n791, MEM_stage_inst_dmem_n790, MEM_stage_inst_dmem_n789, MEM_stage_inst_dmem_n788, MEM_stage_inst_dmem_n787, MEM_stage_inst_dmem_n786, MEM_stage_inst_dmem_n785, MEM_stage_inst_dmem_n784, MEM_stage_inst_dmem_n783, MEM_stage_inst_dmem_n782, MEM_stage_inst_dmem_n781, MEM_stage_inst_dmem_n780, MEM_stage_inst_dmem_n779, MEM_stage_inst_dmem_n778, MEM_stage_inst_dmem_n777, MEM_stage_inst_dmem_n776, MEM_stage_inst_dmem_n775, MEM_stage_inst_dmem_n774, MEM_stage_inst_dmem_n773, MEM_stage_inst_dmem_n772, MEM_stage_inst_dmem_n771, MEM_stage_inst_dmem_n770, MEM_stage_inst_dmem_n769, MEM_stage_inst_dmem_n768, MEM_stage_inst_dmem_n767, MEM_stage_inst_dmem_n766, MEM_stage_inst_dmem_n765, MEM_stage_inst_dmem_n764, MEM_stage_inst_dmem_n763, MEM_stage_inst_dmem_n762, MEM_stage_inst_dmem_n761, MEM_stage_inst_dmem_n760, MEM_stage_inst_dmem_n759, MEM_stage_inst_dmem_n758, MEM_stage_inst_dmem_n757, MEM_stage_inst_dmem_n756, MEM_stage_inst_dmem_n755, MEM_stage_inst_dmem_n754, MEM_stage_inst_dmem_n753, MEM_stage_inst_dmem_n752, MEM_stage_inst_dmem_n751, MEM_stage_inst_dmem_n750, MEM_stage_inst_dmem_n749, MEM_stage_inst_dmem_n748, MEM_stage_inst_dmem_n747, MEM_stage_inst_dmem_n746, MEM_stage_inst_dmem_n745, MEM_stage_inst_dmem_n744, MEM_stage_inst_dmem_n743, MEM_stage_inst_dmem_n742, MEM_stage_inst_dmem_n741, MEM_stage_inst_dmem_n740, MEM_stage_inst_dmem_n739, MEM_stage_inst_dmem_n738, MEM_stage_inst_dmem_n737, MEM_stage_inst_dmem_n736, MEM_stage_inst_dmem_n735, MEM_stage_inst_dmem_n734, MEM_stage_inst_dmem_n733, MEM_stage_inst_dmem_n732, MEM_stage_inst_dmem_n731, MEM_stage_inst_dmem_n730, MEM_stage_inst_dmem_n729, MEM_stage_inst_dmem_n728, MEM_stage_inst_dmem_n727, MEM_stage_inst_dmem_n726, MEM_stage_inst_dmem_n725, MEM_stage_inst_dmem_n724, MEM_stage_inst_dmem_n723, MEM_stage_inst_dmem_n722, MEM_stage_inst_dmem_n721, MEM_stage_inst_dmem_n720, MEM_stage_inst_dmem_n719, MEM_stage_inst_dmem_n718, MEM_stage_inst_dmem_n717, MEM_stage_inst_dmem_n716, MEM_stage_inst_dmem_n715, MEM_stage_inst_dmem_n714, MEM_stage_inst_dmem_n713, MEM_stage_inst_dmem_n712, MEM_stage_inst_dmem_n711, MEM_stage_inst_dmem_n710, MEM_stage_inst_dmem_n709, MEM_stage_inst_dmem_n708, MEM_stage_inst_dmem_n707, MEM_stage_inst_dmem_n706, MEM_stage_inst_dmem_n705, MEM_stage_inst_dmem_n704, MEM_stage_inst_dmem_n703, MEM_stage_inst_dmem_n702, MEM_stage_inst_dmem_n701, MEM_stage_inst_dmem_n700, MEM_stage_inst_dmem_n699, MEM_stage_inst_dmem_n698, MEM_stage_inst_dmem_n697, MEM_stage_inst_dmem_n696, MEM_stage_inst_dmem_n695, MEM_stage_inst_dmem_n694, MEM_stage_inst_dmem_n693, MEM_stage_inst_dmem_n692, MEM_stage_inst_dmem_n691, MEM_stage_inst_dmem_n690, MEM_stage_inst_dmem_n689, MEM_stage_inst_dmem_n688, MEM_stage_inst_dmem_n687, MEM_stage_inst_dmem_n686, MEM_stage_inst_dmem_n685, MEM_stage_inst_dmem_n684, MEM_stage_inst_dmem_n683, MEM_stage_inst_dmem_n682, MEM_stage_inst_dmem_n681, MEM_stage_inst_dmem_n680, MEM_stage_inst_dmem_n679, MEM_stage_inst_dmem_n678, MEM_stage_inst_dmem_n677, MEM_stage_inst_dmem_n676, MEM_stage_inst_dmem_n675, MEM_stage_inst_dmem_n674, MEM_stage_inst_dmem_n673, MEM_stage_inst_dmem_n672, MEM_stage_inst_dmem_n671, MEM_stage_inst_dmem_n670, MEM_stage_inst_dmem_n669, MEM_stage_inst_dmem_n668, MEM_stage_inst_dmem_n667, MEM_stage_inst_dmem_n666, MEM_stage_inst_dmem_n665, MEM_stage_inst_dmem_n664, MEM_stage_inst_dmem_n663, MEM_stage_inst_dmem_n662, MEM_stage_inst_dmem_n661, MEM_stage_inst_dmem_n660, MEM_stage_inst_dmem_n659, MEM_stage_inst_dmem_n658, MEM_stage_inst_dmem_n657, MEM_stage_inst_dmem_n656, MEM_stage_inst_dmem_n655, MEM_stage_inst_dmem_n654, MEM_stage_inst_dmem_n653, MEM_stage_inst_dmem_n652, MEM_stage_inst_dmem_n651, MEM_stage_inst_dmem_n650, MEM_stage_inst_dmem_n649, MEM_stage_inst_dmem_n648, MEM_stage_inst_dmem_n647, MEM_stage_inst_dmem_n646, MEM_stage_inst_dmem_n645, MEM_stage_inst_dmem_n644, MEM_stage_inst_dmem_n643, MEM_stage_inst_dmem_n642, MEM_stage_inst_dmem_n641, MEM_stage_inst_dmem_n640, MEM_stage_inst_dmem_n639, MEM_stage_inst_dmem_n638, MEM_stage_inst_dmem_n637, MEM_stage_inst_dmem_n636, MEM_stage_inst_dmem_n635, MEM_stage_inst_dmem_n634, MEM_stage_inst_dmem_n633, MEM_stage_inst_dmem_n632, MEM_stage_inst_dmem_n631, MEM_stage_inst_dmem_n630, MEM_stage_inst_dmem_n629, MEM_stage_inst_dmem_n628, MEM_stage_inst_dmem_n627, MEM_stage_inst_dmem_n626, MEM_stage_inst_dmem_n625, MEM_stage_inst_dmem_n624, MEM_stage_inst_dmem_n623, MEM_stage_inst_dmem_n622, MEM_stage_inst_dmem_n621, MEM_stage_inst_dmem_n620, MEM_stage_inst_dmem_n619, MEM_stage_inst_dmem_n618, MEM_stage_inst_dmem_n617, MEM_stage_inst_dmem_n616, MEM_stage_inst_dmem_n615, MEM_stage_inst_dmem_n614, MEM_stage_inst_dmem_n613, MEM_stage_inst_dmem_n612, MEM_stage_inst_dmem_n611, MEM_stage_inst_dmem_n610, MEM_stage_inst_dmem_n609, MEM_stage_inst_dmem_n608, MEM_stage_inst_dmem_n607, MEM_stage_inst_dmem_n606, MEM_stage_inst_dmem_n605, MEM_stage_inst_dmem_n604, MEM_stage_inst_dmem_n603, MEM_stage_inst_dmem_n602, MEM_stage_inst_dmem_n601, MEM_stage_inst_dmem_n600, MEM_stage_inst_dmem_n599, MEM_stage_inst_dmem_n598, MEM_stage_inst_dmem_n597, MEM_stage_inst_dmem_n596, MEM_stage_inst_dmem_n595, MEM_stage_inst_dmem_n594, MEM_stage_inst_dmem_n593, MEM_stage_inst_dmem_n592, MEM_stage_inst_dmem_n591, MEM_stage_inst_dmem_n590, MEM_stage_inst_dmem_n589, MEM_stage_inst_dmem_n588, MEM_stage_inst_dmem_n587, MEM_stage_inst_dmem_n586, MEM_stage_inst_dmem_n585, MEM_stage_inst_dmem_n584, MEM_stage_inst_dmem_n583, MEM_stage_inst_dmem_n582, MEM_stage_inst_dmem_n581, MEM_stage_inst_dmem_n580, MEM_stage_inst_dmem_n579, MEM_stage_inst_dmem_n578, MEM_stage_inst_dmem_n577, MEM_stage_inst_dmem_n576, MEM_stage_inst_dmem_n575, MEM_stage_inst_dmem_n574, MEM_stage_inst_dmem_n573, MEM_stage_inst_dmem_n572, MEM_stage_inst_dmem_n571, MEM_stage_inst_dmem_n570, MEM_stage_inst_dmem_n569, MEM_stage_inst_dmem_n568, MEM_stage_inst_dmem_n567, MEM_stage_inst_dmem_n566, MEM_stage_inst_dmem_n565, MEM_stage_inst_dmem_n564, MEM_stage_inst_dmem_n563, MEM_stage_inst_dmem_n562, MEM_stage_inst_dmem_n561, MEM_stage_inst_dmem_n560, MEM_stage_inst_dmem_n559, MEM_stage_inst_dmem_n558, MEM_stage_inst_dmem_n557, MEM_stage_inst_dmem_n556, MEM_stage_inst_dmem_n555, MEM_stage_inst_dmem_n554, MEM_stage_inst_dmem_n553, MEM_stage_inst_dmem_n552, MEM_stage_inst_dmem_n551, MEM_stage_inst_dmem_n550, MEM_stage_inst_dmem_n549, MEM_stage_inst_dmem_n548, MEM_stage_inst_dmem_n547, MEM_stage_inst_dmem_n546, MEM_stage_inst_dmem_n545, MEM_stage_inst_dmem_n544, MEM_stage_inst_dmem_n543, MEM_stage_inst_dmem_n542, MEM_stage_inst_dmem_n541, MEM_stage_inst_dmem_n540, MEM_stage_inst_dmem_n539, MEM_stage_inst_dmem_n538, MEM_stage_inst_dmem_n537, MEM_stage_inst_dmem_n536, MEM_stage_inst_dmem_n535, MEM_stage_inst_dmem_n534, MEM_stage_inst_dmem_n533, MEM_stage_inst_dmem_n532, MEM_stage_inst_dmem_n531, MEM_stage_inst_dmem_n530, MEM_stage_inst_dmem_n529, MEM_stage_inst_dmem_n528, MEM_stage_inst_dmem_n527, MEM_stage_inst_dmem_n526, MEM_stage_inst_dmem_n525, MEM_stage_inst_dmem_n524, MEM_stage_inst_dmem_n523, MEM_stage_inst_dmem_n522, MEM_stage_inst_dmem_n521, MEM_stage_inst_dmem_n520, MEM_stage_inst_dmem_n519, MEM_stage_inst_dmem_n518, MEM_stage_inst_dmem_n517, MEM_stage_inst_dmem_n516, MEM_stage_inst_dmem_n515, MEM_stage_inst_dmem_n514, MEM_stage_inst_dmem_n513, MEM_stage_inst_dmem_n512, MEM_stage_inst_dmem_n511, MEM_stage_inst_dmem_n510, MEM_stage_inst_dmem_n509, MEM_stage_inst_dmem_n508, MEM_stage_inst_dmem_n507, MEM_stage_inst_dmem_n506, MEM_stage_inst_dmem_n505, MEM_stage_inst_dmem_n504, MEM_stage_inst_dmem_n503, MEM_stage_inst_dmem_n502, MEM_stage_inst_dmem_n501, MEM_stage_inst_dmem_n500, MEM_stage_inst_dmem_n499, MEM_stage_inst_dmem_n498, MEM_stage_inst_dmem_n497, MEM_stage_inst_dmem_n496, MEM_stage_inst_dmem_n495, MEM_stage_inst_dmem_n494, MEM_stage_inst_dmem_n493, MEM_stage_inst_dmem_n492, MEM_stage_inst_dmem_n491, MEM_stage_inst_dmem_n490, MEM_stage_inst_dmem_n489, MEM_stage_inst_dmem_n488, MEM_stage_inst_dmem_n487, MEM_stage_inst_dmem_n486, MEM_stage_inst_dmem_n485, MEM_stage_inst_dmem_n484, MEM_stage_inst_dmem_n483, MEM_stage_inst_dmem_n482, MEM_stage_inst_dmem_n481, MEM_stage_inst_dmem_n480, MEM_stage_inst_dmem_n479, MEM_stage_inst_dmem_n478, MEM_stage_inst_dmem_n477, MEM_stage_inst_dmem_n476, MEM_stage_inst_dmem_n475, MEM_stage_inst_dmem_n474, MEM_stage_inst_dmem_n473, MEM_stage_inst_dmem_n472, MEM_stage_inst_dmem_n471, MEM_stage_inst_dmem_n470, MEM_stage_inst_dmem_n469, MEM_stage_inst_dmem_n468, MEM_stage_inst_dmem_n467, MEM_stage_inst_dmem_n466, MEM_stage_inst_dmem_n465, MEM_stage_inst_dmem_n464, MEM_stage_inst_dmem_n463, MEM_stage_inst_dmem_n462, MEM_stage_inst_dmem_n461, MEM_stage_inst_dmem_n460, MEM_stage_inst_dmem_n459, MEM_stage_inst_dmem_n458, MEM_stage_inst_dmem_n457, MEM_stage_inst_dmem_n456, MEM_stage_inst_dmem_n455, MEM_stage_inst_dmem_n454, MEM_stage_inst_dmem_n453, MEM_stage_inst_dmem_n452, MEM_stage_inst_dmem_n451, MEM_stage_inst_dmem_n450, MEM_stage_inst_dmem_n449, MEM_stage_inst_dmem_n448, MEM_stage_inst_dmem_n447, MEM_stage_inst_dmem_n446, MEM_stage_inst_dmem_n445, MEM_stage_inst_dmem_n444, MEM_stage_inst_dmem_n443, MEM_stage_inst_dmem_n442, MEM_stage_inst_dmem_n441, MEM_stage_inst_dmem_n440, MEM_stage_inst_dmem_n439, MEM_stage_inst_dmem_n438, MEM_stage_inst_dmem_n437, MEM_stage_inst_dmem_n436, MEM_stage_inst_dmem_n435, MEM_stage_inst_dmem_n434, MEM_stage_inst_dmem_n433, MEM_stage_inst_dmem_n432, MEM_stage_inst_dmem_n431, MEM_stage_inst_dmem_n430, MEM_stage_inst_dmem_n429, MEM_stage_inst_dmem_n428, MEM_stage_inst_dmem_n427, MEM_stage_inst_dmem_n426, MEM_stage_inst_dmem_n425, MEM_stage_inst_dmem_n424, MEM_stage_inst_dmem_n423, MEM_stage_inst_dmem_n422, MEM_stage_inst_dmem_n421, MEM_stage_inst_dmem_n420, MEM_stage_inst_dmem_n419, MEM_stage_inst_dmem_n418, MEM_stage_inst_dmem_n417, MEM_stage_inst_dmem_n416, MEM_stage_inst_dmem_n415, MEM_stage_inst_dmem_n414, MEM_stage_inst_dmem_n413, MEM_stage_inst_dmem_n412, MEM_stage_inst_dmem_n411, MEM_stage_inst_dmem_n410, MEM_stage_inst_dmem_n409, MEM_stage_inst_dmem_n408, MEM_stage_inst_dmem_n407, MEM_stage_inst_dmem_n406, MEM_stage_inst_dmem_n405, MEM_stage_inst_dmem_n404, MEM_stage_inst_dmem_n403, MEM_stage_inst_dmem_n402, MEM_stage_inst_dmem_n401, MEM_stage_inst_dmem_n400, MEM_stage_inst_dmem_n399, MEM_stage_inst_dmem_n398, MEM_stage_inst_dmem_n397, MEM_stage_inst_dmem_n396, MEM_stage_inst_dmem_n395, MEM_stage_inst_dmem_n394, MEM_stage_inst_dmem_n393, MEM_stage_inst_dmem_n392, MEM_stage_inst_dmem_n391, MEM_stage_inst_dmem_n390, MEM_stage_inst_dmem_n389, MEM_stage_inst_dmem_n388, MEM_stage_inst_dmem_n387, MEM_stage_inst_dmem_n386, MEM_stage_inst_dmem_n385, MEM_stage_inst_dmem_n384, MEM_stage_inst_dmem_n383, MEM_stage_inst_dmem_n382, MEM_stage_inst_dmem_n381, MEM_stage_inst_dmem_n380, MEM_stage_inst_dmem_n379, MEM_stage_inst_dmem_n378, MEM_stage_inst_dmem_n377, MEM_stage_inst_dmem_n376, MEM_stage_inst_dmem_n375, MEM_stage_inst_dmem_n374, MEM_stage_inst_dmem_n373, MEM_stage_inst_dmem_n372, MEM_stage_inst_dmem_n371, MEM_stage_inst_dmem_n370, MEM_stage_inst_dmem_n369, MEM_stage_inst_dmem_n368, MEM_stage_inst_dmem_n367, MEM_stage_inst_dmem_n366, MEM_stage_inst_dmem_n365, MEM_stage_inst_dmem_n364, MEM_stage_inst_dmem_n363, MEM_stage_inst_dmem_n362, MEM_stage_inst_dmem_n361, MEM_stage_inst_dmem_n360, MEM_stage_inst_dmem_n359, MEM_stage_inst_dmem_n358, MEM_stage_inst_dmem_n357, MEM_stage_inst_dmem_n356, MEM_stage_inst_dmem_n355, MEM_stage_inst_dmem_n354, MEM_stage_inst_dmem_n353, MEM_stage_inst_dmem_n352, MEM_stage_inst_dmem_n351, MEM_stage_inst_dmem_n350, MEM_stage_inst_dmem_n349, MEM_stage_inst_dmem_n348, MEM_stage_inst_dmem_n347, MEM_stage_inst_dmem_n346, MEM_stage_inst_dmem_n345, MEM_stage_inst_dmem_n344, MEM_stage_inst_dmem_n343, MEM_stage_inst_dmem_n342, MEM_stage_inst_dmem_n341, MEM_stage_inst_dmem_n340, MEM_stage_inst_dmem_n339, MEM_stage_inst_dmem_n338, MEM_stage_inst_dmem_n337, MEM_stage_inst_dmem_n336, MEM_stage_inst_dmem_n335, MEM_stage_inst_dmem_n334, MEM_stage_inst_dmem_n333, MEM_stage_inst_dmem_n332, MEM_stage_inst_dmem_n331, MEM_stage_inst_dmem_n330, MEM_stage_inst_dmem_n329, MEM_stage_inst_dmem_n328, MEM_stage_inst_dmem_n327, MEM_stage_inst_dmem_n326, MEM_stage_inst_dmem_n325, MEM_stage_inst_dmem_n324, MEM_stage_inst_dmem_n323, MEM_stage_inst_dmem_n322, MEM_stage_inst_dmem_n321, MEM_stage_inst_dmem_n320, MEM_stage_inst_dmem_n319, MEM_stage_inst_dmem_n318, MEM_stage_inst_dmem_n317, MEM_stage_inst_dmem_n316, MEM_stage_inst_dmem_n315, MEM_stage_inst_dmem_n314, MEM_stage_inst_dmem_n313, MEM_stage_inst_dmem_n312, MEM_stage_inst_dmem_n311, MEM_stage_inst_dmem_n310, MEM_stage_inst_dmem_n309, MEM_stage_inst_dmem_n308, MEM_stage_inst_dmem_n307, MEM_stage_inst_dmem_n306, MEM_stage_inst_dmem_n305, MEM_stage_inst_dmem_n304, MEM_stage_inst_dmem_n303, MEM_stage_inst_dmem_n302, MEM_stage_inst_dmem_n301, MEM_stage_inst_dmem_n300, MEM_stage_inst_dmem_n299, MEM_stage_inst_dmem_n298, MEM_stage_inst_dmem_n297, MEM_stage_inst_dmem_n296, MEM_stage_inst_dmem_n295, MEM_stage_inst_dmem_n294, MEM_stage_inst_dmem_n293, MEM_stage_inst_dmem_n292, MEM_stage_inst_dmem_n291, MEM_stage_inst_dmem_n290, MEM_stage_inst_dmem_n289, MEM_stage_inst_dmem_n288, MEM_stage_inst_dmem_n287, MEM_stage_inst_dmem_n286, MEM_stage_inst_dmem_n285, MEM_stage_inst_dmem_n284, MEM_stage_inst_dmem_n283, MEM_stage_inst_dmem_n282, MEM_stage_inst_dmem_n281, MEM_stage_inst_dmem_n280, MEM_stage_inst_dmem_n279, MEM_stage_inst_dmem_n278, MEM_stage_inst_dmem_n277, MEM_stage_inst_dmem_n276, MEM_stage_inst_dmem_n275, MEM_stage_inst_dmem_n274, MEM_stage_inst_dmem_n273, MEM_stage_inst_dmem_n272, MEM_stage_inst_dmem_n271, MEM_stage_inst_dmem_n270, MEM_stage_inst_dmem_n269, MEM_stage_inst_dmem_n268, MEM_stage_inst_dmem_n267, MEM_stage_inst_dmem_n266, MEM_stage_inst_dmem_n265, MEM_stage_inst_dmem_n264, MEM_stage_inst_dmem_n263, MEM_stage_inst_dmem_n262, MEM_stage_inst_dmem_n261, MEM_stage_inst_dmem_n260, MEM_stage_inst_dmem_n259, MEM_stage_inst_dmem_n258, MEM_stage_inst_dmem_n257, MEM_stage_inst_dmem_n256, MEM_stage_inst_dmem_n255, MEM_stage_inst_dmem_n254, MEM_stage_inst_dmem_n253, MEM_stage_inst_dmem_n252, MEM_stage_inst_dmem_n251, MEM_stage_inst_dmem_n250, MEM_stage_inst_dmem_n249, MEM_stage_inst_dmem_n248, MEM_stage_inst_dmem_n247, MEM_stage_inst_dmem_n246, MEM_stage_inst_dmem_n245, MEM_stage_inst_dmem_n244, MEM_stage_inst_dmem_n243, MEM_stage_inst_dmem_n242, MEM_stage_inst_dmem_n241, MEM_stage_inst_dmem_n240, MEM_stage_inst_dmem_n239, MEM_stage_inst_dmem_n238, MEM_stage_inst_dmem_n237, MEM_stage_inst_dmem_n236, MEM_stage_inst_dmem_n235, MEM_stage_inst_dmem_n234, MEM_stage_inst_dmem_n233, MEM_stage_inst_dmem_n232, MEM_stage_inst_dmem_n231, MEM_stage_inst_dmem_n230, MEM_stage_inst_dmem_n229, MEM_stage_inst_dmem_n228, MEM_stage_inst_dmem_n227, MEM_stage_inst_dmem_n226, MEM_stage_inst_dmem_n225, MEM_stage_inst_dmem_n224, MEM_stage_inst_dmem_n223, MEM_stage_inst_dmem_n116, MEM_stage_inst_dmem_n115, MEM_stage_inst_dmem_n114, MEM_stage_inst_dmem_n113, MEM_stage_inst_dmem_n112, MEM_stage_inst_dmem_n111, MEM_stage_inst_dmem_n109, MEM_stage_inst_dmem_n105, MEM_stage_inst_dmem_n104, MEM_stage_inst_dmem_n103, MEM_stage_inst_dmem_n102, MEM_stage_inst_dmem_n101, MEM_stage_inst_dmem_n100, MEM_stage_inst_dmem_n96, MEM_stage_inst_dmem_n77, MEM_stage_inst_dmem_n76, MEM_stage_inst_dmem_n75, MEM_stage_inst_dmem_n74, MEM_stage_inst_dmem_n73, MEM_stage_inst_dmem_n72, MEM_stage_inst_dmem_n71, MEM_stage_inst_dmem_n70, MEM_stage_inst_dmem_n69, MEM_stage_inst_dmem_n68, MEM_stage_inst_dmem_n67, MEM_stage_inst_dmem_n66, MEM_stage_inst_dmem_n65, MEM_stage_inst_dmem_n64, MEM_stage_inst_dmem_n63, MEM_stage_inst_dmem_n62, MEM_stage_inst_dmem_n61, MEM_stage_inst_dmem_n60, MEM_stage_inst_dmem_n59, MEM_stage_inst_dmem_n58, MEM_stage_inst_dmem_n57, MEM_stage_inst_dmem_n56, MEM_stage_inst_dmem_n55, MEM_stage_inst_dmem_n54, MEM_stage_inst_dmem_n53, MEM_stage_inst_dmem_n52, MEM_stage_inst_dmem_n51, MEM_stage_inst_dmem_n50, MEM_stage_inst_dmem_n49, MEM_stage_inst_dmem_n48, MEM_stage_inst_dmem_n47, MEM_stage_inst_dmem_n46, MEM_stage_inst_dmem_n45, MEM_stage_inst_dmem_n44, MEM_stage_inst_dmem_n43, MEM_stage_inst_dmem_n42, MEM_stage_inst_dmem_n41, MEM_stage_inst_dmem_n40, MEM_stage_inst_dmem_n39, MEM_stage_inst_dmem_n38, MEM_stage_inst_dmem_n37, MEM_stage_inst_dmem_n36, MEM_stage_inst_dmem_n35, MEM_stage_inst_dmem_n34, MEM_stage_inst_dmem_n33, MEM_stage_inst_dmem_n32, MEM_stage_inst_dmem_n31, MEM_stage_inst_dmem_n30, MEM_stage_inst_dmem_n29, MEM_stage_inst_dmem_n28, MEM_stage_inst_dmem_n27, MEM_stage_inst_dmem_n26, MEM_stage_inst_dmem_n25, MEM_stage_inst_dmem_n24, MEM_stage_inst_dmem_n23, MEM_stage_inst_dmem_n22, MEM_stage_inst_dmem_n21, MEM_stage_inst_dmem_n20, MEM_stage_inst_dmem_n19, MEM_stage_inst_dmem_n18, MEM_stage_inst_dmem_n17, MEM_stage_inst_dmem_n16, MEM_stage_inst_dmem_n15, MEM_stage_inst_dmem_n14, MEM_stage_inst_dmem_n13, MEM_stage_inst_dmem_n12, MEM_stage_inst_dmem_n11, MEM_stage_inst_dmem_n10, MEM_stage_inst_dmem_n9, MEM_stage_inst_dmem_n8, MEM_stage_inst_dmem_n7, MEM_stage_inst_dmem_n6, MEM_stage_inst_dmem_n5, MEM_stage_inst_dmem_n4, MEM_stage_inst_dmem_n3, MEM_stage_inst_dmem_n2, MEM_stage_inst_dmem_n1;

INV_X1 U1873 ( .A(rst), .ZN(n1739) );
BUF_X1 U1874 ( .A(n3521), .Z(n3520) );
INV_X1 U1875 ( .A(n1742), .ZN(n1740) );
INV_X2 U1876 ( .A(n1740), .ZN(n1741) );
BUF_X1 U1877 ( .A(n3521), .Z(n1742) );
BUF_X4 U1878 ( .A(n3521), .Z(n3518) );
INV_X1 U1880 ( .A(rst), .ZN(n3521) );
BUF_X1 U1881 ( .A(n1741), .Z(n3517) );
AND2_X1 U1882 ( .A1(n2516), .A2(n2515), .ZN(n2517) );
OR2_X1 U1883 ( .A1(n2518), .A2(n2517), .ZN(n2577) );
OR2_X1 U1884 ( .A1(ID_pipeline_reg_out_35), .A2(ID_pipeline_reg_out_27), .ZN(n2360) );
AND2_X1 U1885 ( .A1(n2840), .A2(n2839), .ZN(n2841) );
AND2_X1 U1886 ( .A1(n3008), .A2(n3007), .ZN(n3009) );
AND2_X1 U1887 ( .A1(n2577), .A2(n2576), .ZN(n2578) );
AND2_X1 U1888 ( .A1(n2961), .A2(n2960), .ZN(n2962) );
INV_X1 U1889 ( .A(n3104), .ZN(n3037) );
INV_X1 U1890 ( .A(n3026), .ZN(n2998) );
OR2_X1 U1891 ( .A1(n2842), .A2(n2841), .ZN(n2864) );
INV_X1 U1892 ( .A(n2871), .ZN(n3034) );
INV_X1 U1893 ( .A(n3022), .ZN(n2976) );
OR2_X1 U1894 ( .A1(n2904), .A2(n2903), .ZN(n2961) );
OR2_X1 U1895 ( .A1(n2668), .A2(n2667), .ZN(n2711) );
OR2_X1 U1896 ( .A1(n3061), .A2(n3060), .ZN(n3090) );
OR2_X1 U1897 ( .A1(n2866), .A2(n2865), .ZN(n2902) );
INV_X1 U1898 ( .A(n3108), .ZN(n3045) );
OR2_X1 U1899 ( .A1(n3092), .A2(n3091), .ZN(n3096) );
AND2_X1 U1900 ( .A1(n2757), .A2(n2756), .ZN(n2758) );
INV_X1 U1901 ( .A(n2447), .ZN(n2454) );
INV_X1 U1902 ( .A(n3024), .ZN(n2978) );
AND2_X1 U1903 ( .A1(n2711), .A2(n2710), .ZN(n2712) );
INV_X1 U1904 ( .A(n2538), .ZN(n2747) );
INV_X1 U1905 ( .A(n3080), .ZN(n2884) );
INV_X1 U1906 ( .A(n3075), .ZN(n3115) );
INV_X1 U1907 ( .A(n1738), .ZN(n1751) );
OR2_X1 U1908 ( .A1(n2759), .A2(n2758), .ZN(n2778) );
OR2_X1 U1909 ( .A1(n2713), .A2(n2712), .ZN(n2757) );
OR2_X1 U1910 ( .A1(n2631), .A2(n2630), .ZN(n2666) );
INV_X1 U1911 ( .A(n3119), .ZN(n2936) );
INV_X1 U1912 ( .A(n2874), .ZN(n3042) );
INV_X1 U1913 ( .A(n1778), .ZN(n1763) );
AND2_X1 U1914 ( .A1(n1798), .A2(n1797), .ZN(n1800) );
AND2_X1 U1915 ( .A1(n2079), .A2(n2078), .ZN(n2056) );
INV_X1 U1916 ( .A(n2595), .ZN(n2598) );
AND2_X1 U1917 ( .A1(n2350), .A2(n2349), .ZN(n2351) );
OR2_X1 U1918 ( .A1(n2061), .A2(n2060), .ZN(n2064) );
INV_X1 U1919 ( .A(n2609), .ZN(n2772) );
INV_X1 U1920 ( .A(n3078), .ZN(n2746) );
INV_X1 U1921 ( .A(n2325), .ZN(n2326) );
INV_X1 U1922 ( .A(n3446), .ZN(n3447) );
INV_X1 U1923 ( .A(n2357), .ZN(n2331) );
INV_X1 U1924 ( .A(n3167), .ZN(n3140) );
INV_X1 U1925 ( .A(n3144), .ZN(n2118) );
INV_X1 U1926 ( .A(n2680), .ZN(n2600) );
INV_X1 U1927 ( .A(n2344), .ZN(n2353) );
AND2_X1 U1928 ( .A1(n1822), .A2(n1821), .ZN(n3163) );
BUF_X1 U1929 ( .A(n1739), .Z(n3519) );
AND2_X1 U1930 ( .A1(MEM_stage_inst_mem_read_data_15), .A2(n3518), .ZN(MEM_stage_inst_N23) );
AND2_X1 U1931 ( .A1(MEM_stage_inst_mem_read_data_0), .A2(n3518), .ZN(MEM_stage_inst_N8) );
AND2_X1 U1932 ( .A1(EX_pipeline_reg_out_0), .A2(n3518), .ZN(MEM_stage_inst_N3) );
AND2_X1 U1933 ( .A1(EX_pipeline_reg_out_37), .A2(n3518), .ZN(MEM_stage_inst_N39) );
AND2_X1 U1934 ( .A1(EX_pipeline_reg_out_36), .A2(n3518), .ZN(MEM_stage_inst_N38) );
AND2_X1 U1935 ( .A1(ID_pipeline_reg_out_4), .A2(n3518), .ZN(EX_stage_inst_N7) );
AND2_X1 U1936 ( .A1(EX_pipeline_reg_out_4), .A2(n3518), .ZN(MEM_stage_inst_N7) );
AND2_X1 U1937 ( .A1(EX_pipeline_reg_out_30), .A2(n3518), .ZN(MEM_stage_inst_N32) );
AND2_X1 U1938 ( .A1(EX_pipeline_reg_out_32), .A2(n3518), .ZN(MEM_stage_inst_N34) );
AND2_X1 U1939 ( .A1(EX_pipeline_reg_out_34), .A2(n3518), .ZN(MEM_stage_inst_N36) );
AND2_X1 U1940 ( .A1(EX_pipeline_reg_out_33), .A2(n3521), .ZN(MEM_stage_inst_N35) );
AND2_X1 U1941 ( .A1(EX_pipeline_reg_out_35), .A2(n3518), .ZN(MEM_stage_inst_N37) );
AND2_X1 U1942 ( .A1(EX_pipeline_reg_out_31), .A2(n3521), .ZN(MEM_stage_inst_N33) );
AND2_X1 U1943 ( .A1(ID_pipeline_reg_out_7), .A2(n3518), .ZN(EX_stage_inst_N10) );
AND2_X1 U1944 ( .A1(n3518), .A2(mem_op_dest_2), .ZN(MEM_stage_inst_N6) );
NAND2_X1 U1945 ( .A1(ID_stage_inst_instruction_reg_15), .A2(ID_stage_inst_instruction_reg_12), .ZN(n1746) );
NAND2_X1 U1946 ( .A1(ID_stage_inst_instruction_reg_13), .A2(n3510), .ZN(n1745) );
NOR2_X1 U1947 ( .A1(n1746), .A2(n1745), .ZN(n1738) );
NAND2_X1 U1948 ( .A1(branch_offset_imm_5), .A2(n1751), .ZN(n1748) );
NAND2_X1 U1949 ( .A1(n1738), .A2(ID_stage_inst_instruction_reg_11), .ZN(n1747) );
NAND2_X1 U1950 ( .A1(n1748), .A2(n1747), .ZN(n1778) );
NAND2_X1 U1951 ( .A1(branch_offset_imm_3), .A2(n1751), .ZN(n1750) );
NAND2_X1 U1952 ( .A1(n1738), .A2(ID_stage_inst_instruction_reg_9), .ZN(n1749) );
NAND2_X1 U1953 ( .A1(n1750), .A2(n1749), .ZN(n1781) );
NAND2_X1 U1954 ( .A1(branch_offset_imm_4), .A2(n1751), .ZN(n1753) );
NAND2_X1 U1955 ( .A1(n1738), .A2(ID_stage_inst_instruction_reg_10), .ZN(n1752) );
NAND2_X1 U1956 ( .A1(n1753), .A2(n1752), .ZN(n1777) );
INV_X1 U1957 ( .A(n1777), .ZN(n1764) );
OR2_X1 U1958 ( .A1(n1781), .A2(n1764), .ZN(n1758) );
NOR2_X2 U1959 ( .A1(n1778), .A2(n1758), .ZN(n2306) );
NAND2_X1 U1960 ( .A1(register_file_inst_reg_array_18), .A2(n2306), .ZN(n1755) );
NAND2_X1 U1961 ( .A1(n1778), .A2(n1781), .ZN(n1757) );
NOR2_X2 U1962 ( .A1(n1764), .A2(n1757), .ZN(n2307) );
NAND2_X1 U1963 ( .A1(register_file_inst_reg_array_98), .A2(n2307), .ZN(n1754) );
NAND2_X1 U1964 ( .A1(n1755), .A2(n1754), .ZN(n1768) );
NOR2_X1 U1965 ( .A1(n1781), .A2(n1777), .ZN(n1756) );
NAND2_X1 U1966 ( .A1(n1756), .A2(n1778), .ZN(n2310) );
NOR2_X1 U1967 ( .A1(n2310), .A2(n3494), .ZN(n1762) );
NOR2_X2 U1968 ( .A1(n1777), .A2(n1757), .ZN(n2311) );
NAND2_X1 U1969 ( .A1(register_file_inst_reg_array_66), .A2(n2311), .ZN(n1760) );
NOR2_X2 U1970 ( .A1(n1763), .A2(n1758), .ZN(n2312) );
NAND2_X1 U1971 ( .A1(register_file_inst_reg_array_82), .A2(n2312), .ZN(n1759) );
NAND2_X1 U1972 ( .A1(n1760), .A2(n1759), .ZN(n1761) );
NOR2_X1 U1973 ( .A1(n1762), .A2(n1761), .ZN(n1766) );
NAND2_X1 U1974 ( .A1(n1763), .A2(n1781), .ZN(n1769) );
NOR2_X2 U1975 ( .A1(n1764), .A2(n1769), .ZN(n2317) );
NAND2_X1 U1976 ( .A1(register_file_inst_reg_array_34), .A2(n2317), .ZN(n1765) );
NAND2_X1 U1977 ( .A1(n1766), .A2(n1765), .ZN(n1767) );
NOR2_X1 U1978 ( .A1(n1768), .A2(n1767), .ZN(n1771) );
NOR2_X2 U1979 ( .A1(n1777), .A2(n1769), .ZN(n2322) );
NAND2_X1 U1980 ( .A1(n2322), .A2(register_file_inst_reg_array_2), .ZN(n1770) );
NAND2_X1 U1981 ( .A1(n1771), .A2(n1770), .ZN(reg_read_data_2_2) );
NAND2_X1 U1982 ( .A1(ID_stage_inst_instruction_reg_15), .A2(n3487), .ZN(n1774) );
NOR2_X1 U1983 ( .A1(ID_stage_inst_instruction_reg_13), .A2(n1774), .ZN(n2030) );
XOR2_X1 U1984 ( .A(ID_stage_inst_instruction_reg_14), .B(n2030), .Z(n1773) );
NOR2_X1 U1985 ( .A1(ID_stage_inst_instruction_reg_15), .A2(n3487), .ZN(n1772) );
NOR2_X1 U1986 ( .A1(n1773), .A2(n1772), .ZN(n1776) );
NAND2_X1 U1987 ( .A1(ID_stage_inst_instruction_reg_13), .A2(n1774), .ZN(n1775) );
NAND2_X1 U1988 ( .A1(n1776), .A2(n1775), .ZN(n1782) );
NAND2_X1 U1989 ( .A1(n1782), .A2(n1777), .ZN(n1797) );
XOR2_X1 U1990 ( .A(ex_op_dest_1), .B(n1797), .Z(n1780) );
NAND2_X1 U1991 ( .A1(n1782), .A2(n1778), .ZN(n1798) );
XOR2_X1 U1992 ( .A(ex_op_dest_2), .B(n1798), .Z(n1779) );
NAND2_X1 U1993 ( .A1(n1780), .A2(n1779), .ZN(n1784) );
NAND2_X1 U1994 ( .A1(n1782), .A2(n1781), .ZN(n1799) );
XNOR2_X1 U1995 ( .A(n1799), .B(ex_op_dest_0), .ZN(n1783) );
NOR2_X1 U1996 ( .A1(n1784), .A2(n1783), .ZN(n1790) );
XNOR2_X1 U1997 ( .A(mem_op_dest_2), .B(n1798), .ZN(n1788) );
XOR2_X1 U1998 ( .A(mem_op_dest_1), .B(n1797), .Z(n1786) );
XOR2_X1 U1999 ( .A(mem_op_dest_0), .B(n1799), .Z(n1785) );
NAND2_X1 U2000 ( .A1(n1786), .A2(n1785), .ZN(n1787) );
NOR2_X1 U2001 ( .A1(n1788), .A2(n1787), .ZN(n1789) );
NOR2_X1 U2002 ( .A1(n1790), .A2(n1789), .ZN(n1796) );
XNOR2_X1 U2003 ( .A(reg_write_dest_0), .B(n1799), .ZN(n1792) );
XOR2_X1 U2004 ( .A(n3484), .B(n1797), .Z(n1791) );
NOR2_X1 U2005 ( .A1(n1792), .A2(n1791), .ZN(n1794) );
XNOR2_X1 U2006 ( .A(n3475), .B(n1798), .ZN(n1793) );
NAND2_X1 U2007 ( .A1(n1794), .A2(n1793), .ZN(n1795) );
NAND2_X1 U2008 ( .A1(n1796), .A2(n1795), .ZN(n1802) );
NAND2_X1 U2009 ( .A1(n1800), .A2(n1799), .ZN(n1801) );
NAND2_X1 U2010 ( .A1(n1802), .A2(n1801), .ZN(n1822) );
XOR2_X1 U2011 ( .A(n3480), .B(reg_write_dest_1), .Z(n1804) );
XOR2_X1 U2012 ( .A(n3479), .B(reg_write_dest_2), .Z(n1803) );
NAND2_X1 U2013 ( .A1(n1804), .A2(n1803), .ZN(n1806) );
XOR2_X1 U2014 ( .A(reg_read_addr_1_0), .B(reg_write_dest_0), .Z(n1805) );
NOR2_X1 U2015 ( .A1(n1806), .A2(n1805), .ZN(n1812) );
XOR2_X1 U2016 ( .A(n3480), .B(ex_op_dest_1), .Z(n1808) );
XOR2_X1 U2017 ( .A(n3479), .B(ex_op_dest_2), .Z(n1807) );
NAND2_X1 U2018 ( .A1(n1808), .A2(n1807), .ZN(n1810) );
XOR2_X1 U2019 ( .A(reg_read_addr_1_0), .B(ex_op_dest_0), .Z(n1809) );
NOR2_X1 U2020 ( .A1(n1810), .A2(n1809), .ZN(n1811) );
NOR2_X1 U2021 ( .A1(n1812), .A2(n1811), .ZN(n1818) );
XNOR2_X1 U2022 ( .A(n3480), .B(mem_op_dest_1), .ZN(n1814) );
XNOR2_X1 U2023 ( .A(n3479), .B(mem_op_dest_2), .ZN(n1813) );
NOR2_X1 U2024 ( .A1(n1814), .A2(n1813), .ZN(n1816) );
XNOR2_X1 U2025 ( .A(mem_op_dest_0), .B(reg_read_addr_1_0), .ZN(n1815) );
NAND2_X1 U2026 ( .A1(n1816), .A2(n1815), .ZN(n1817) );
NAND2_X1 U2027 ( .A1(n1818), .A2(n1817), .ZN(n1820) );
NOR2_X1 U2028 ( .A1(reg_read_addr_1_0), .A2(reg_read_addr_1_2), .ZN(n1825) );
NAND2_X1 U2029 ( .A1(n3480), .A2(n1825), .ZN(n1819) );
NAND2_X1 U2030 ( .A1(n1820), .A2(n1819), .ZN(n1821) );
NAND2_X1 U2031 ( .A1(ID_stage_inst_instruction_reg_12), .A2(n3163), .ZN(n2350) );
NAND2_X1 U2032 ( .A1(ID_stage_inst_instruction_reg_13), .A2(n3163), .ZN(n2346) );
NAND2_X1 U2033 ( .A1(n2350), .A2(n2346), .ZN(n2333) );
INV_X1 U2034 ( .A(n2333), .ZN(n1823) );
NAND2_X1 U2035 ( .A1(ID_stage_inst_instruction_reg_14), .A2(n3163), .ZN(n2344) );
NOR2_X1 U2036 ( .A1(n1823), .A2(n2344), .ZN(n2341) );
NAND2_X1 U2037 ( .A1(ID_stage_inst_instruction_reg_15), .A2(n3163), .ZN(n2349) );
INV_X1 U2038 ( .A(n2349), .ZN(n2336) );
NAND2_X1 U2039 ( .A1(n2336), .A2(n3518), .ZN(n2345) );
NOR2_X1 U2040 ( .A1(n2341), .A2(n2345), .ZN(n1824) );
NAND2_X1 U2041 ( .A1(n1823), .A2(n2344), .ZN(n2329) );
NAND2_X1 U2042 ( .A1(n1824), .A2(n2329), .ZN(n2325) );
AND2_X1 U2043 ( .A1(reg_read_data_2_2), .A2(n2325), .ZN(ID_stage_inst_ex_alu_src2_2) );
AND2_X1 U2044 ( .A1(n3518), .A2(mem_op_dest_0), .ZN(MEM_stage_inst_N4) );
AND2_X1 U2045 ( .A1(n3518), .A2(ex_op_dest_1), .ZN(EX_stage_inst_N5) );
AND2_X1 U2046 ( .A1(n3518), .A2(mem_op_dest_1), .ZN(MEM_stage_inst_N5) );
AND2_X1 U2047 ( .A1(n3518), .A2(ex_op_dest_2), .ZN(EX_stage_inst_N6) );
AND2_X1 U2048 ( .A1(ID_pipeline_reg_out_0), .A2(n3518), .ZN(EX_stage_inst_N3) );
AND2_X1 U2049 ( .A1(ID_pipeline_reg_out_21), .A2(n3518), .ZN(EX_stage_inst_N24) );
AND2_X1 U2050 ( .A1(ID_pipeline_reg_out_20), .A2(n3518), .ZN(EX_stage_inst_N23) );
AND2_X1 U2051 ( .A1(ID_pipeline_reg_out_15), .A2(n3518), .ZN(EX_stage_inst_N18) );
AND2_X1 U2052 ( .A1(ID_pipeline_reg_out_19), .A2(n3518), .ZN(EX_stage_inst_N22) );
AND2_X1 U2053 ( .A1(ID_pipeline_reg_out_9), .A2(n3518), .ZN(EX_stage_inst_N12) );
AND2_X1 U2054 ( .A1(ID_pipeline_reg_out_16), .A2(n3518), .ZN(EX_stage_inst_N19) );
AND2_X1 U2055 ( .A1(ID_pipeline_reg_out_18), .A2(n3518), .ZN(EX_stage_inst_N21) );
AND2_X1 U2056 ( .A1(n3519), .A2(ex_op_dest_0), .ZN(EX_stage_inst_N4) );
AND2_X1 U2057 ( .A1(ID_pipeline_reg_out_8), .A2(n3518), .ZN(EX_stage_inst_N11) );
AND2_X1 U2058 ( .A1(ID_pipeline_reg_out_10), .A2(n3518), .ZN(EX_stage_inst_N13) );
AND2_X1 U2059 ( .A1(ID_pipeline_reg_out_12), .A2(n3518), .ZN(EX_stage_inst_N15) );
AND2_X1 U2060 ( .A1(MEM_stage_inst_mem_read_data_2), .A2(n3521), .ZN(MEM_stage_inst_N10) );
AND2_X1 U2061 ( .A1(MEM_stage_inst_mem_read_data_4), .A2(n3521), .ZN(MEM_stage_inst_N12) );
AND2_X1 U2062 ( .A1(MEM_stage_inst_mem_read_data_10), .A2(n3521), .ZN(MEM_stage_inst_N18) );
AND2_X1 U2063 ( .A1(MEM_stage_inst_mem_read_data_13), .A2(n3521), .ZN(MEM_stage_inst_N21) );
AND2_X1 U2064 ( .A1(MEM_stage_inst_mem_read_data_1), .A2(n3518), .ZN(MEM_stage_inst_N9) );
AND2_X1 U2065 ( .A1(MEM_stage_inst_mem_read_data_3), .A2(n3518), .ZN(MEM_stage_inst_N11) );
AND2_X1 U2066 ( .A1(MEM_stage_inst_mem_read_data_5), .A2(n3518), .ZN(MEM_stage_inst_N13) );
AND2_X1 U2067 ( .A1(MEM_stage_inst_mem_read_data_6), .A2(n3518), .ZN(MEM_stage_inst_N14) );
AND2_X1 U2068 ( .A1(MEM_stage_inst_mem_read_data_7), .A2(n3518), .ZN(MEM_stage_inst_N15) );
AND2_X1 U2069 ( .A1(MEM_stage_inst_mem_read_data_8), .A2(n3518), .ZN(MEM_stage_inst_N16) );
AND2_X1 U2070 ( .A1(MEM_stage_inst_mem_read_data_9), .A2(n3518), .ZN(MEM_stage_inst_N17) );
AND2_X1 U2071 ( .A1(MEM_stage_inst_mem_read_data_11), .A2(n3518), .ZN(MEM_stage_inst_N19) );
AND2_X1 U2072 ( .A1(MEM_stage_inst_mem_read_data_12), .A2(n3518), .ZN(MEM_stage_inst_N20) );
AND2_X1 U2073 ( .A1(MEM_stage_inst_mem_read_data_14), .A2(n3518), .ZN(MEM_stage_inst_N22) );
INV_X1 U2074 ( .A(n3163), .ZN(n3176) );
NOR2_X1 U2075 ( .A1(n3176), .A2(n3515), .ZN(ID_stage_inst_ir_dest_with_bubble_1) );
AND2_X1 U2076 ( .A1(ID_stage_inst_instruction_reg_9), .A2(n3163), .ZN(ID_stage_inst_ir_dest_with_bubble_0) );
AND2_X1 U2077 ( .A1(ID_stage_inst_instruction_reg_11), .A2(n3163), .ZN(ID_stage_inst_ir_dest_with_bubble_2) );
AND2_X1 U2078 ( .A1(reg_read_addr_1_1), .A2(n1825), .ZN(n2009) );
NAND2_X1 U2079 ( .A1(register_file_inst_reg_array_31), .A2(n2009), .ZN(n1840) );
NAND2_X1 U2080 ( .A1(reg_read_addr_1_0), .A2(reg_read_addr_1_1), .ZN(n1826) );
NOR2_X2 U2081 ( .A1(n3479), .A2(n1826), .ZN(n2010) );
NAND2_X1 U2082 ( .A1(n2010), .A2(register_file_inst_reg_array_111), .ZN(n1828) );
NOR2_X2 U2083 ( .A1(reg_read_addr_1_2), .A2(n1826), .ZN(n2011) );
NAND2_X1 U2084 ( .A1(n2011), .A2(register_file_inst_reg_array_47), .ZN(n1827) );
NAND2_X1 U2085 ( .A1(n1828), .A2(n1827), .ZN(n1838) );
NOR2_X1 U2086 ( .A1(n3479), .A2(reg_read_addr_1_0), .ZN(n1829) );
NAND2_X1 U2087 ( .A1(n1829), .A2(n3480), .ZN(n2014) );
NOR2_X1 U2088 ( .A1(n3492), .A2(n2014), .ZN(n1833) );
NAND2_X1 U2089 ( .A1(reg_read_addr_1_0), .A2(n3480), .ZN(n1834) );
NOR2_X2 U2090 ( .A1(n3479), .A2(n1834), .ZN(n2015) );
NAND2_X1 U2091 ( .A1(n2015), .A2(register_file_inst_reg_array_79), .ZN(n1831) );
AND2_X1 U2092 ( .A1(reg_read_addr_1_1), .A2(n1829), .ZN(n2016) );
NAND2_X1 U2093 ( .A1(n2016), .A2(register_file_inst_reg_array_95), .ZN(n1830) );
NAND2_X1 U2094 ( .A1(n1831), .A2(n1830), .ZN(n1832) );
NOR2_X1 U2095 ( .A1(n1833), .A2(n1832), .ZN(n1836) );
NOR2_X2 U2096 ( .A1(reg_read_addr_1_2), .A2(n1834), .ZN(n2021) );
NAND2_X1 U2097 ( .A1(n2021), .A2(register_file_inst_reg_array_15), .ZN(n1835) );
NAND2_X1 U2098 ( .A1(n1836), .A2(n1835), .ZN(n1837) );
NOR2_X1 U2099 ( .A1(n1838), .A2(n1837), .ZN(n1839) );
NAND2_X1 U2100 ( .A1(n1840), .A2(n1839), .ZN(reg_read_data_1_15) );
NAND2_X1 U2101 ( .A1(register_file_inst_reg_array_25), .A2(n2009), .ZN(n1852) );
NAND2_X1 U2102 ( .A1(n2010), .A2(register_file_inst_reg_array_105), .ZN(n1842) );
NAND2_X1 U2103 ( .A1(n2011), .A2(register_file_inst_reg_array_41), .ZN(n1841) );
NAND2_X1 U2104 ( .A1(n1842), .A2(n1841), .ZN(n1850) );
NOR2_X1 U2105 ( .A1(n3493), .A2(n2014), .ZN(n1846) );
NAND2_X1 U2106 ( .A1(n2015), .A2(register_file_inst_reg_array_73), .ZN(n1844) );
NAND2_X1 U2107 ( .A1(n2016), .A2(register_file_inst_reg_array_89), .ZN(n1843) );
NAND2_X1 U2108 ( .A1(n1844), .A2(n1843), .ZN(n1845) );
NOR2_X1 U2109 ( .A1(n1846), .A2(n1845), .ZN(n1848) );
NAND2_X1 U2110 ( .A1(n2021), .A2(register_file_inst_reg_array_9), .ZN(n1847) );
NAND2_X1 U2111 ( .A1(n1848), .A2(n1847), .ZN(n1849) );
NOR2_X1 U2112 ( .A1(n1850), .A2(n1849), .ZN(n1851) );
NAND2_X1 U2113 ( .A1(n1852), .A2(n1851), .ZN(reg_read_data_1_9) );
NAND2_X1 U2114 ( .A1(register_file_inst_reg_array_18), .A2(n2009), .ZN(n1864) );
NAND2_X1 U2115 ( .A1(n2010), .A2(register_file_inst_reg_array_98), .ZN(n1854) );
NAND2_X1 U2116 ( .A1(n2011), .A2(register_file_inst_reg_array_34), .ZN(n1853) );
NAND2_X1 U2117 ( .A1(n1854), .A2(n1853), .ZN(n1862) );
NOR2_X1 U2118 ( .A1(n3494), .A2(n2014), .ZN(n1858) );
NAND2_X1 U2119 ( .A1(n2015), .A2(register_file_inst_reg_array_66), .ZN(n1856) );
NAND2_X1 U2120 ( .A1(n2016), .A2(register_file_inst_reg_array_82), .ZN(n1855) );
NAND2_X1 U2121 ( .A1(n1856), .A2(n1855), .ZN(n1857) );
NOR2_X1 U2122 ( .A1(n1858), .A2(n1857), .ZN(n1860) );
NAND2_X1 U2123 ( .A1(n2021), .A2(register_file_inst_reg_array_2), .ZN(n1859) );
NAND2_X1 U2124 ( .A1(n1860), .A2(n1859), .ZN(n1861) );
NOR2_X1 U2125 ( .A1(n1862), .A2(n1861), .ZN(n1863) );
NAND2_X1 U2126 ( .A1(n1864), .A2(n1863), .ZN(reg_read_data_1_2) );
NAND2_X1 U2127 ( .A1(register_file_inst_reg_array_16), .A2(n2009), .ZN(n1876) );
NAND2_X1 U2128 ( .A1(n2010), .A2(register_file_inst_reg_array_96), .ZN(n1866) );
NAND2_X1 U2129 ( .A1(n2011), .A2(register_file_inst_reg_array_32), .ZN(n1865) );
NAND2_X1 U2130 ( .A1(n1866), .A2(n1865), .ZN(n1874) );
NOR2_X1 U2131 ( .A1(n3491), .A2(n2014), .ZN(n1870) );
NAND2_X1 U2132 ( .A1(n2015), .A2(register_file_inst_reg_array_64), .ZN(n1868) );
NAND2_X1 U2133 ( .A1(n2016), .A2(register_file_inst_reg_array_80), .ZN(n1867) );
NAND2_X1 U2134 ( .A1(n1868), .A2(n1867), .ZN(n1869) );
NOR2_X1 U2135 ( .A1(n1870), .A2(n1869), .ZN(n1872) );
NAND2_X1 U2136 ( .A1(n2021), .A2(register_file_inst_reg_array_0), .ZN(n1871) );
NAND2_X1 U2137 ( .A1(n1872), .A2(n1871), .ZN(n1873) );
NOR2_X1 U2138 ( .A1(n1874), .A2(n1873), .ZN(n1875) );
NAND2_X1 U2139 ( .A1(n1876), .A2(n1875), .ZN(reg_read_data_1_0) );
NAND2_X1 U2140 ( .A1(register_file_inst_reg_array_28), .A2(n2009), .ZN(n1888) );
NAND2_X1 U2141 ( .A1(n2010), .A2(register_file_inst_reg_array_108), .ZN(n1878) );
NAND2_X1 U2142 ( .A1(n2011), .A2(register_file_inst_reg_array_44), .ZN(n1877) );
NAND2_X1 U2143 ( .A1(n1878), .A2(n1877), .ZN(n1886) );
NOR2_X1 U2144 ( .A1(n3495), .A2(n2014), .ZN(n1882) );
NAND2_X1 U2145 ( .A1(n2015), .A2(register_file_inst_reg_array_76), .ZN(n1880) );
NAND2_X1 U2146 ( .A1(n2016), .A2(register_file_inst_reg_array_92), .ZN(n1879) );
NAND2_X1 U2147 ( .A1(n1880), .A2(n1879), .ZN(n1881) );
NOR2_X1 U2148 ( .A1(n1882), .A2(n1881), .ZN(n1884) );
NAND2_X1 U2149 ( .A1(n2021), .A2(register_file_inst_reg_array_12), .ZN(n1883) );
NAND2_X1 U2150 ( .A1(n1884), .A2(n1883), .ZN(n1885) );
NOR2_X1 U2151 ( .A1(n1886), .A2(n1885), .ZN(n1887) );
NAND2_X1 U2152 ( .A1(n1888), .A2(n1887), .ZN(reg_read_data_1_12) );
NAND2_X1 U2153 ( .A1(register_file_inst_reg_array_20), .A2(n2009), .ZN(n1900) );
NAND2_X1 U2154 ( .A1(n2010), .A2(register_file_inst_reg_array_100), .ZN(n1890) );
NAND2_X1 U2155 ( .A1(n2011), .A2(register_file_inst_reg_array_36), .ZN(n1889) );
NAND2_X1 U2156 ( .A1(n1890), .A2(n1889), .ZN(n1898) );
NOR2_X1 U2157 ( .A1(n3496), .A2(n2014), .ZN(n1894) );
NAND2_X1 U2158 ( .A1(n2015), .A2(register_file_inst_reg_array_68), .ZN(n1892) );
NAND2_X1 U2159 ( .A1(n2016), .A2(register_file_inst_reg_array_84), .ZN(n1891) );
NAND2_X1 U2160 ( .A1(n1892), .A2(n1891), .ZN(n1893) );
NOR2_X1 U2161 ( .A1(n1894), .A2(n1893), .ZN(n1896) );
NAND2_X1 U2162 ( .A1(n2021), .A2(register_file_inst_reg_array_4), .ZN(n1895) );
NAND2_X1 U2163 ( .A1(n1896), .A2(n1895), .ZN(n1897) );
NOR2_X1 U2164 ( .A1(n1898), .A2(n1897), .ZN(n1899) );
NAND2_X1 U2165 ( .A1(n1900), .A2(n1899), .ZN(reg_read_data_1_4) );
NAND2_X1 U2166 ( .A1(register_file_inst_reg_array_21), .A2(n2009), .ZN(n1912) );
NAND2_X1 U2167 ( .A1(n2010), .A2(register_file_inst_reg_array_101), .ZN(n1902) );
NAND2_X1 U2168 ( .A1(n2011), .A2(register_file_inst_reg_array_37), .ZN(n1901) );
NAND2_X1 U2169 ( .A1(n1902), .A2(n1901), .ZN(n1910) );
NOR2_X1 U2170 ( .A1(n3497), .A2(n2014), .ZN(n1906) );
NAND2_X1 U2171 ( .A1(n2015), .A2(register_file_inst_reg_array_69), .ZN(n1904) );
NAND2_X1 U2172 ( .A1(n2016), .A2(register_file_inst_reg_array_85), .ZN(n1903) );
NAND2_X1 U2173 ( .A1(n1904), .A2(n1903), .ZN(n1905) );
NOR2_X1 U2174 ( .A1(n1906), .A2(n1905), .ZN(n1908) );
NAND2_X1 U2175 ( .A1(n2021), .A2(register_file_inst_reg_array_5), .ZN(n1907) );
NAND2_X1 U2176 ( .A1(n1908), .A2(n1907), .ZN(n1909) );
NOR2_X1 U2177 ( .A1(n1910), .A2(n1909), .ZN(n1911) );
NAND2_X1 U2178 ( .A1(n1912), .A2(n1911), .ZN(reg_read_data_1_5) );
NAND2_X1 U2179 ( .A1(register_file_inst_reg_array_27), .A2(n2009), .ZN(n1924) );
NAND2_X1 U2180 ( .A1(n2010), .A2(register_file_inst_reg_array_107), .ZN(n1914) );
NAND2_X1 U2181 ( .A1(n2011), .A2(register_file_inst_reg_array_43), .ZN(n1913) );
NAND2_X1 U2182 ( .A1(n1914), .A2(n1913), .ZN(n1922) );
NOR2_X1 U2183 ( .A1(n3498), .A2(n2014), .ZN(n1918) );
NAND2_X1 U2184 ( .A1(n2015), .A2(register_file_inst_reg_array_75), .ZN(n1916) );
NAND2_X1 U2185 ( .A1(n2016), .A2(register_file_inst_reg_array_91), .ZN(n1915) );
NAND2_X1 U2186 ( .A1(n1916), .A2(n1915), .ZN(n1917) );
NOR2_X1 U2187 ( .A1(n1918), .A2(n1917), .ZN(n1920) );
NAND2_X1 U2188 ( .A1(n2021), .A2(register_file_inst_reg_array_11), .ZN(n1919) );
NAND2_X1 U2189 ( .A1(n1920), .A2(n1919), .ZN(n1921) );
NOR2_X1 U2190 ( .A1(n1922), .A2(n1921), .ZN(n1923) );
NAND2_X1 U2191 ( .A1(n1924), .A2(n1923), .ZN(reg_read_data_1_11) );
NAND2_X1 U2192 ( .A1(register_file_inst_reg_array_17), .A2(n2009), .ZN(n1936) );
NAND2_X1 U2193 ( .A1(n2010), .A2(register_file_inst_reg_array_97), .ZN(n1926) );
NAND2_X1 U2194 ( .A1(n2011), .A2(register_file_inst_reg_array_33), .ZN(n1925) );
NAND2_X1 U2195 ( .A1(n1926), .A2(n1925), .ZN(n1934) );
NOR2_X1 U2196 ( .A1(n3499), .A2(n2014), .ZN(n1930) );
NAND2_X1 U2197 ( .A1(n2015), .A2(register_file_inst_reg_array_65), .ZN(n1928) );
NAND2_X1 U2198 ( .A1(n2016), .A2(register_file_inst_reg_array_81), .ZN(n1927) );
NAND2_X1 U2199 ( .A1(n1928), .A2(n1927), .ZN(n1929) );
NOR2_X1 U2200 ( .A1(n1930), .A2(n1929), .ZN(n1932) );
NAND2_X1 U2201 ( .A1(n2021), .A2(register_file_inst_reg_array_1), .ZN(n1931) );
NAND2_X1 U2202 ( .A1(n1932), .A2(n1931), .ZN(n1933) );
NOR2_X1 U2203 ( .A1(n1934), .A2(n1933), .ZN(n1935) );
NAND2_X1 U2204 ( .A1(n1936), .A2(n1935), .ZN(reg_read_data_1_1) );
NAND2_X1 U2205 ( .A1(register_file_inst_reg_array_24), .A2(n2009), .ZN(n1948) );
NAND2_X1 U2206 ( .A1(n2010), .A2(register_file_inst_reg_array_104), .ZN(n1938) );
NAND2_X1 U2207 ( .A1(n2011), .A2(register_file_inst_reg_array_40), .ZN(n1937) );
NAND2_X1 U2208 ( .A1(n1938), .A2(n1937), .ZN(n1946) );
NOR2_X1 U2209 ( .A1(n3500), .A2(n2014), .ZN(n1942) );
NAND2_X1 U2210 ( .A1(n2015), .A2(register_file_inst_reg_array_72), .ZN(n1940) );
NAND2_X1 U2211 ( .A1(n2016), .A2(register_file_inst_reg_array_88), .ZN(n1939) );
NAND2_X1 U2212 ( .A1(n1940), .A2(n1939), .ZN(n1941) );
NOR2_X1 U2213 ( .A1(n1942), .A2(n1941), .ZN(n1944) );
NAND2_X1 U2214 ( .A1(n2021), .A2(register_file_inst_reg_array_8), .ZN(n1943) );
NAND2_X1 U2215 ( .A1(n1944), .A2(n1943), .ZN(n1945) );
NOR2_X1 U2216 ( .A1(n1946), .A2(n1945), .ZN(n1947) );
NAND2_X1 U2217 ( .A1(n1948), .A2(n1947), .ZN(reg_read_data_1_8) );
NAND2_X1 U2218 ( .A1(register_file_inst_reg_array_30), .A2(n2009), .ZN(n1960) );
NAND2_X1 U2219 ( .A1(n2010), .A2(register_file_inst_reg_array_110), .ZN(n1950) );
NAND2_X1 U2220 ( .A1(n2011), .A2(register_file_inst_reg_array_46), .ZN(n1949) );
NAND2_X1 U2221 ( .A1(n1950), .A2(n1949), .ZN(n1958) );
NOR2_X1 U2222 ( .A1(n3501), .A2(n2014), .ZN(n1954) );
NAND2_X1 U2223 ( .A1(n2015), .A2(register_file_inst_reg_array_78), .ZN(n1952) );
NAND2_X1 U2224 ( .A1(n2016), .A2(register_file_inst_reg_array_94), .ZN(n1951) );
NAND2_X1 U2225 ( .A1(n1952), .A2(n1951), .ZN(n1953) );
NOR2_X1 U2226 ( .A1(n1954), .A2(n1953), .ZN(n1956) );
NAND2_X1 U2227 ( .A1(n2021), .A2(register_file_inst_reg_array_14), .ZN(n1955) );
NAND2_X1 U2228 ( .A1(n1956), .A2(n1955), .ZN(n1957) );
NOR2_X1 U2229 ( .A1(n1958), .A2(n1957), .ZN(n1959) );
NAND2_X1 U2230 ( .A1(n1960), .A2(n1959), .ZN(reg_read_data_1_14) );
NAND2_X1 U2231 ( .A1(register_file_inst_reg_array_29), .A2(n2009), .ZN(n1972) );
NAND2_X1 U2232 ( .A1(n2010), .A2(register_file_inst_reg_array_109), .ZN(n1962) );
NAND2_X1 U2233 ( .A1(n2011), .A2(register_file_inst_reg_array_45), .ZN(n1961) );
NAND2_X1 U2234 ( .A1(n1962), .A2(n1961), .ZN(n1970) );
NOR2_X1 U2235 ( .A1(n3502), .A2(n2014), .ZN(n1966) );
NAND2_X1 U2236 ( .A1(n2015), .A2(register_file_inst_reg_array_77), .ZN(n1964) );
NAND2_X1 U2237 ( .A1(n2016), .A2(register_file_inst_reg_array_93), .ZN(n1963) );
NAND2_X1 U2238 ( .A1(n1964), .A2(n1963), .ZN(n1965) );
NOR2_X1 U2239 ( .A1(n1966), .A2(n1965), .ZN(n1968) );
NAND2_X1 U2240 ( .A1(n2021), .A2(register_file_inst_reg_array_13), .ZN(n1967) );
NAND2_X1 U2241 ( .A1(n1968), .A2(n1967), .ZN(n1969) );
NOR2_X1 U2242 ( .A1(n1970), .A2(n1969), .ZN(n1971) );
NAND2_X1 U2243 ( .A1(n1972), .A2(n1971), .ZN(reg_read_data_1_13) );
NAND2_X1 U2244 ( .A1(register_file_inst_reg_array_22), .A2(n2009), .ZN(n1984) );
NAND2_X1 U2245 ( .A1(n2010), .A2(register_file_inst_reg_array_102), .ZN(n1974) );
NAND2_X1 U2246 ( .A1(n2011), .A2(register_file_inst_reg_array_38), .ZN(n1973) );
NAND2_X1 U2247 ( .A1(n1974), .A2(n1973), .ZN(n1982) );
NOR2_X1 U2248 ( .A1(n3503), .A2(n2014), .ZN(n1978) );
NAND2_X1 U2249 ( .A1(n2015), .A2(register_file_inst_reg_array_70), .ZN(n1976) );
NAND2_X1 U2250 ( .A1(n2016), .A2(register_file_inst_reg_array_86), .ZN(n1975) );
NAND2_X1 U2251 ( .A1(n1976), .A2(n1975), .ZN(n1977) );
NOR2_X1 U2252 ( .A1(n1978), .A2(n1977), .ZN(n1980) );
NAND2_X1 U2253 ( .A1(n2021), .A2(register_file_inst_reg_array_6), .ZN(n1979) );
NAND2_X1 U2254 ( .A1(n1980), .A2(n1979), .ZN(n1981) );
NOR2_X1 U2255 ( .A1(n1982), .A2(n1981), .ZN(n1983) );
NAND2_X1 U2256 ( .A1(n1984), .A2(n1983), .ZN(reg_read_data_1_6) );
NAND2_X1 U2257 ( .A1(register_file_inst_reg_array_26), .A2(n2009), .ZN(n1996) );
NAND2_X1 U2258 ( .A1(n2010), .A2(register_file_inst_reg_array_106), .ZN(n1986) );
NAND2_X1 U2259 ( .A1(n2011), .A2(register_file_inst_reg_array_42), .ZN(n1985) );
NAND2_X1 U2260 ( .A1(n1986), .A2(n1985), .ZN(n1994) );
NOR2_X1 U2261 ( .A1(n3504), .A2(n2014), .ZN(n1990) );
NAND2_X1 U2262 ( .A1(n2015), .A2(register_file_inst_reg_array_74), .ZN(n1988) );
NAND2_X1 U2263 ( .A1(n2016), .A2(register_file_inst_reg_array_90), .ZN(n1987) );
NAND2_X1 U2264 ( .A1(n1988), .A2(n1987), .ZN(n1989) );
NOR2_X1 U2265 ( .A1(n1990), .A2(n1989), .ZN(n1992) );
NAND2_X1 U2266 ( .A1(n2021), .A2(register_file_inst_reg_array_10), .ZN(n1991) );
NAND2_X1 U2267 ( .A1(n1992), .A2(n1991), .ZN(n1993) );
NOR2_X1 U2268 ( .A1(n1994), .A2(n1993), .ZN(n1995) );
NAND2_X1 U2269 ( .A1(n1996), .A2(n1995), .ZN(reg_read_data_1_10) );
NAND2_X1 U2270 ( .A1(register_file_inst_reg_array_23), .A2(n2009), .ZN(n2008) );
NAND2_X1 U2271 ( .A1(n2010), .A2(register_file_inst_reg_array_103), .ZN(n1998) );
NAND2_X1 U2272 ( .A1(n2011), .A2(register_file_inst_reg_array_39), .ZN(n1997) );
NAND2_X1 U2273 ( .A1(n1998), .A2(n1997), .ZN(n2006) );
NOR2_X1 U2274 ( .A1(n3505), .A2(n2014), .ZN(n2002) );
NAND2_X1 U2275 ( .A1(n2015), .A2(register_file_inst_reg_array_71), .ZN(n2000) );
NAND2_X1 U2276 ( .A1(n2016), .A2(register_file_inst_reg_array_87), .ZN(n1999) );
NAND2_X1 U2277 ( .A1(n2000), .A2(n1999), .ZN(n2001) );
NOR2_X1 U2278 ( .A1(n2002), .A2(n2001), .ZN(n2004) );
NAND2_X1 U2279 ( .A1(n2021), .A2(register_file_inst_reg_array_7), .ZN(n2003) );
NAND2_X1 U2280 ( .A1(n2004), .A2(n2003), .ZN(n2005) );
NOR2_X1 U2281 ( .A1(n2006), .A2(n2005), .ZN(n2007) );
NAND2_X1 U2282 ( .A1(n2008), .A2(n2007), .ZN(reg_read_data_1_7) );
NAND2_X1 U2283 ( .A1(register_file_inst_reg_array_19), .A2(n2009), .ZN(n2027) );
NAND2_X1 U2284 ( .A1(n2010), .A2(register_file_inst_reg_array_99), .ZN(n2013) );
NAND2_X1 U2285 ( .A1(n2011), .A2(register_file_inst_reg_array_35), .ZN(n2012) );
NAND2_X1 U2286 ( .A1(n2013), .A2(n2012), .ZN(n2025) );
NOR2_X1 U2287 ( .A1(n3506), .A2(n2014), .ZN(n2020) );
NAND2_X1 U2288 ( .A1(n2015), .A2(register_file_inst_reg_array_67), .ZN(n2018) );
NAND2_X1 U2289 ( .A1(n2016), .A2(register_file_inst_reg_array_83), .ZN(n2017) );
NAND2_X1 U2290 ( .A1(n2018), .A2(n2017), .ZN(n2019) );
NOR2_X1 U2291 ( .A1(n2020), .A2(n2019), .ZN(n2023) );
NAND2_X1 U2292 ( .A1(n2021), .A2(register_file_inst_reg_array_3), .ZN(n2022) );
NAND2_X1 U2293 ( .A1(n2023), .A2(n2022), .ZN(n2024) );
NOR2_X1 U2294 ( .A1(n2025), .A2(n2024), .ZN(n2026) );
NAND2_X1 U2295 ( .A1(n2027), .A2(n2026), .ZN(reg_read_data_1_3) );
NAND2_X1 U2296 ( .A1(n3176), .A2(pc_7_), .ZN(n2067) );
NOR2_X1 U2297 ( .A1(ID_stage_inst_ir_dest_with_bubble_0), .A2(ID_stage_inst_ir_dest_with_bubble_2), .ZN(n2046) );
NOR2_X1 U2298 ( .A1(reg_read_data_1_15), .A2(reg_read_data_1_9), .ZN(n2029) );
NOR2_X1 U2299 ( .A1(reg_read_data_1_2), .A2(reg_read_data_1_0), .ZN(n2028) );
NAND2_X1 U2300 ( .A1(n2029), .A2(n2028), .ZN(n2044) );
NAND2_X1 U2301 ( .A1(ID_stage_inst_instruction_reg_14), .A2(n2030), .ZN(n2031) );
NOR2_X1 U2302 ( .A1(n2031), .A2(reg_read_data_1_4), .ZN(n2033) );
NOR2_X1 U2303 ( .A1(reg_read_data_1_5), .A2(reg_read_data_1_11), .ZN(n2032) );
NAND2_X1 U2304 ( .A1(n2033), .A2(n2032), .ZN(n2034) );
NOR2_X1 U2305 ( .A1(reg_read_data_1_12), .A2(n2034), .ZN(n2042) );
NOR2_X1 U2306 ( .A1(reg_read_data_1_1), .A2(reg_read_data_1_8), .ZN(n2036) );
NOR2_X1 U2307 ( .A1(reg_read_data_1_14), .A2(reg_read_data_1_13), .ZN(n2035) );
NAND2_X1 U2308 ( .A1(n2036), .A2(n2035), .ZN(n2040) );
NOR2_X1 U2309 ( .A1(reg_read_data_1_6), .A2(reg_read_data_1_10), .ZN(n2038) );
NOR2_X1 U2310 ( .A1(reg_read_data_1_7), .A2(reg_read_data_1_3), .ZN(n2037) );
NAND2_X1 U2311 ( .A1(n2038), .A2(n2037), .ZN(n2039) );
NOR2_X1 U2312 ( .A1(n2040), .A2(n2039), .ZN(n2041) );
NAND2_X1 U2313 ( .A1(n2042), .A2(n2041), .ZN(n2043) );
NOR2_X1 U2314 ( .A1(n2044), .A2(n2043), .ZN(n2045) );
NAND2_X1 U2315 ( .A1(n2046), .A2(n2045), .ZN(n2047) );
OR2_X1 U2316 ( .A1(ID_stage_inst_ir_dest_with_bubble_1), .A2(n2047), .ZN(n2049) );
NOR2_X1 U2317 ( .A1(n3509), .A2(n2049), .ZN(n2062) );
AND2_X1 U2318 ( .A1(n2062), .A2(pc_6_), .ZN(n2061) );
AND2_X1 U2319 ( .A1(n2062), .A2(pc_5_), .ZN(n2059) );
NOR2_X1 U2320 ( .A1(n2049), .A2(n3512), .ZN(n2055) );
AND2_X1 U2321 ( .A1(pc_4_), .A2(n2055), .ZN(n2057) );
NOR2_X1 U2322 ( .A1(n2049), .A2(n3513), .ZN(n2052) );
AND2_X1 U2323 ( .A1(pc_3_), .A2(n2052), .ZN(n2054) );
NOR2_X1 U2324 ( .A1(n2049), .A2(n3514), .ZN(n2048) );
AND2_X1 U2325 ( .A1(pc_1_), .A2(n2048), .ZN(n2051) );
XOR2_X1 U2326 ( .A(pc_1_), .B(n2048), .Z(n2114) );
OR2_X1 U2327 ( .A1(branch_offset_imm_0), .A2(n2049), .ZN(n2092) );
AND2_X1 U2328 ( .A1(pc_0_), .A2(n2092), .ZN(n2113) );
AND2_X1 U2329 ( .A1(n2114), .A2(n2113), .ZN(n2050) );
OR2_X1 U2330 ( .A1(n2051), .A2(n2050), .ZN(n2088) );
AND2_X1 U2331 ( .A1(n2088), .A2(pc_2_), .ZN(n2084) );
XOR2_X1 U2332 ( .A(pc_3_), .B(n2052), .Z(n2083) );
AND2_X1 U2333 ( .A1(n2084), .A2(n2083), .ZN(n2053) );
OR2_X1 U2334 ( .A1(n2054), .A2(n2053), .ZN(n2079) );
XOR2_X1 U2335 ( .A(pc_4_), .B(n2055), .Z(n2078) );
OR2_X1 U2336 ( .A1(n2057), .A2(n2056), .ZN(n2074) );
XOR2_X1 U2337 ( .A(n2062), .B(pc_5_), .Z(n2073) );
AND2_X1 U2338 ( .A1(n2074), .A2(n2073), .ZN(n2058) );
OR2_X1 U2339 ( .A1(n2059), .A2(n2058), .ZN(n2069) );
XOR2_X1 U2340 ( .A(n2062), .B(pc_6_), .Z(n2068) );
AND2_X1 U2341 ( .A1(n2069), .A2(n2068), .ZN(n2060) );
XOR2_X1 U2342 ( .A(n2062), .B(pc_7_), .Z(n2063) );
XOR2_X1 U2343 ( .A(n2064), .B(n2063), .Z(n2065) );
NAND2_X1 U2344 ( .A1(n2065), .A2(n3163), .ZN(n2066) );
NAND2_X1 U2345 ( .A1(n2067), .A2(n2066), .ZN(n1727) );
NAND2_X1 U2346 ( .A1(n3176), .A2(pc_6_), .ZN(n2072) );
XOR2_X1 U2347 ( .A(n2069), .B(n2068), .Z(n2070) );
NAND2_X1 U2348 ( .A1(n2070), .A2(n3163), .ZN(n2071) );
NAND2_X1 U2349 ( .A1(n2072), .A2(n2071), .ZN(n1728) );
NAND2_X1 U2350 ( .A1(n3176), .A2(pc_5_), .ZN(n2077) );
XOR2_X1 U2351 ( .A(n2074), .B(n2073), .Z(n2075) );
NAND2_X1 U2352 ( .A1(n2075), .A2(n3163), .ZN(n2076) );
NAND2_X1 U2353 ( .A1(n2077), .A2(n2076), .ZN(n1729) );
NAND2_X1 U2354 ( .A1(n3176), .A2(pc_4_), .ZN(n2082) );
XOR2_X1 U2355 ( .A(n2079), .B(n2078), .Z(n2080) );
NAND2_X1 U2356 ( .A1(n2080), .A2(n3163), .ZN(n2081) );
NAND2_X1 U2357 ( .A1(n2082), .A2(n2081), .ZN(n1730) );
NAND2_X1 U2358 ( .A1(n3176), .A2(pc_3_), .ZN(n2087) );
XOR2_X1 U2359 ( .A(n2084), .B(n2083), .Z(n2085) );
NAND2_X1 U2360 ( .A1(n2085), .A2(n3163), .ZN(n2086) );
NAND2_X1 U2361 ( .A1(n2087), .A2(n2086), .ZN(n1731) );
NAND2_X1 U2362 ( .A1(n3176), .A2(pc_2_), .ZN(n2091) );
XOR2_X1 U2363 ( .A(n2088), .B(pc_2_), .Z(n2089) );
NAND2_X1 U2364 ( .A1(n2089), .A2(n3163), .ZN(n2090) );
NAND2_X1 U2365 ( .A1(n2091), .A2(n2090), .ZN(n1732) );
NAND2_X1 U2366 ( .A1(n3176), .A2(pc_0_), .ZN(n2095) );
XOR2_X1 U2367 ( .A(pc_0_), .B(n2092), .Z(n2093) );
NAND2_X1 U2368 ( .A1(n2093), .A2(n3163), .ZN(n2094) );
NAND2_X1 U2369 ( .A1(n2095), .A2(n2094), .ZN(n1734) );
NAND2_X1 U2370 ( .A1(branch_offset_imm_5), .A2(n3176), .ZN(n2099) );
NOR2_X1 U2371 ( .A1(n3176), .A2(pc_6_), .ZN(n2111) );
NOR2_X1 U2372 ( .A1(pc_7_), .A2(pc_5_), .ZN(n2105) );
NOR2_X1 U2373 ( .A1(pc_4_), .A2(pc_3_), .ZN(n2096) );
AND2_X1 U2374 ( .A1(n2105), .A2(n2096), .ZN(n2097) );
NAND2_X1 U2375 ( .A1(n2111), .A2(n2097), .ZN(n3144) );
NAND2_X1 U2376 ( .A1(pc_1_), .A2(n2118), .ZN(n3153) );
INV_X1 U2377 ( .A(n3153), .ZN(n2098) );
NAND2_X1 U2378 ( .A1(pc_2_), .A2(n2098), .ZN(n3141) );
NAND2_X1 U2379 ( .A1(n2099), .A2(n3141), .ZN(n1722) );
OR2_X1 U2380 ( .A1(pc_1_), .A2(n3481), .ZN(n2100) );
NAND2_X1 U2381 ( .A1(n2118), .A2(n2100), .ZN(n2102) );
NAND2_X1 U2382 ( .A1(branch_offset_imm_3), .A2(n3176), .ZN(n2101) );
NAND2_X1 U2383 ( .A1(n2102), .A2(n2101), .ZN(n1724) );
NAND2_X1 U2384 ( .A1(pc_2_), .A2(n2118), .ZN(n2103) );
OR2_X1 U2385 ( .A1(pc_1_), .A2(n2103), .ZN(n3143) );
NAND2_X1 U2386 ( .A1(branch_offset_imm_1), .A2(n3176), .ZN(n2104) );
NAND2_X1 U2387 ( .A1(n3143), .A2(n2104), .ZN(n1725) );
NAND2_X1 U2388 ( .A1(n2105), .A2(n3481), .ZN(n2109) );
NOR2_X1 U2389 ( .A1(pc_1_), .A2(pc_0_), .ZN(n2107) );
NOR2_X1 U2390 ( .A1(pc_4_), .A2(n3511), .ZN(n2106) );
NAND2_X1 U2391 ( .A1(n2107), .A2(n2106), .ZN(n2108) );
NOR2_X1 U2392 ( .A1(n2109), .A2(n2108), .ZN(n2110) );
NAND2_X1 U2393 ( .A1(n2111), .A2(n2110), .ZN(n3167) );
NAND2_X1 U2394 ( .A1(n3176), .A2(branch_offset_imm_0), .ZN(n2112) );
NAND2_X1 U2395 ( .A1(n3167), .A2(n2112), .ZN(n1726) );
NAND2_X1 U2396 ( .A1(n3176), .A2(pc_1_), .ZN(n2117) );
XOR2_X1 U2397 ( .A(n2114), .B(n2113), .Z(n2115) );
NAND2_X1 U2398 ( .A1(n2115), .A2(n3163), .ZN(n2116) );
NAND2_X1 U2399 ( .A1(n2117), .A2(n2116), .ZN(n1733) );
NAND2_X1 U2400 ( .A1(branch_offset_imm_4), .A2(n3176), .ZN(n2119) );
NAND2_X1 U2401 ( .A1(pc_0_), .A2(n2118), .ZN(n3131) );
INV_X1 U2402 ( .A(n3131), .ZN(n3180) );
NAND2_X1 U2403 ( .A1(pc_1_), .A2(n3180), .ZN(n3173) );
NAND2_X1 U2404 ( .A1(n2119), .A2(n3173), .ZN(n1723) );
NAND2_X1 U2405 ( .A1(register_file_inst_reg_array_23), .A2(n2306), .ZN(n2121) );
NAND2_X1 U2406 ( .A1(register_file_inst_reg_array_103), .A2(n2307), .ZN(n2120) );
NAND2_X1 U2407 ( .A1(n2121), .A2(n2120), .ZN(n2129) );
NOR2_X1 U2408 ( .A1(n2310), .A2(n3505), .ZN(n2125) );
NAND2_X1 U2409 ( .A1(register_file_inst_reg_array_71), .A2(n2311), .ZN(n2123) );
NAND2_X1 U2410 ( .A1(register_file_inst_reg_array_87), .A2(n2312), .ZN(n2122) );
NAND2_X1 U2411 ( .A1(n2123), .A2(n2122), .ZN(n2124) );
NOR2_X1 U2412 ( .A1(n2125), .A2(n2124), .ZN(n2127) );
NAND2_X1 U2413 ( .A1(register_file_inst_reg_array_39), .A2(n2317), .ZN(n2126) );
NAND2_X1 U2414 ( .A1(n2127), .A2(n2126), .ZN(n2128) );
NOR2_X1 U2415 ( .A1(n2129), .A2(n2128), .ZN(n2131) );
NAND2_X1 U2416 ( .A1(n2322), .A2(register_file_inst_reg_array_7), .ZN(n2130) );
NAND2_X1 U2417 ( .A1(n2131), .A2(n2130), .ZN(reg_read_data_2_7) );
NAND2_X1 U2418 ( .A1(n2325), .A2(reg_read_data_2_7), .ZN(n2132) );
NAND2_X1 U2419 ( .A1(branch_offset_imm_5), .A2(n2326), .ZN(n2262) );
NAND2_X1 U2420 ( .A1(n2132), .A2(n2262), .ZN(ID_stage_inst_ex_alu_src2_7) );
NAND2_X1 U2421 ( .A1(register_file_inst_reg_array_25), .A2(n2306), .ZN(n2134) );
NAND2_X1 U2422 ( .A1(register_file_inst_reg_array_105), .A2(n2307), .ZN(n2133) );
NAND2_X1 U2423 ( .A1(n2134), .A2(n2133), .ZN(n2142) );
NOR2_X1 U2424 ( .A1(n2310), .A2(n3493), .ZN(n2138) );
NAND2_X1 U2425 ( .A1(register_file_inst_reg_array_73), .A2(n2311), .ZN(n2136) );
NAND2_X1 U2426 ( .A1(register_file_inst_reg_array_89), .A2(n2312), .ZN(n2135) );
NAND2_X1 U2427 ( .A1(n2136), .A2(n2135), .ZN(n2137) );
NOR2_X1 U2428 ( .A1(n2138), .A2(n2137), .ZN(n2140) );
NAND2_X1 U2429 ( .A1(register_file_inst_reg_array_41), .A2(n2317), .ZN(n2139) );
NAND2_X1 U2430 ( .A1(n2140), .A2(n2139), .ZN(n2141) );
NOR2_X1 U2431 ( .A1(n2142), .A2(n2141), .ZN(n2144) );
NAND2_X1 U2432 ( .A1(n2322), .A2(register_file_inst_reg_array_9), .ZN(n2143) );
NAND2_X1 U2433 ( .A1(n2144), .A2(n2143), .ZN(reg_read_data_2_9) );
NAND2_X1 U2434 ( .A1(n2325), .A2(reg_read_data_2_9), .ZN(n2145) );
NAND2_X1 U2435 ( .A1(n2145), .A2(n2262), .ZN(ID_stage_inst_ex_alu_src2_9) );
NAND2_X1 U2436 ( .A1(register_file_inst_reg_array_28), .A2(n2306), .ZN(n2147) );
NAND2_X1 U2437 ( .A1(register_file_inst_reg_array_108), .A2(n2307), .ZN(n2146) );
NAND2_X1 U2438 ( .A1(n2147), .A2(n2146), .ZN(n2155) );
NOR2_X1 U2439 ( .A1(n2310), .A2(n3495), .ZN(n2151) );
NAND2_X1 U2440 ( .A1(register_file_inst_reg_array_76), .A2(n2311), .ZN(n2149) );
NAND2_X1 U2441 ( .A1(register_file_inst_reg_array_92), .A2(n2312), .ZN(n2148) );
NAND2_X1 U2442 ( .A1(n2149), .A2(n2148), .ZN(n2150) );
NOR2_X1 U2443 ( .A1(n2151), .A2(n2150), .ZN(n2153) );
NAND2_X1 U2444 ( .A1(register_file_inst_reg_array_44), .A2(n2317), .ZN(n2152) );
NAND2_X1 U2445 ( .A1(n2153), .A2(n2152), .ZN(n2154) );
NOR2_X1 U2446 ( .A1(n2155), .A2(n2154), .ZN(n2157) );
NAND2_X1 U2447 ( .A1(n2322), .A2(register_file_inst_reg_array_12), .ZN(n2156) );
NAND2_X1 U2448 ( .A1(n2157), .A2(n2156), .ZN(reg_read_data_2_12) );
NAND2_X1 U2449 ( .A1(n2325), .A2(reg_read_data_2_12), .ZN(n2158) );
NAND2_X1 U2450 ( .A1(n2158), .A2(n2262), .ZN(ID_stage_inst_ex_alu_src2_12) );
NAND2_X1 U2451 ( .A1(register_file_inst_reg_array_27), .A2(n2306), .ZN(n2160) );
NAND2_X1 U2452 ( .A1(register_file_inst_reg_array_107), .A2(n2307), .ZN(n2159) );
NAND2_X1 U2453 ( .A1(n2160), .A2(n2159), .ZN(n2168) );
NOR2_X1 U2454 ( .A1(n2310), .A2(n3498), .ZN(n2164) );
NAND2_X1 U2455 ( .A1(register_file_inst_reg_array_75), .A2(n2311), .ZN(n2162) );
NAND2_X1 U2456 ( .A1(register_file_inst_reg_array_91), .A2(n2312), .ZN(n2161) );
NAND2_X1 U2457 ( .A1(n2162), .A2(n2161), .ZN(n2163) );
NOR2_X1 U2458 ( .A1(n2164), .A2(n2163), .ZN(n2166) );
NAND2_X1 U2459 ( .A1(register_file_inst_reg_array_43), .A2(n2317), .ZN(n2165) );
NAND2_X1 U2460 ( .A1(n2166), .A2(n2165), .ZN(n2167) );
NOR2_X1 U2461 ( .A1(n2168), .A2(n2167), .ZN(n2170) );
NAND2_X1 U2462 ( .A1(n2322), .A2(register_file_inst_reg_array_11), .ZN(n2169) );
NAND2_X1 U2463 ( .A1(n2170), .A2(n2169), .ZN(reg_read_data_2_11) );
NAND2_X1 U2464 ( .A1(n2325), .A2(reg_read_data_2_11), .ZN(n2171) );
NAND2_X1 U2465 ( .A1(n2171), .A2(n2262), .ZN(ID_stage_inst_ex_alu_src2_11) );
NAND2_X1 U2466 ( .A1(register_file_inst_reg_array_30), .A2(n2306), .ZN(n2173) );
NAND2_X1 U2467 ( .A1(register_file_inst_reg_array_110), .A2(n2307), .ZN(n2172) );
NAND2_X1 U2468 ( .A1(n2173), .A2(n2172), .ZN(n2181) );
NOR2_X1 U2469 ( .A1(n2310), .A2(n3501), .ZN(n2177) );
NAND2_X1 U2470 ( .A1(register_file_inst_reg_array_78), .A2(n2311), .ZN(n2175) );
NAND2_X1 U2471 ( .A1(register_file_inst_reg_array_94), .A2(n2312), .ZN(n2174) );
NAND2_X1 U2472 ( .A1(n2175), .A2(n2174), .ZN(n2176) );
NOR2_X1 U2473 ( .A1(n2177), .A2(n2176), .ZN(n2179) );
NAND2_X1 U2474 ( .A1(register_file_inst_reg_array_46), .A2(n2317), .ZN(n2178) );
NAND2_X1 U2475 ( .A1(n2179), .A2(n2178), .ZN(n2180) );
NOR2_X1 U2476 ( .A1(n2181), .A2(n2180), .ZN(n2183) );
NAND2_X1 U2477 ( .A1(n2322), .A2(register_file_inst_reg_array_14), .ZN(n2182) );
NAND2_X1 U2478 ( .A1(n2183), .A2(n2182), .ZN(reg_read_data_2_14) );
NAND2_X1 U2479 ( .A1(n2325), .A2(reg_read_data_2_14), .ZN(n2184) );
NAND2_X1 U2480 ( .A1(n2184), .A2(n2262), .ZN(ID_stage_inst_ex_alu_src2_14) );
NAND2_X1 U2481 ( .A1(register_file_inst_reg_array_26), .A2(n2306), .ZN(n2186) );
NAND2_X1 U2482 ( .A1(register_file_inst_reg_array_106), .A2(n2307), .ZN(n2185) );
NAND2_X1 U2483 ( .A1(n2186), .A2(n2185), .ZN(n2194) );
NOR2_X1 U2484 ( .A1(n2310), .A2(n3504), .ZN(n2190) );
NAND2_X1 U2485 ( .A1(register_file_inst_reg_array_74), .A2(n2311), .ZN(n2188) );
NAND2_X1 U2486 ( .A1(register_file_inst_reg_array_90), .A2(n2312), .ZN(n2187) );
NAND2_X1 U2487 ( .A1(n2188), .A2(n2187), .ZN(n2189) );
NOR2_X1 U2488 ( .A1(n2190), .A2(n2189), .ZN(n2192) );
NAND2_X1 U2489 ( .A1(register_file_inst_reg_array_42), .A2(n2317), .ZN(n2191) );
NAND2_X1 U2490 ( .A1(n2192), .A2(n2191), .ZN(n2193) );
NOR2_X1 U2491 ( .A1(n2194), .A2(n2193), .ZN(n2196) );
NAND2_X1 U2492 ( .A1(n2322), .A2(register_file_inst_reg_array_10), .ZN(n2195) );
NAND2_X1 U2493 ( .A1(n2196), .A2(n2195), .ZN(reg_read_data_2_10) );
NAND2_X1 U2494 ( .A1(n2325), .A2(reg_read_data_2_10), .ZN(n2197) );
NAND2_X1 U2495 ( .A1(n2197), .A2(n2262), .ZN(ID_stage_inst_ex_alu_src2_10) );
NAND2_X1 U2496 ( .A1(register_file_inst_reg_array_24), .A2(n2306), .ZN(n2199) );
NAND2_X1 U2497 ( .A1(register_file_inst_reg_array_104), .A2(n2307), .ZN(n2198) );
NAND2_X1 U2498 ( .A1(n2199), .A2(n2198), .ZN(n2207) );
NOR2_X1 U2499 ( .A1(n2310), .A2(n3500), .ZN(n2203) );
NAND2_X1 U2500 ( .A1(register_file_inst_reg_array_72), .A2(n2311), .ZN(n2201) );
NAND2_X1 U2501 ( .A1(register_file_inst_reg_array_88), .A2(n2312), .ZN(n2200) );
NAND2_X1 U2502 ( .A1(n2201), .A2(n2200), .ZN(n2202) );
NOR2_X1 U2503 ( .A1(n2203), .A2(n2202), .ZN(n2205) );
NAND2_X1 U2504 ( .A1(register_file_inst_reg_array_40), .A2(n2317), .ZN(n2204) );
NAND2_X1 U2505 ( .A1(n2205), .A2(n2204), .ZN(n2206) );
NOR2_X1 U2506 ( .A1(n2207), .A2(n2206), .ZN(n2209) );
NAND2_X1 U2507 ( .A1(n2322), .A2(register_file_inst_reg_array_8), .ZN(n2208) );
NAND2_X1 U2508 ( .A1(n2209), .A2(n2208), .ZN(reg_read_data_2_8) );
NAND2_X1 U2509 ( .A1(n2325), .A2(reg_read_data_2_8), .ZN(n2210) );
NAND2_X1 U2510 ( .A1(n2210), .A2(n2262), .ZN(ID_stage_inst_ex_alu_src2_8) );
NAND2_X1 U2511 ( .A1(register_file_inst_reg_array_22), .A2(n2306), .ZN(n2212) );
NAND2_X1 U2512 ( .A1(register_file_inst_reg_array_102), .A2(n2307), .ZN(n2211) );
NAND2_X1 U2513 ( .A1(n2212), .A2(n2211), .ZN(n2220) );
NOR2_X1 U2514 ( .A1(n2310), .A2(n3503), .ZN(n2216) );
NAND2_X1 U2515 ( .A1(register_file_inst_reg_array_70), .A2(n2311), .ZN(n2214) );
NAND2_X1 U2516 ( .A1(register_file_inst_reg_array_86), .A2(n2312), .ZN(n2213) );
NAND2_X1 U2517 ( .A1(n2214), .A2(n2213), .ZN(n2215) );
NOR2_X1 U2518 ( .A1(n2216), .A2(n2215), .ZN(n2218) );
NAND2_X1 U2519 ( .A1(register_file_inst_reg_array_38), .A2(n2317), .ZN(n2217) );
NAND2_X1 U2520 ( .A1(n2218), .A2(n2217), .ZN(n2219) );
NOR2_X1 U2521 ( .A1(n2220), .A2(n2219), .ZN(n2222) );
NAND2_X1 U2522 ( .A1(n2322), .A2(register_file_inst_reg_array_6), .ZN(n2221) );
NAND2_X1 U2523 ( .A1(n2222), .A2(n2221), .ZN(reg_read_data_2_6) );
NAND2_X1 U2524 ( .A1(n2325), .A2(reg_read_data_2_6), .ZN(n2223) );
NAND2_X1 U2525 ( .A1(n2223), .A2(n2262), .ZN(ID_stage_inst_ex_alu_src2_6) );
NAND2_X1 U2526 ( .A1(register_file_inst_reg_array_29), .A2(n2306), .ZN(n2225) );
NAND2_X1 U2527 ( .A1(register_file_inst_reg_array_109), .A2(n2307), .ZN(n2224) );
NAND2_X1 U2528 ( .A1(n2225), .A2(n2224), .ZN(n2233) );
NOR2_X1 U2529 ( .A1(n2310), .A2(n3502), .ZN(n2229) );
NAND2_X1 U2530 ( .A1(register_file_inst_reg_array_77), .A2(n2311), .ZN(n2227) );
NAND2_X1 U2531 ( .A1(register_file_inst_reg_array_93), .A2(n2312), .ZN(n2226) );
NAND2_X1 U2532 ( .A1(n2227), .A2(n2226), .ZN(n2228) );
NOR2_X1 U2533 ( .A1(n2229), .A2(n2228), .ZN(n2231) );
NAND2_X1 U2534 ( .A1(register_file_inst_reg_array_45), .A2(n2317), .ZN(n2230) );
NAND2_X1 U2535 ( .A1(n2231), .A2(n2230), .ZN(n2232) );
NOR2_X1 U2536 ( .A1(n2233), .A2(n2232), .ZN(n2235) );
NAND2_X1 U2537 ( .A1(n2322), .A2(register_file_inst_reg_array_13), .ZN(n2234) );
NAND2_X1 U2538 ( .A1(n2235), .A2(n2234), .ZN(reg_read_data_2_13) );
NAND2_X1 U2539 ( .A1(n2325), .A2(reg_read_data_2_13), .ZN(n2236) );
NAND2_X1 U2540 ( .A1(n2236), .A2(n2262), .ZN(ID_stage_inst_ex_alu_src2_13) );
NAND2_X1 U2541 ( .A1(register_file_inst_reg_array_21), .A2(n2306), .ZN(n2238) );
NAND2_X1 U2542 ( .A1(register_file_inst_reg_array_101), .A2(n2307), .ZN(n2237) );
NAND2_X1 U2543 ( .A1(n2238), .A2(n2237), .ZN(n2246) );
NOR2_X1 U2544 ( .A1(n2310), .A2(n3497), .ZN(n2242) );
NAND2_X1 U2545 ( .A1(register_file_inst_reg_array_69), .A2(n2311), .ZN(n2240) );
NAND2_X1 U2546 ( .A1(register_file_inst_reg_array_85), .A2(n2312), .ZN(n2239) );
NAND2_X1 U2547 ( .A1(n2240), .A2(n2239), .ZN(n2241) );
NOR2_X1 U2548 ( .A1(n2242), .A2(n2241), .ZN(n2244) );
NAND2_X1 U2549 ( .A1(register_file_inst_reg_array_37), .A2(n2317), .ZN(n2243) );
NAND2_X1 U2550 ( .A1(n2244), .A2(n2243), .ZN(n2245) );
NOR2_X1 U2551 ( .A1(n2246), .A2(n2245), .ZN(n2248) );
NAND2_X1 U2552 ( .A1(n2322), .A2(register_file_inst_reg_array_5), .ZN(n2247) );
NAND2_X1 U2553 ( .A1(n2248), .A2(n2247), .ZN(reg_read_data_2_5) );
NAND2_X1 U2554 ( .A1(n2325), .A2(reg_read_data_2_5), .ZN(n2249) );
NAND2_X1 U2555 ( .A1(n2249), .A2(n2262), .ZN(ID_stage_inst_ex_alu_src2_5) );
NAND2_X1 U2556 ( .A1(register_file_inst_reg_array_31), .A2(n2306), .ZN(n2251) );
NAND2_X1 U2557 ( .A1(register_file_inst_reg_array_111), .A2(n2307), .ZN(n2250) );
NAND2_X1 U2558 ( .A1(n2251), .A2(n2250), .ZN(n2259) );
NOR2_X1 U2559 ( .A1(n2310), .A2(n3492), .ZN(n2255) );
NAND2_X1 U2560 ( .A1(register_file_inst_reg_array_79), .A2(n2311), .ZN(n2253) );
NAND2_X1 U2561 ( .A1(register_file_inst_reg_array_95), .A2(n2312), .ZN(n2252) );
NAND2_X1 U2562 ( .A1(n2253), .A2(n2252), .ZN(n2254) );
NOR2_X1 U2563 ( .A1(n2255), .A2(n2254), .ZN(n2257) );
NAND2_X1 U2564 ( .A1(register_file_inst_reg_array_47), .A2(n2317), .ZN(n2256) );
NAND2_X1 U2565 ( .A1(n2257), .A2(n2256), .ZN(n2258) );
NOR2_X1 U2566 ( .A1(n2259), .A2(n2258), .ZN(n2261) );
NAND2_X1 U2567 ( .A1(n2322), .A2(register_file_inst_reg_array_15), .ZN(n2260) );
NAND2_X1 U2568 ( .A1(n2261), .A2(n2260), .ZN(reg_read_data_2_15) );
NAND2_X1 U2569 ( .A1(n2325), .A2(reg_read_data_2_15), .ZN(n2263) );
NAND2_X1 U2570 ( .A1(n2263), .A2(n2262), .ZN(ID_stage_inst_ex_alu_src2_15) );
NAND2_X1 U2571 ( .A1(register_file_inst_reg_array_20), .A2(n2306), .ZN(n2265) );
NAND2_X1 U2572 ( .A1(register_file_inst_reg_array_100), .A2(n2307), .ZN(n2264) );
NAND2_X1 U2573 ( .A1(n2265), .A2(n2264), .ZN(n2273) );
NOR2_X1 U2574 ( .A1(n2310), .A2(n3496), .ZN(n2269) );
NAND2_X1 U2575 ( .A1(register_file_inst_reg_array_68), .A2(n2311), .ZN(n2267) );
NAND2_X1 U2576 ( .A1(register_file_inst_reg_array_84), .A2(n2312), .ZN(n2266) );
NAND2_X1 U2577 ( .A1(n2267), .A2(n2266), .ZN(n2268) );
NOR2_X1 U2578 ( .A1(n2269), .A2(n2268), .ZN(n2271) );
NAND2_X1 U2579 ( .A1(register_file_inst_reg_array_36), .A2(n2317), .ZN(n2270) );
NAND2_X1 U2580 ( .A1(n2271), .A2(n2270), .ZN(n2272) );
NOR2_X1 U2581 ( .A1(n2273), .A2(n2272), .ZN(n2275) );
NAND2_X1 U2582 ( .A1(n2322), .A2(register_file_inst_reg_array_4), .ZN(n2274) );
NAND2_X1 U2583 ( .A1(n2275), .A2(n2274), .ZN(reg_read_data_2_4) );
NAND2_X1 U2584 ( .A1(n2325), .A2(reg_read_data_2_4), .ZN(n2277) );
NAND2_X1 U2585 ( .A1(branch_offset_imm_4), .A2(n2326), .ZN(n2276) );
NAND2_X1 U2586 ( .A1(n2277), .A2(n2276), .ZN(ID_stage_inst_ex_alu_src2_4) );
NAND2_X1 U2587 ( .A1(register_file_inst_reg_array_96), .A2(n2307), .ZN(n2279) );
NAND2_X1 U2588 ( .A1(register_file_inst_reg_array_16), .A2(n2306), .ZN(n2278) );
NAND2_X1 U2589 ( .A1(n2279), .A2(n2278), .ZN(n2287) );
NOR2_X1 U2590 ( .A1(n3491), .A2(n2310), .ZN(n2283) );
NAND2_X1 U2591 ( .A1(n2311), .A2(register_file_inst_reg_array_64), .ZN(n2281) );
NAND2_X1 U2592 ( .A1(n2312), .A2(register_file_inst_reg_array_80), .ZN(n2280) );
NAND2_X1 U2593 ( .A1(n2281), .A2(n2280), .ZN(n2282) );
NOR2_X1 U2594 ( .A1(n2283), .A2(n2282), .ZN(n2285) );
NAND2_X1 U2595 ( .A1(n2317), .A2(register_file_inst_reg_array_32), .ZN(n2284) );
NAND2_X1 U2596 ( .A1(n2285), .A2(n2284), .ZN(n2286) );
NOR2_X1 U2597 ( .A1(n2287), .A2(n2286), .ZN(n2289) );
NAND2_X1 U2598 ( .A1(register_file_inst_reg_array_0), .A2(n2322), .ZN(n2288) );
NAND2_X1 U2599 ( .A1(n2289), .A2(n2288), .ZN(reg_read_data_2_0) );
NAND2_X1 U2600 ( .A1(n2325), .A2(reg_read_data_2_0), .ZN(n2291) );
NAND2_X1 U2601 ( .A1(n2326), .A2(branch_offset_imm_0), .ZN(n2290) );
NAND2_X1 U2602 ( .A1(n2291), .A2(n2290), .ZN(ID_stage_inst_ex_alu_src2_0) );
NAND2_X1 U2603 ( .A1(register_file_inst_reg_array_19), .A2(n2306), .ZN(n2293) );
NAND2_X1 U2604 ( .A1(register_file_inst_reg_array_99), .A2(n2307), .ZN(n2292) );
NAND2_X1 U2605 ( .A1(n2293), .A2(n2292), .ZN(n2301) );
NOR2_X1 U2606 ( .A1(n2310), .A2(n3506), .ZN(n2297) );
NAND2_X1 U2607 ( .A1(register_file_inst_reg_array_67), .A2(n2311), .ZN(n2295) );
NAND2_X1 U2608 ( .A1(register_file_inst_reg_array_83), .A2(n2312), .ZN(n2294) );
NAND2_X1 U2609 ( .A1(n2295), .A2(n2294), .ZN(n2296) );
NOR2_X1 U2610 ( .A1(n2297), .A2(n2296), .ZN(n2299) );
NAND2_X1 U2611 ( .A1(register_file_inst_reg_array_35), .A2(n2317), .ZN(n2298) );
NAND2_X1 U2612 ( .A1(n2299), .A2(n2298), .ZN(n2300) );
NOR2_X1 U2613 ( .A1(n2301), .A2(n2300), .ZN(n2303) );
NAND2_X1 U2614 ( .A1(n2322), .A2(register_file_inst_reg_array_3), .ZN(n2302) );
NAND2_X1 U2615 ( .A1(n2303), .A2(n2302), .ZN(reg_read_data_2_3) );
NAND2_X1 U2616 ( .A1(n2325), .A2(reg_read_data_2_3), .ZN(n2305) );
NAND2_X1 U2617 ( .A1(branch_offset_imm_3), .A2(n2326), .ZN(n2304) );
NAND2_X1 U2618 ( .A1(n2305), .A2(n2304), .ZN(ID_stage_inst_ex_alu_src2_3) );
NAND2_X1 U2619 ( .A1(register_file_inst_reg_array_17), .A2(n2306), .ZN(n2309) );
NAND2_X1 U2620 ( .A1(register_file_inst_reg_array_97), .A2(n2307), .ZN(n2308) );
NAND2_X1 U2621 ( .A1(n2309), .A2(n2308), .ZN(n2321) );
NOR2_X1 U2622 ( .A1(n2310), .A2(n3499), .ZN(n2316) );
NAND2_X1 U2623 ( .A1(register_file_inst_reg_array_65), .A2(n2311), .ZN(n2314) );
NAND2_X1 U2624 ( .A1(register_file_inst_reg_array_81), .A2(n2312), .ZN(n2313) );
NAND2_X1 U2625 ( .A1(n2314), .A2(n2313), .ZN(n2315) );
NOR2_X1 U2626 ( .A1(n2316), .A2(n2315), .ZN(n2319) );
NAND2_X1 U2627 ( .A1(register_file_inst_reg_array_33), .A2(n2317), .ZN(n2318) );
NAND2_X1 U2628 ( .A1(n2319), .A2(n2318), .ZN(n2320) );
NOR2_X1 U2629 ( .A1(n2321), .A2(n2320), .ZN(n2324) );
NAND2_X1 U2630 ( .A1(n2322), .A2(register_file_inst_reg_array_1), .ZN(n2323) );
NAND2_X1 U2631 ( .A1(n2324), .A2(n2323), .ZN(reg_read_data_2_1) );
NAND2_X1 U2632 ( .A1(n2325), .A2(reg_read_data_2_1), .ZN(n2328) );
NAND2_X1 U2633 ( .A1(branch_offset_imm_1), .A2(n2326), .ZN(n2327) );
NAND2_X1 U2634 ( .A1(n2328), .A2(n2327), .ZN(ID_stage_inst_ex_alu_src2_1) );
NOR2_X1 U2635 ( .A1(n2329), .A2(n2349), .ZN(n2338) );
NAND2_X1 U2636 ( .A1(n2338), .A2(n3518), .ZN(n2343) );
NOR2_X1 U2637 ( .A1(rst), .A2(n2336), .ZN(n2340) );
NAND2_X1 U2638 ( .A1(n2344), .A2(n2346), .ZN(n2330) );
NAND2_X1 U2639 ( .A1(n2340), .A2(n2330), .ZN(n2357) );
NAND2_X1 U2640 ( .A1(n2331), .A2(n2350), .ZN(n2332) );
NAND2_X1 U2641 ( .A1(n2343), .A2(n2332), .ZN(ID_stage_inst_ex_alu_cmd_0) );
NOR2_X1 U2642 ( .A1(n2350), .A2(n2346), .ZN(n2352) );
NOR2_X1 U2643 ( .A1(n2344), .A2(n2333), .ZN(n2334) );
NOR2_X1 U2644 ( .A1(n2352), .A2(n2334), .ZN(n2335) );
NOR2_X1 U2645 ( .A1(n2336), .A2(n2335), .ZN(n2337) );
NOR2_X1 U2646 ( .A1(n2338), .A2(n2337), .ZN(n2339) );
NOR2_X1 U2647 ( .A1(rst), .A2(n2339), .ZN(ID_stage_inst_ex_alu_cmd_1) );
NAND2_X1 U2648 ( .A1(n2341), .A2(n2340), .ZN(n2342) );
NAND2_X1 U2649 ( .A1(n2343), .A2(n2342), .ZN(ID_stage_inst_ex_alu_cmd_2) );
NOR2_X1 U2650 ( .A1(n2346), .A2(n2345), .ZN(n2347) );
NAND2_X1 U2651 ( .A1(n2347), .A2(n2350), .ZN(n2348) );
NOR2_X1 U2652 ( .A1(n2353), .A2(n2348), .ZN(ID_stage_inst_write_back_result_mux) );
NOR2_X1 U2653 ( .A1(n2352), .A2(n2351), .ZN(n2355) );
NOR2_X1 U2654 ( .A1(n2353), .A2(rst), .ZN(n2354) );
NAND2_X1 U2655 ( .A1(n2355), .A2(n2354), .ZN(n2356) );
NAND2_X1 U2656 ( .A1(n2357), .A2(n2356), .ZN(ID_stage_inst_write_back_en) );
AND2_X1 U2657 ( .A1(EX_pipeline_reg_out_22), .A2(n3518), .ZN(MEM_stage_inst_N24) );
AND2_X1 U2658 ( .A1(EX_pipeline_reg_out_23), .A2(n3521), .ZN(MEM_stage_inst_N25) );
AND2_X1 U2659 ( .A1(EX_pipeline_reg_out_24), .A2(n3518), .ZN(MEM_stage_inst_N26) );
AND2_X1 U2660 ( .A1(EX_pipeline_reg_out_25), .A2(n3518), .ZN(MEM_stage_inst_N27) );
AND2_X1 U2661 ( .A1(EX_pipeline_reg_out_26), .A2(n3518), .ZN(MEM_stage_inst_N28) );
AND2_X1 U2662 ( .A1(EX_pipeline_reg_out_27), .A2(n3521), .ZN(MEM_stage_inst_N29) );
AND2_X1 U2663 ( .A1(EX_pipeline_reg_out_28), .A2(n3518), .ZN(MEM_stage_inst_N30) );
AND2_X1 U2664 ( .A1(EX_pipeline_reg_out_29), .A2(n3518), .ZN(MEM_stage_inst_N31) );
AND2_X1 U2665 ( .A1(ID_pipeline_reg_out_5), .A2(n3521), .ZN(EX_stage_inst_N8) );
AND2_X1 U2666 ( .A1(ID_pipeline_reg_out_6), .A2(n3521), .ZN(EX_stage_inst_N9) );
AND2_X1 U2667 ( .A1(ID_pipeline_reg_out_11), .A2(n3521), .ZN(EX_stage_inst_N14) );
AND2_X1 U2668 ( .A1(ID_pipeline_reg_out_13), .A2(n3521), .ZN(EX_stage_inst_N16) );
AND2_X1 U2669 ( .A1(ID_pipeline_reg_out_14), .A2(n3521), .ZN(EX_stage_inst_N17) );
AND2_X1 U2670 ( .A1(ID_pipeline_reg_out_17), .A2(n3521), .ZN(EX_stage_inst_N20) );
NOR2_X1 U2671 ( .A1(ID_pipeline_reg_out_29), .A2(ID_pipeline_reg_out_31), .ZN(n2366) );
NOR2_X1 U2672 ( .A1(ID_pipeline_reg_out_34), .A2(ID_pipeline_reg_out_33), .ZN(n2359) );
NOR2_X1 U2673 ( .A1(ID_pipeline_reg_out_36), .A2(ID_pipeline_reg_out_32), .ZN(n2358) );
NAND2_X1 U2674 ( .A1(n2359), .A2(n2358), .ZN(n2364) );
NOR2_X1 U2675 ( .A1(ID_pipeline_reg_out_30), .A2(ID_pipeline_reg_out_28), .ZN(n2362) );
NOR2_X1 U2676 ( .A1(ID_pipeline_reg_out_37), .A2(n2360), .ZN(n2361) );
NAND2_X1 U2677 ( .A1(n2362), .A2(n2361), .ZN(n2363) );
NOR2_X1 U2678 ( .A1(n2364), .A2(n2363), .ZN(n2365) );
NAND2_X1 U2679 ( .A1(n2366), .A2(n2365), .ZN(n2412) );
NAND2_X1 U2680 ( .A1(ID_pipeline_reg_out_55), .A2(ID_pipeline_reg_out_56), .ZN(n2367) );
NOR2_X1 U2681 ( .A1(n2412), .A2(n2367), .ZN(n2814) );
NAND2_X1 U2682 ( .A1(n2814), .A2(n3473), .ZN(n3080) );
NOR2_X1 U2683 ( .A1(rst), .A2(n3080), .ZN(n2854) );
NOR2_X1 U2684 ( .A1(n3485), .A2(n3474), .ZN(n2539) );
NAND2_X1 U2685 ( .A1(n2854), .A2(n2539), .ZN(n2417) );
NAND2_X1 U2686 ( .A1(n3488), .A2(ID_pipeline_reg_out_55), .ZN(n3026) );
NOR2_X1 U2687 ( .A1(ID_pipeline_reg_out_38), .A2(ID_pipeline_reg_out_54), .ZN(n2368) );
NOR2_X1 U2688 ( .A1(n2998), .A2(n2368), .ZN(n2369) );
NOR2_X1 U2689 ( .A1(n3472), .A2(n2369), .ZN(n2373) );
NOR2_X1 U2690 ( .A1(ID_pipeline_reg_out_22), .A2(ID_pipeline_reg_out_54), .ZN(n2370) );
NOR2_X1 U2691 ( .A1(n2998), .A2(n2370), .ZN(n2371) );
NOR2_X1 U2692 ( .A1(n3486), .A2(n2371), .ZN(n2372) );
NOR2_X1 U2693 ( .A1(n2373), .A2(n2372), .ZN(n2375) );
NOR2_X1 U2694 ( .A1(n3472), .A2(n3486), .ZN(n2419) );
OR2_X1 U2695 ( .A1(ID_pipeline_reg_out_55), .A2(n3488), .ZN(n2448) );
NAND2_X1 U2696 ( .A1(n3473), .A2(n2448), .ZN(n2548) );
NOR2_X1 U2697 ( .A1(n2419), .A2(n2548), .ZN(n2374) );
NOR2_X1 U2698 ( .A1(n2375), .A2(n2374), .ZN(n2410) );
NAND2_X1 U2699 ( .A1(n2814), .A2(n3474), .ZN(n2645) );
NAND2_X1 U2700 ( .A1(n3471), .A2(ID_pipeline_reg_out_24), .ZN(n3104) );
NOR2_X1 U2701 ( .A1(n3478), .A2(ID_pipeline_reg_out_22), .ZN(n2722) );
NAND2_X1 U2702 ( .A1(n2722), .A2(ID_pipeline_reg_out_44), .ZN(n2801) );
NOR2_X2 U2703 ( .A1(ID_pipeline_reg_out_22), .A2(ID_pipeline_reg_out_23), .ZN(n2874) );
NAND2_X1 U2704 ( .A1(n2874), .A2(ID_pipeline_reg_out_42), .ZN(n2376) );
NAND2_X1 U2705 ( .A1(n2801), .A2(n2376), .ZN(n2378) );
NOR2_X1 U2706 ( .A1(n3472), .A2(ID_pipeline_reg_out_23), .ZN(n3108) );
NAND2_X1 U2707 ( .A1(ID_pipeline_reg_out_43), .A2(n3108), .ZN(n2719) );
NAND2_X1 U2708 ( .A1(ID_pipeline_reg_out_22), .A2(ID_pipeline_reg_out_23), .ZN(n3046) );
INV_X1 U2709 ( .A(n3046), .ZN(n2943) );
NAND2_X1 U2710 ( .A1(n2943), .A2(ID_pipeline_reg_out_45), .ZN(n2878) );
NAND2_X1 U2711 ( .A1(n2719), .A2(n2878), .ZN(n2377) );
NOR2_X1 U2712 ( .A1(n2378), .A2(n2377), .ZN(n2611) );
NAND2_X1 U2713 ( .A1(n3037), .A2(n2611), .ZN(n2395) );
NAND2_X1 U2714 ( .A1(ID_pipeline_reg_out_53), .A2(ID_pipeline_reg_out_22), .ZN(n2380) );
NAND2_X1 U2715 ( .A1(ID_pipeline_reg_out_52), .A2(n3472), .ZN(n2379) );
NAND2_X1 U2716 ( .A1(n2380), .A2(n2379), .ZN(n2491) );
NAND2_X1 U2717 ( .A1(ID_pipeline_reg_out_23), .A2(n2491), .ZN(n2382) );
NAND2_X1 U2718 ( .A1(n2874), .A2(ID_pipeline_reg_out_50), .ZN(n2381) );
NAND2_X1 U2719 ( .A1(n2382), .A2(n2381), .ZN(n2384) );
NOR2_X1 U2720 ( .A1(n3045), .A2(n3483), .ZN(n2383) );
NOR2_X1 U2721 ( .A1(n2384), .A2(n2383), .ZN(n2968) );
NAND2_X1 U2722 ( .A1(ID_pipeline_reg_out_24), .A2(n2968), .ZN(n2393) );
NAND2_X1 U2723 ( .A1(ID_pipeline_reg_out_22), .A2(n3490), .ZN(n2385) );
NAND2_X1 U2724 ( .A1(n3478), .A2(n2385), .ZN(n2387) );
NOR2_X1 U2725 ( .A1(ID_pipeline_reg_out_22), .A2(ID_pipeline_reg_out_46), .ZN(n2386) );
NOR2_X1 U2726 ( .A1(n2387), .A2(n2386), .ZN(n2391) );
NAND2_X1 U2727 ( .A1(n2722), .A2(ID_pipeline_reg_out_48), .ZN(n2389) );
NAND2_X1 U2728 ( .A1(n2943), .A2(ID_pipeline_reg_out_49), .ZN(n2388) );
NAND2_X1 U2729 ( .A1(n2389), .A2(n2388), .ZN(n2390) );
NOR2_X1 U2730 ( .A1(n2391), .A2(n2390), .ZN(n2610) );
NAND2_X1 U2731 ( .A1(n2610), .A2(n3476), .ZN(n2392) );
NAND2_X1 U2732 ( .A1(n2393), .A2(n2392), .ZN(n2815) );
NAND2_X1 U2733 ( .A1(ID_pipeline_reg_out_25), .A2(n2815), .ZN(n2394) );
NAND2_X1 U2734 ( .A1(n2395), .A2(n2394), .ZN(n2396) );
NOR2_X1 U2735 ( .A1(n2645), .A2(n2396), .ZN(n2405) );
NAND2_X1 U2736 ( .A1(n3476), .A2(n3471), .ZN(n3075) );
INV_X1 U2737 ( .A(n2722), .ZN(n3041) );
NOR2_X1 U2738 ( .A1(ID_pipeline_reg_out_40), .A2(n3041), .ZN(n2400) );
NOR2_X1 U2739 ( .A1(ID_pipeline_reg_out_39), .A2(n3472), .ZN(n2525) );
NOR2_X1 U2740 ( .A1(ID_pipeline_reg_out_22), .A2(ID_pipeline_reg_out_38), .ZN(n2397) );
NOR2_X1 U2741 ( .A1(n2525), .A2(n2397), .ZN(n2398) );
NOR2_X1 U2742 ( .A1(ID_pipeline_reg_out_23), .A2(n2398), .ZN(n2399) );
NOR2_X1 U2743 ( .A1(n2400), .A2(n2399), .ZN(n2402) );
NAND2_X1 U2744 ( .A1(n2943), .A2(n3482), .ZN(n2401) );
NAND2_X1 U2745 ( .A1(n2402), .A2(n2401), .ZN(n2403) );
NAND2_X1 U2746 ( .A1(n3115), .A2(n2403), .ZN(n2404) );
NAND2_X1 U2747 ( .A1(n2405), .A2(n2404), .ZN(n2408) );
NOR2_X2 U2748 ( .A1(ID_pipeline_reg_out_55), .A2(ID_pipeline_reg_out_56), .ZN(n3098) );
XOR2_X1 U2749 ( .A(ID_pipeline_reg_out_38), .B(ID_pipeline_reg_out_22), .Z(n2406) );
NAND2_X1 U2750 ( .A1(n3098), .A2(n2406), .ZN(n2407) );
NAND2_X1 U2751 ( .A1(n2408), .A2(n2407), .ZN(n2409) );
NOR2_X1 U2752 ( .A1(n2410), .A2(n2409), .ZN(n2414) );
NAND2_X1 U2753 ( .A1(n3474), .A2(n3471), .ZN(n2812) );
OR2_X1 U2754 ( .A1(n3473), .A2(n2448), .ZN(n2411) );
OR2_X1 U2755 ( .A1(n2412), .A2(n2411), .ZN(n2806) );
NOR2_X1 U2756 ( .A1(n2812), .A2(n2806), .ZN(n2609) );
NOR2_X1 U2757 ( .A1(ID_pipeline_reg_out_24), .A2(n2772), .ZN(n2725) );
NOR2_X1 U2758 ( .A1(n3042), .A2(n3486), .ZN(n2795) );
NAND2_X1 U2759 ( .A1(n2725), .A2(n2795), .ZN(n2413) );
NAND2_X1 U2760 ( .A1(n2414), .A2(n2413), .ZN(n2415) );
NAND2_X1 U2761 ( .A1(n2415), .A2(n3518), .ZN(n2416) );
NAND2_X1 U2762 ( .A1(n2417), .A2(n2416), .ZN(EX_stage_inst_N25) );
AND2_X1 U2763 ( .A1(n3472), .A2(ID_pipeline_reg_out_39), .ZN(n2418) );
NOR2_X1 U2764 ( .A1(n2419), .A2(n2418), .ZN(n2585) );
NOR2_X1 U2765 ( .A1(ID_pipeline_reg_out_23), .A2(n2585), .ZN(n2981) );
NAND2_X1 U2766 ( .A1(n2725), .A2(n2981), .ZN(n2446) );
NOR2_X1 U2767 ( .A1(n3041), .A2(n3507), .ZN(n2828) );
NAND2_X1 U2768 ( .A1(ID_pipeline_reg_out_44), .A2(n3108), .ZN(n2421) );
NAND2_X1 U2769 ( .A1(ID_pipeline_reg_out_43), .A2(n2874), .ZN(n2420) );
NAND2_X1 U2770 ( .A1(n2421), .A2(n2420), .ZN(n2422) );
NOR2_X1 U2771 ( .A1(n2828), .A2(n2422), .ZN(n2423) );
NAND2_X1 U2772 ( .A1(n2943), .A2(ID_pipeline_reg_out_46), .ZN(n2912) );
NAND2_X1 U2773 ( .A1(n2423), .A2(n2912), .ZN(n2638) );
NOR2_X1 U2774 ( .A1(n3476), .A2(n2638), .ZN(n2431) );
NOR2_X1 U2775 ( .A1(ID_pipeline_reg_out_42), .A2(n3472), .ZN(n2654) );
NOR2_X1 U2776 ( .A1(ID_pipeline_reg_out_22), .A2(ID_pipeline_reg_out_41), .ZN(n2424) );
NOR2_X1 U2777 ( .A1(n2654), .A2(n2424), .ZN(n2425) );
NOR2_X1 U2778 ( .A1(n2425), .A2(n3478), .ZN(n2428) );
NOR2_X1 U2779 ( .A1(n3472), .A2(n3508), .ZN(n2657) );
NOR2_X1 U2780 ( .A1(ID_pipeline_reg_out_23), .A2(ID_pipeline_reg_out_39), .ZN(n2447) );
NOR2_X1 U2781 ( .A1(n3108), .A2(n2447), .ZN(n2426) );
NOR2_X1 U2782 ( .A1(n2657), .A2(n2426), .ZN(n2427) );
NOR2_X1 U2783 ( .A1(n2428), .A2(n2427), .ZN(n2429) );
NOR2_X1 U2784 ( .A1(ID_pipeline_reg_out_24), .A2(n2429), .ZN(n2430) );
NOR2_X1 U2785 ( .A1(n2431), .A2(n2430), .ZN(n2432) );
NOR2_X1 U2786 ( .A1(ID_pipeline_reg_out_25), .A2(n2432), .ZN(n2433) );
NOR2_X1 U2787 ( .A1(n2645), .A2(n2433), .ZN(n2444) );
NAND2_X1 U2788 ( .A1(n3472), .A2(n3483), .ZN(n2434) );
NAND2_X1 U2789 ( .A1(n3478), .A2(n2434), .ZN(n2436) );
NOR2_X1 U2790 ( .A1(ID_pipeline_reg_out_52), .A2(n3472), .ZN(n2435) );
NOR2_X1 U2791 ( .A1(n2436), .A2(n2435), .ZN(n2467) );
NOR2_X1 U2792 ( .A1(n3485), .A2(n3041), .ZN(n2437) );
NOR2_X1 U2793 ( .A1(n2467), .A2(n2437), .ZN(n3014) );
NAND2_X1 U2794 ( .A1(ID_pipeline_reg_out_24), .A2(n3014), .ZN(n2442) );
NAND2_X1 U2795 ( .A1(n2874), .A2(ID_pipeline_reg_out_47), .ZN(n2826) );
NAND2_X1 U2796 ( .A1(n2722), .A2(ID_pipeline_reg_out_49), .ZN(n2438) );
NAND2_X1 U2797 ( .A1(n2826), .A2(n2438), .ZN(n2440) );
NAND2_X1 U2798 ( .A1(n2943), .A2(ID_pipeline_reg_out_50), .ZN(n3112) );
NAND2_X1 U2799 ( .A1(n3108), .A2(ID_pipeline_reg_out_48), .ZN(n2913) );
NAND2_X1 U2800 ( .A1(n3112), .A2(n2913), .ZN(n2439) );
NOR2_X1 U2801 ( .A1(n2440), .A2(n2439), .ZN(n2639) );
NAND2_X1 U2802 ( .A1(n2639), .A2(n3476), .ZN(n2441) );
NAND2_X1 U2803 ( .A1(n2442), .A2(n2441), .ZN(n2846) );
NAND2_X1 U2804 ( .A1(n2846), .A2(ID_pipeline_reg_out_25), .ZN(n2443) );
NAND2_X1 U2805 ( .A1(n2444), .A2(n2443), .ZN(n2445) );
NAND2_X1 U2806 ( .A1(n2446), .A2(n2445), .ZN(n2463) );
NOR2_X2 U2807 ( .A1(ID_pipeline_reg_out_54), .A2(n2448), .ZN(n3022) );
NAND2_X1 U2808 ( .A1(ID_pipeline_reg_out_23), .A2(ID_pipeline_reg_out_39), .ZN(n2449) );
NAND2_X1 U2809 ( .A1(n3022), .A2(n2449), .ZN(n2452) );
NAND2_X1 U2810 ( .A1(n2449), .A2(n3473), .ZN(n2450) );
NAND2_X1 U2811 ( .A1(n2998), .A2(n2450), .ZN(n2451) );
NAND2_X1 U2812 ( .A1(n2452), .A2(n2451), .ZN(n2453) );
NAND2_X1 U2813 ( .A1(n2454), .A2(n2453), .ZN(n2461) );
INV_X1 U2814 ( .A(n3473), .ZN(n3093) );
XOR2_X1 U2815 ( .A(n3093), .B(ID_pipeline_reg_out_23), .Z(n2514) );
XOR2_X1 U2816 ( .A(n2514), .B(ID_pipeline_reg_out_39), .Z(n2516) );
AND2_X1 U2817 ( .A1(ID_pipeline_reg_out_38), .A2(n3093), .ZN(n2458) );
XOR2_X1 U2818 ( .A(ID_pipeline_reg_out_38), .B(n3093), .Z(n2456) );
XOR2_X1 U2819 ( .A(n3093), .B(ID_pipeline_reg_out_22), .Z(n2455) );
AND2_X1 U2820 ( .A1(n2456), .A2(n2455), .ZN(n2457) );
OR2_X1 U2821 ( .A1(n2458), .A2(n2457), .ZN(n2515) );
XOR2_X1 U2822 ( .A(n2516), .B(n2515), .Z(n2459) );
NAND2_X1 U2823 ( .A1(n3098), .A2(n2459), .ZN(n2460) );
NAND2_X1 U2824 ( .A1(n2461), .A2(n2460), .ZN(n2462) );
NOR2_X1 U2825 ( .A1(n2463), .A2(n2462), .ZN(n2464) );
NOR2_X1 U2826 ( .A1(rst), .A2(n2464), .ZN(n2474) );
NAND2_X1 U2827 ( .A1(n2539), .A2(n3476), .ZN(n2538) );
XOR2_X1 U2828 ( .A(n3474), .B(ID_pipeline_reg_out_23), .Z(n2465) );
NAND2_X1 U2829 ( .A1(n3041), .A2(n2465), .ZN(n2466) );
NAND2_X1 U2830 ( .A1(ID_pipeline_reg_out_53), .A2(n2466), .ZN(n2469) );
NAND2_X1 U2831 ( .A1(n2467), .A2(n3474), .ZN(n2468) );
NAND2_X1 U2832 ( .A1(n2469), .A2(n2468), .ZN(n2675) );
NAND2_X1 U2833 ( .A1(ID_pipeline_reg_out_24), .A2(n2675), .ZN(n2470) );
NAND2_X1 U2834 ( .A1(n2538), .A2(n2470), .ZN(n2472) );
NOR2_X1 U2835 ( .A1(ID_pipeline_reg_out_26), .A2(ID_pipeline_reg_out_24), .ZN(n2684) );
INV_X1 U2836 ( .A(n2684), .ZN(n2596) );
NOR2_X1 U2837 ( .A1(n2596), .A2(n2639), .ZN(n2471) );
NOR2_X1 U2838 ( .A1(n2472), .A2(n2471), .ZN(n2850) );
NAND2_X1 U2839 ( .A1(n2854), .A2(ID_pipeline_reg_out_25), .ZN(n2677) );
NOR2_X1 U2840 ( .A1(n2850), .A2(n2677), .ZN(n2473) );
NOR2_X1 U2841 ( .A1(n2474), .A2(n2473), .ZN(n2475) );
AND2_X1 U2842 ( .A1(n3471), .A2(n2539), .ZN(n2792) );
NAND2_X1 U2843 ( .A1(n2854), .A2(n2792), .ZN(n2680) );
NAND2_X1 U2844 ( .A1(n2475), .A2(n2680), .ZN(EX_stage_inst_N26) );
NAND2_X1 U2845 ( .A1(ID_pipeline_reg_out_24), .A2(n3474), .ZN(n2477) );
NOR2_X1 U2846 ( .A1(n2491), .A2(ID_pipeline_reg_out_23), .ZN(n2476) );
NOR2_X1 U2847 ( .A1(n2477), .A2(n2476), .ZN(n2478) );
NOR2_X1 U2848 ( .A1(n2539), .A2(n2478), .ZN(n2481) );
NOR2_X1 U2849 ( .A1(n3485), .A2(ID_pipeline_reg_out_26), .ZN(n3078) );
NAND2_X1 U2850 ( .A1(ID_pipeline_reg_out_23), .A2(n2746), .ZN(n2479) );
NOR2_X1 U2851 ( .A1(n2479), .A2(n3476), .ZN(n2480) );
NOR2_X1 U2852 ( .A1(n2481), .A2(n2480), .ZN(n2490) );
NOR2_X1 U2853 ( .A1(n3046), .A2(n3483), .ZN(n2488) );
NAND2_X1 U2854 ( .A1(ID_pipeline_reg_out_50), .A2(n2722), .ZN(n2486) );
NOR2_X1 U2855 ( .A1(ID_pipeline_reg_out_49), .A2(n3472), .ZN(n2483) );
NOR2_X1 U2856 ( .A1(ID_pipeline_reg_out_22), .A2(ID_pipeline_reg_out_48), .ZN(n2482) );
NOR2_X1 U2857 ( .A1(n2483), .A2(n2482), .ZN(n2484) );
NAND2_X1 U2858 ( .A1(n2484), .A2(n3478), .ZN(n2485) );
NAND2_X1 U2859 ( .A1(n2486), .A2(n2485), .ZN(n2487) );
NOR2_X1 U2860 ( .A1(n2488), .A2(n2487), .ZN(n2691) );
NOR2_X1 U2861 ( .A1(n2691), .A2(n2596), .ZN(n2489) );
NOR2_X1 U2862 ( .A1(n2490), .A2(n2489), .ZN(n2885) );
NOR2_X1 U2863 ( .A1(n2885), .A2(n2677), .ZN(n2536) );
NAND2_X1 U2864 ( .A1(n3478), .A2(n2491), .ZN(n3065) );
NAND2_X1 U2865 ( .A1(ID_pipeline_reg_out_24), .A2(n3065), .ZN(n2493) );
NAND2_X1 U2866 ( .A1(n2691), .A2(n3476), .ZN(n2492) );
NAND2_X1 U2867 ( .A1(n2493), .A2(n2492), .ZN(n2890) );
NAND2_X1 U2868 ( .A1(ID_pipeline_reg_out_25), .A2(n2890), .ZN(n2508) );
NOR2_X1 U2869 ( .A1(ID_pipeline_reg_out_41), .A2(n3045), .ZN(n2497) );
NOR2_X1 U2870 ( .A1(ID_pipeline_reg_out_22), .A2(ID_pipeline_reg_out_42), .ZN(n2602) );
NOR2_X1 U2871 ( .A1(ID_pipeline_reg_out_43), .A2(n3472), .ZN(n2494) );
NOR2_X1 U2872 ( .A1(n2602), .A2(n2494), .ZN(n2495) );
NOR2_X1 U2873 ( .A1(n2495), .A2(n3478), .ZN(n2496) );
NOR2_X1 U2874 ( .A1(n2497), .A2(n2496), .ZN(n2499) );
NAND2_X1 U2875 ( .A1(n2874), .A2(n3508), .ZN(n2498) );
NAND2_X1 U2876 ( .A1(n2499), .A2(n2498), .ZN(n2500) );
NAND2_X1 U2877 ( .A1(n3476), .A2(n2500), .ZN(n2505) );
NAND2_X1 U2878 ( .A1(n3108), .A2(ID_pipeline_reg_out_45), .ZN(n2800) );
NAND2_X1 U2879 ( .A1(n2943), .A2(ID_pipeline_reg_out_47), .ZN(n2501) );
NAND2_X1 U2880 ( .A1(n2800), .A2(n2501), .ZN(n2503) );
NAND2_X1 U2881 ( .A1(n2874), .A2(ID_pipeline_reg_out_44), .ZN(n2718) );
NAND2_X1 U2882 ( .A1(n2722), .A2(ID_pipeline_reg_out_46), .ZN(n2877) );
NAND2_X1 U2883 ( .A1(n2718), .A2(n2877), .ZN(n2502) );
NOR2_X1 U2884 ( .A1(n2503), .A2(n2502), .ZN(n2692) );
NAND2_X1 U2885 ( .A1(n2692), .A2(ID_pipeline_reg_out_24), .ZN(n2504) );
NAND2_X1 U2886 ( .A1(n2505), .A2(n2504), .ZN(n2506) );
NAND2_X1 U2887 ( .A1(n3471), .A2(n2506), .ZN(n2507) );
NAND2_X1 U2888 ( .A1(n2508), .A2(n2507), .ZN(n2509) );
NOR2_X1 U2889 ( .A1(n2645), .A2(n2509), .ZN(n2523) );
NAND2_X1 U2890 ( .A1(n3022), .A2(n3476), .ZN(n2512) );
NAND2_X1 U2891 ( .A1(n3476), .A2(n3473), .ZN(n2510) );
NAND2_X1 U2892 ( .A1(n2998), .A2(n2510), .ZN(n2511) );
NAND2_X1 U2893 ( .A1(n2512), .A2(n2511), .ZN(n2513) );
NAND2_X1 U2894 ( .A1(ID_pipeline_reg_out_40), .A2(n2513), .ZN(n2521) );
AND2_X1 U2895 ( .A1(n2514), .A2(ID_pipeline_reg_out_39), .ZN(n2518) );
XOR2_X1 U2896 ( .A(n3093), .B(ID_pipeline_reg_out_24), .Z(n2575) );
XOR2_X1 U2897 ( .A(n2575), .B(ID_pipeline_reg_out_40), .Z(n2576) );
XOR2_X1 U2898 ( .A(n2577), .B(n2576), .Z(n2519) );
NAND2_X1 U2899 ( .A1(n3098), .A2(n2519), .ZN(n2520) );
NAND2_X1 U2900 ( .A1(n2521), .A2(n2520), .ZN(n2522) );
NOR2_X1 U2901 ( .A1(n2523), .A2(n2522), .ZN(n2529) );
NAND2_X1 U2902 ( .A1(n2722), .A2(ID_pipeline_reg_out_38), .ZN(n2527) );
NOR2_X1 U2903 ( .A1(ID_pipeline_reg_out_22), .A2(ID_pipeline_reg_out_40), .ZN(n2524) );
NOR2_X1 U2904 ( .A1(n2525), .A2(n2524), .ZN(n2604) );
NAND2_X1 U2905 ( .A1(n2604), .A2(n3478), .ZN(n2526) );
NAND2_X1 U2906 ( .A1(n2527), .A2(n2526), .ZN(n3032) );
NAND2_X1 U2907 ( .A1(n2725), .A2(n3032), .ZN(n2528) );
NAND2_X1 U2908 ( .A1(n2529), .A2(n2528), .ZN(n2533) );
NOR2_X1 U2909 ( .A1(ID_pipeline_reg_out_40), .A2(n2976), .ZN(n2530) );
NAND2_X1 U2910 ( .A1(ID_pipeline_reg_out_54), .A2(n2998), .ZN(n3024) );
NOR2_X1 U2911 ( .A1(n2530), .A2(n2978), .ZN(n2531) );
NOR2_X1 U2912 ( .A1(n3476), .A2(n2531), .ZN(n2532) );
NOR2_X1 U2913 ( .A1(n2533), .A2(n2532), .ZN(n2534) );
NOR2_X1 U2914 ( .A1(rst), .A2(n2534), .ZN(n2535) );
NOR2_X1 U2915 ( .A1(n2536), .A2(n2535), .ZN(n2537) );
NAND2_X1 U2916 ( .A1(n2537), .A2(n2680), .ZN(EX_stage_inst_N27) );
NOR2_X1 U2917 ( .A1(n3476), .A2(n2746), .ZN(n2688) );
NOR2_X1 U2918 ( .A1(n2747), .A2(n2688), .ZN(n2595) );
NAND2_X1 U2919 ( .A1(n2539), .A2(n2874), .ZN(n3076) );
NAND2_X1 U2920 ( .A1(n2595), .A2(n3076), .ZN(n2545) );
NAND2_X1 U2921 ( .A1(ID_pipeline_reg_out_50), .A2(n3108), .ZN(n2541) );
NAND2_X1 U2922 ( .A1(ID_pipeline_reg_out_52), .A2(n2943), .ZN(n2540) );
NAND2_X1 U2923 ( .A1(n2541), .A2(n2540), .ZN(n2543) );
NAND2_X1 U2924 ( .A1(n2722), .A2(ID_pipeline_reg_out_51), .ZN(n3109) );
NAND2_X1 U2925 ( .A1(n2874), .A2(ID_pipeline_reg_out_49), .ZN(n2911) );
NAND2_X1 U2926 ( .A1(n3109), .A2(n2911), .ZN(n2542) );
NOR2_X1 U2927 ( .A1(n2543), .A2(n2542), .ZN(n2737) );
NOR2_X1 U2928 ( .A1(n2737), .A2(n2596), .ZN(n2544) );
NOR2_X1 U2929 ( .A1(n2545), .A2(n2544), .ZN(n2926) );
NOR2_X1 U2930 ( .A1(n2926), .A2(n2677), .ZN(n2546) );
NOR2_X1 U2931 ( .A1(n2546), .A2(n2600), .ZN(n2594) );
NOR2_X1 U2932 ( .A1(n3471), .A2(n3482), .ZN(n2547) );
NOR2_X1 U2933 ( .A1(n2548), .A2(n2547), .ZN(n2556) );
NOR2_X1 U2934 ( .A1(ID_pipeline_reg_out_41), .A2(ID_pipeline_reg_out_54), .ZN(n2549) );
NOR2_X1 U2935 ( .A1(n2998), .A2(n2549), .ZN(n2550) );
NOR2_X1 U2936 ( .A1(n3471), .A2(n2550), .ZN(n2554) );
NOR2_X1 U2937 ( .A1(ID_pipeline_reg_out_25), .A2(ID_pipeline_reg_out_54), .ZN(n2551) );
NOR2_X1 U2938 ( .A1(n2998), .A2(n2551), .ZN(n2552) );
NOR2_X1 U2939 ( .A1(n3482), .A2(n2552), .ZN(n2553) );
NOR2_X1 U2940 ( .A1(n2554), .A2(n2553), .ZN(n2555) );
NOR2_X1 U2941 ( .A1(n2556), .A2(n2555), .ZN(n2584) );
NOR2_X1 U2942 ( .A1(ID_pipeline_reg_out_43), .A2(n3041), .ZN(n2558) );
NOR2_X1 U2943 ( .A1(ID_pipeline_reg_out_41), .A2(n3042), .ZN(n2557) );
NOR2_X1 U2944 ( .A1(n2558), .A2(n2557), .ZN(n2562) );
NOR2_X1 U2945 ( .A1(ID_pipeline_reg_out_42), .A2(n3045), .ZN(n2560) );
NOR2_X1 U2946 ( .A1(ID_pipeline_reg_out_44), .A2(n3046), .ZN(n2559) );
NOR2_X1 U2947 ( .A1(n2560), .A2(n2559), .ZN(n2561) );
NAND2_X1 U2948 ( .A1(n2562), .A2(n2561), .ZN(n2563) );
NAND2_X1 U2949 ( .A1(n3115), .A2(n2563), .ZN(n2569) );
NAND2_X1 U2950 ( .A1(ID_pipeline_reg_out_48), .A2(n2943), .ZN(n2565) );
NAND2_X1 U2951 ( .A1(ID_pipeline_reg_out_45), .A2(n2874), .ZN(n2564) );
NAND2_X1 U2952 ( .A1(n2565), .A2(n2564), .ZN(n2567) );
NAND2_X1 U2953 ( .A1(n2722), .A2(ID_pipeline_reg_out_47), .ZN(n2910) );
NAND2_X1 U2954 ( .A1(n3108), .A2(ID_pipeline_reg_out_46), .ZN(n2825) );
NAND2_X1 U2955 ( .A1(n2910), .A2(n2825), .ZN(n2566) );
NOR2_X1 U2956 ( .A1(n2567), .A2(n2566), .ZN(n2738) );
NAND2_X1 U2957 ( .A1(n3037), .A2(n2738), .ZN(n2568) );
NAND2_X1 U2958 ( .A1(n2569), .A2(n2568), .ZN(n2570) );
NOR2_X1 U2959 ( .A1(n2645), .A2(n2570), .ZN(n2574) );
NAND2_X1 U2960 ( .A1(ID_pipeline_reg_out_53), .A2(n2874), .ZN(n3122) );
NAND2_X1 U2961 ( .A1(ID_pipeline_reg_out_24), .A2(n3122), .ZN(n2572) );
NAND2_X1 U2962 ( .A1(n2737), .A2(n3476), .ZN(n2571) );
NAND2_X1 U2963 ( .A1(n2572), .A2(n2571), .ZN(n2931) );
NAND2_X1 U2964 ( .A1(ID_pipeline_reg_out_25), .A2(n2931), .ZN(n2573) );
NAND2_X1 U2965 ( .A1(n2574), .A2(n2573), .ZN(n2582) );
AND2_X1 U2966 ( .A1(n2575), .A2(ID_pipeline_reg_out_40), .ZN(n2579) );
OR2_X1 U2967 ( .A1(n2579), .A2(n2578), .ZN(n2629) );
XOR2_X1 U2968 ( .A(n3093), .B(ID_pipeline_reg_out_25), .Z(n2627) );
XOR2_X1 U2969 ( .A(n2627), .B(ID_pipeline_reg_out_41), .Z(n2628) );
XOR2_X1 U2970 ( .A(n2629), .B(n2628), .Z(n2580) );
NAND2_X1 U2971 ( .A1(n3098), .A2(n2580), .ZN(n2581) );
NAND2_X1 U2972 ( .A1(n2582), .A2(n2581), .ZN(n2583) );
NOR2_X1 U2973 ( .A1(n2584), .A2(n2583), .ZN(n2591) );
NOR2_X1 U2974 ( .A1(n3042), .A2(n3482), .ZN(n2587) );
NOR2_X1 U2975 ( .A1(n2585), .A2(n3478), .ZN(n2586) );
NOR2_X1 U2976 ( .A1(n2587), .A2(n2586), .ZN(n2589) );
NAND2_X1 U2977 ( .A1(n2657), .A2(n3478), .ZN(n2588) );
NAND2_X1 U2978 ( .A1(n2589), .A2(n2588), .ZN(n2920) );
NAND2_X1 U2979 ( .A1(n2725), .A2(n2920), .ZN(n2590) );
NAND2_X1 U2980 ( .A1(n2591), .A2(n2590), .ZN(n2592) );
NAND2_X1 U2981 ( .A1(n2592), .A2(n3518), .ZN(n2593) );
NAND2_X1 U2982 ( .A1(n2594), .A2(n2593), .ZN(EX_stage_inst_N28) );
NOR2_X1 U2983 ( .A1(n2968), .A2(n2596), .ZN(n2597) );
NOR2_X1 U2984 ( .A1(n2598), .A2(n2597), .ZN(n2972) );
NOR2_X1 U2985 ( .A1(n2972), .A2(n2677), .ZN(n2599) );
NOR2_X1 U2986 ( .A1(n2600), .A2(n2599), .ZN(n2637) );
NOR2_X1 U2987 ( .A1(n3472), .A2(ID_pipeline_reg_out_41), .ZN(n2601) );
NOR2_X1 U2988 ( .A1(n2602), .A2(n2601), .ZN(n2603) );
NOR2_X1 U2989 ( .A1(ID_pipeline_reg_out_23), .A2(n2603), .ZN(n2606) );
NOR2_X1 U2990 ( .A1(n2604), .A2(n3478), .ZN(n2605) );
NOR2_X1 U2991 ( .A1(n2606), .A2(n2605), .ZN(n2794) );
NOR2_X1 U2992 ( .A1(ID_pipeline_reg_out_24), .A2(n2794), .ZN(n2608) );
NOR2_X1 U2993 ( .A1(n2795), .A2(n3476), .ZN(n2607) );
NOR2_X1 U2994 ( .A1(n2608), .A2(n2607), .ZN(n2935) );
NAND2_X1 U2995 ( .A1(n2609), .A2(n2935), .ZN(n2618) );
INV_X1 U2996 ( .A(n2645), .ZN(n2745) );
NOR2_X1 U2997 ( .A1(n2610), .A2(n3104), .ZN(n2613) );
NOR2_X1 U2998 ( .A1(n2611), .A2(n3075), .ZN(n2612) );
NOR2_X1 U2999 ( .A1(n2613), .A2(n2612), .ZN(n2615) );
NOR2_X1 U3000 ( .A1(n3471), .A2(ID_pipeline_reg_out_24), .ZN(n2871) );
OR2_X1 U3001 ( .A1(n3034), .A2(n2968), .ZN(n2614) );
NAND2_X1 U3002 ( .A1(n2615), .A2(n2614), .ZN(n2616) );
NAND2_X1 U3003 ( .A1(n2745), .A2(n2616), .ZN(n2617) );
NAND2_X1 U3004 ( .A1(n2618), .A2(n2617), .ZN(n2626) );
NAND2_X1 U3005 ( .A1(ID_pipeline_reg_out_26), .A2(ID_pipeline_reg_out_42), .ZN(n2620) );
NAND2_X1 U3006 ( .A1(n3022), .A2(n2620), .ZN(n2619) );
NAND2_X1 U3007 ( .A1(n3024), .A2(n2619), .ZN(n2622) );
NOR2_X1 U3008 ( .A1(n3026), .A2(n2620), .ZN(n2621) );
NOR2_X1 U3009 ( .A1(n2622), .A2(n2621), .ZN(n2624) );
NOR2_X1 U3010 ( .A1(ID_pipeline_reg_out_42), .A2(ID_pipeline_reg_out_26), .ZN(n2623) );
NOR2_X1 U3011 ( .A1(n2624), .A2(n2623), .ZN(n2625) );
NOR2_X1 U3012 ( .A1(n2626), .A2(n2625), .ZN(n2634) );
AND2_X1 U3013 ( .A1(n2627), .A2(ID_pipeline_reg_out_41), .ZN(n2631) );
AND2_X1 U3014 ( .A1(n2629), .A2(n2628), .ZN(n2630) );
XOR2_X1 U3015 ( .A(n3093), .B(ID_pipeline_reg_out_26), .Z(n2664) );
XOR2_X1 U3016 ( .A(n2664), .B(ID_pipeline_reg_out_42), .Z(n2665) );
XOR2_X1 U3017 ( .A(n2666), .B(n2665), .Z(n2632) );
NAND2_X1 U3018 ( .A1(n3098), .A2(n2632), .ZN(n2633) );
NAND2_X1 U3019 ( .A1(n2634), .A2(n2633), .ZN(n2635) );
NAND2_X1 U3020 ( .A1(n3521), .A2(n2635), .ZN(n2636) );
NAND2_X1 U3021 ( .A1(n2637), .A2(n2636), .ZN(EX_stage_inst_N29) );
NAND2_X1 U3022 ( .A1(n3115), .A2(n2638), .ZN(n2641) );
OR2_X1 U3023 ( .A1(n3104), .A2(n2639), .ZN(n2640) );
NAND2_X1 U3024 ( .A1(n2641), .A2(n2640), .ZN(n2643) );
NOR2_X1 U3025 ( .A1(n3014), .A2(n3034), .ZN(n2642) );
NOR2_X1 U3026 ( .A1(n2643), .A2(n2642), .ZN(n2644) );
NOR2_X1 U3027 ( .A1(n2645), .A2(n2644), .ZN(n2673) );
NAND2_X1 U3028 ( .A1(ID_pipeline_reg_out_27), .A2(ID_pipeline_reg_out_43), .ZN(n2647) );
NAND2_X1 U3029 ( .A1(n3022), .A2(n2647), .ZN(n2646) );
NAND2_X1 U3030 ( .A1(n3024), .A2(n2646), .ZN(n2649) );
NOR2_X1 U3031 ( .A1(n3026), .A2(n2647), .ZN(n2648) );
NOR2_X1 U3032 ( .A1(n2649), .A2(n2648), .ZN(n2651) );
NOR2_X1 U3033 ( .A1(ID_pipeline_reg_out_27), .A2(ID_pipeline_reg_out_43), .ZN(n2650) );
NOR2_X1 U3034 ( .A1(n2651), .A2(n2650), .ZN(n2663) );
NOR2_X1 U3035 ( .A1(n3476), .A2(n2772), .ZN(n2717) );
NAND2_X1 U3036 ( .A1(n2981), .A2(n2717), .ZN(n2661) );
NOR2_X1 U3037 ( .A1(n3041), .A2(n3482), .ZN(n2656) );
NAND2_X1 U3038 ( .A1(n3472), .A2(n3489), .ZN(n2652) );
NAND2_X1 U3039 ( .A1(n3478), .A2(n2652), .ZN(n2653) );
NOR2_X1 U3040 ( .A1(n2654), .A2(n2653), .ZN(n2655) );
NOR2_X1 U3041 ( .A1(n2656), .A2(n2655), .ZN(n2659) );
NAND2_X1 U3042 ( .A1(n2657), .A2(ID_pipeline_reg_out_23), .ZN(n2658) );
NAND2_X1 U3043 ( .A1(n2659), .A2(n2658), .ZN(n2993) );
NAND2_X1 U3044 ( .A1(n2725), .A2(n2993), .ZN(n2660) );
NAND2_X1 U3045 ( .A1(n2661), .A2(n2660), .ZN(n2662) );
NOR2_X1 U3046 ( .A1(n2663), .A2(n2662), .ZN(n2671) );
AND2_X1 U3047 ( .A1(n2664), .A2(ID_pipeline_reg_out_42), .ZN(n2668) );
AND2_X1 U3048 ( .A1(n2666), .A2(n2665), .ZN(n2667) );
XOR2_X1 U3049 ( .A(n3093), .B(ID_pipeline_reg_out_27), .Z(n2709) );
XOR2_X1 U3050 ( .A(n2709), .B(ID_pipeline_reg_out_43), .Z(n2710) );
XOR2_X1 U3051 ( .A(n2711), .B(n2710), .Z(n2669) );
NAND2_X1 U3052 ( .A1(n3098), .A2(n2669), .ZN(n2670) );
NAND2_X1 U3053 ( .A1(n2671), .A2(n2670), .ZN(n2672) );
NOR2_X1 U3054 ( .A1(n2673), .A2(n2672), .ZN(n2674) );
NOR2_X1 U3055 ( .A1(rst), .A2(n2674), .ZN(n2679) );
AND2_X1 U3056 ( .A1(n3476), .A2(n2675), .ZN(n2676) );
NOR2_X1 U3057 ( .A1(n2688), .A2(n2676), .ZN(n3018) );
NOR2_X1 U3058 ( .A1(n3018), .A2(n2677), .ZN(n2678) );
NOR2_X1 U3059 ( .A1(n2679), .A2(n2678), .ZN(n2681) );
NAND2_X1 U3060 ( .A1(n2681), .A2(n2680), .ZN(EX_stage_inst_N30) );
NAND2_X1 U3061 ( .A1(n2747), .A2(n3478), .ZN(n2686) );
NAND2_X1 U3062 ( .A1(ID_pipeline_reg_out_23), .A2(ID_pipeline_reg_out_53), .ZN(n2682) );
NAND2_X1 U3063 ( .A1(n3065), .A2(n2682), .ZN(n2683) );
NAND2_X1 U3064 ( .A1(n2684), .A2(n2683), .ZN(n2685) );
NAND2_X1 U3065 ( .A1(n2686), .A2(n2685), .ZN(n2687) );
NOR2_X1 U3066 ( .A1(n2688), .A2(n2687), .ZN(n3070) );
NOR2_X1 U3067 ( .A1(n3070), .A2(n3471), .ZN(n2689) );
NOR2_X1 U3068 ( .A1(n2792), .A2(n2689), .ZN(n2690) );
NOR2_X1 U3069 ( .A1(n3080), .A2(n2690), .ZN(n2708) );
NAND2_X1 U3070 ( .A1(n2691), .A2(n3037), .ZN(n2694) );
NAND2_X1 U3071 ( .A1(n2692), .A2(n3115), .ZN(n2693) );
NAND2_X1 U3072 ( .A1(n2694), .A2(n2693), .ZN(n2697) );
NOR2_X1 U3073 ( .A1(ID_pipeline_reg_out_24), .A2(n3065), .ZN(n2695) );
NOR2_X1 U3074 ( .A1(n3471), .A2(n2695), .ZN(n2696) );
NOR2_X1 U3075 ( .A1(n2697), .A2(n2696), .ZN(n2698) );
NAND2_X1 U3076 ( .A1(n2745), .A2(n2698), .ZN(n2706) );
NAND2_X1 U3077 ( .A1(ID_pipeline_reg_out_28), .A2(ID_pipeline_reg_out_44), .ZN(n2699) );
NAND2_X1 U3078 ( .A1(n3022), .A2(n2699), .ZN(n2702) );
NAND2_X1 U3079 ( .A1(n2699), .A2(n3473), .ZN(n2700) );
NAND2_X1 U3080 ( .A1(n2998), .A2(n2700), .ZN(n2701) );
NAND2_X1 U3081 ( .A1(n2702), .A2(n2701), .ZN(n2704) );
OR2_X1 U3082 ( .A1(ID_pipeline_reg_out_44), .A2(ID_pipeline_reg_out_28), .ZN(n2703) );
NAND2_X1 U3083 ( .A1(n2704), .A2(n2703), .ZN(n2705) );
NAND2_X1 U3084 ( .A1(n2706), .A2(n2705), .ZN(n2707) );
NOR2_X1 U3085 ( .A1(n2708), .A2(n2707), .ZN(n2716) );
AND2_X1 U3086 ( .A1(n2709), .A2(ID_pipeline_reg_out_43), .ZN(n2713) );
XOR2_X1 U3087 ( .A(n3093), .B(ID_pipeline_reg_out_28), .Z(n2755) );
XOR2_X1 U3088 ( .A(n2755), .B(ID_pipeline_reg_out_44), .Z(n2756) );
XOR2_X1 U3089 ( .A(n2757), .B(n2756), .Z(n2714) );
NAND2_X1 U3090 ( .A1(n3098), .A2(n2714), .ZN(n2715) );
NAND2_X1 U3091 ( .A1(n2716), .A2(n2715), .ZN(n2729) );
NAND2_X1 U3092 ( .A1(n2717), .A2(n3032), .ZN(n2727) );
NOR2_X1 U3093 ( .A1(n3482), .A2(n3046), .ZN(n2721) );
NAND2_X1 U3094 ( .A1(n2719), .A2(n2718), .ZN(n2720) );
NOR2_X1 U3095 ( .A1(n2721), .A2(n2720), .ZN(n2724) );
NAND2_X1 U3096 ( .A1(ID_pipeline_reg_out_42), .A2(n2722), .ZN(n2723) );
NAND2_X1 U3097 ( .A1(n2724), .A2(n2723), .ZN(n3033) );
NAND2_X1 U3098 ( .A1(n2725), .A2(n3033), .ZN(n2726) );
NAND2_X1 U3099 ( .A1(n2727), .A2(n2726), .ZN(n2728) );
NOR2_X1 U3100 ( .A1(n2729), .A2(n2728), .ZN(n2730) );
NOR2_X1 U3101 ( .A1(rst), .A2(n2730), .ZN(EX_stage_inst_N31) );
NAND2_X1 U3102 ( .A1(ID_pipeline_reg_out_29), .A2(ID_pipeline_reg_out_45), .ZN(n2732) );
NAND2_X1 U3103 ( .A1(n3022), .A2(n2732), .ZN(n2731) );
NAND2_X1 U3104 ( .A1(n3024), .A2(n2731), .ZN(n2734) );
NOR2_X1 U3105 ( .A1(n3026), .A2(n2732), .ZN(n2733) );
NOR2_X1 U3106 ( .A1(n2734), .A2(n2733), .ZN(n2736) );
NOR2_X1 U3107 ( .A1(ID_pipeline_reg_out_29), .A2(ID_pipeline_reg_out_45), .ZN(n2735) );
NOR2_X1 U3108 ( .A1(n2736), .A2(n2735), .ZN(n2754) );
NAND2_X1 U3109 ( .A1(n2737), .A2(n3037), .ZN(n2740) );
NAND2_X1 U3110 ( .A1(n2738), .A2(n3115), .ZN(n2739) );
NAND2_X1 U3111 ( .A1(n2740), .A2(n2739), .ZN(n2743) );
NOR2_X1 U3112 ( .A1(ID_pipeline_reg_out_24), .A2(n3122), .ZN(n2741) );
NOR2_X1 U3113 ( .A1(n3471), .A2(n2741), .ZN(n2742) );
NOR2_X1 U3114 ( .A1(n2743), .A2(n2742), .ZN(n2744) );
NAND2_X1 U3115 ( .A1(n2745), .A2(n2744), .ZN(n2752) );
NOR2_X1 U3116 ( .A1(n3471), .A2(n2746), .ZN(n2853) );
NOR2_X1 U3117 ( .A1(n2853), .A2(n2792), .ZN(n2749) );
NAND2_X1 U3118 ( .A1(n2874), .A2(n2747), .ZN(n2748) );
NAND2_X1 U3119 ( .A1(n2749), .A2(n2748), .ZN(n2750) );
NAND2_X1 U3120 ( .A1(n2884), .A2(n2750), .ZN(n2751) );
NAND2_X1 U3121 ( .A1(n2752), .A2(n2751), .ZN(n2753) );
NOR2_X1 U3122 ( .A1(n2754), .A2(n2753), .ZN(n2762) );
AND2_X1 U3123 ( .A1(n2755), .A2(ID_pipeline_reg_out_44), .ZN(n2759) );
XOR2_X1 U3124 ( .A(n3093), .B(ID_pipeline_reg_out_29), .Z(n2776) );
XOR2_X1 U3125 ( .A(n2776), .B(ID_pipeline_reg_out_45), .Z(n2777) );
XOR2_X1 U3126 ( .A(n2778), .B(n2777), .Z(n2760) );
NAND2_X1 U3127 ( .A1(n3098), .A2(n2760), .ZN(n2761) );
NAND2_X1 U3128 ( .A1(n2762), .A2(n2761), .ZN(n2774) );
OR2_X1 U3129 ( .A1(n3476), .A2(n2920), .ZN(n2771) );
NAND2_X1 U3130 ( .A1(n2943), .A2(ID_pipeline_reg_out_42), .ZN(n2767) );
NOR2_X1 U3131 ( .A1(ID_pipeline_reg_out_44), .A2(n3472), .ZN(n2763) );
NOR2_X1 U3132 ( .A1(ID_pipeline_reg_out_23), .A2(n2763), .ZN(n2765) );
NAND2_X1 U3133 ( .A1(n3507), .A2(n3472), .ZN(n2764) );
NAND2_X1 U3134 ( .A1(n2765), .A2(n2764), .ZN(n2766) );
NAND2_X1 U3135 ( .A1(n2767), .A2(n2766), .ZN(n2769) );
NOR2_X1 U3136 ( .A1(n3041), .A2(n3489), .ZN(n2768) );
NOR2_X1 U3137 ( .A1(n2769), .A2(n2768), .ZN(n2916) );
NAND2_X1 U3138 ( .A1(n2916), .A2(n3476), .ZN(n2770) );
NAND2_X1 U3139 ( .A1(n2771), .A2(n2770), .ZN(n3103) );
NOR2_X1 U3140 ( .A1(n3103), .A2(n2772), .ZN(n2773) );
NOR2_X1 U3141 ( .A1(n2774), .A2(n2773), .ZN(n2775) );
NOR2_X1 U3142 ( .A1(rst), .A2(n2775), .ZN(EX_stage_inst_N32) );
NAND2_X1 U3143 ( .A1(n2884), .A2(n2853), .ZN(n2907) );
AND2_X1 U3144 ( .A1(n2776), .A2(ID_pipeline_reg_out_45), .ZN(n2780) );
AND2_X1 U3145 ( .A1(n2778), .A2(n2777), .ZN(n2779) );
OR2_X1 U3146 ( .A1(n2780), .A2(n2779), .ZN(n2840) );
XOR2_X1 U3147 ( .A(n3093), .B(ID_pipeline_reg_out_30), .Z(n2838) );
XOR2_X1 U3148 ( .A(n2838), .B(ID_pipeline_reg_out_46), .Z(n2839) );
XOR2_X1 U3149 ( .A(n2840), .B(n2839), .Z(n2781) );
NAND2_X1 U3150 ( .A1(n3098), .A2(n2781), .ZN(n2782) );
NAND2_X1 U3151 ( .A1(n2907), .A2(n2782), .ZN(n2790) );
NAND2_X1 U3152 ( .A1(ID_pipeline_reg_out_30), .A2(ID_pipeline_reg_out_46), .ZN(n2784) );
NAND2_X1 U3153 ( .A1(n3022), .A2(n2784), .ZN(n2783) );
NAND2_X1 U3154 ( .A1(n3024), .A2(n2783), .ZN(n2786) );
NOR2_X1 U3155 ( .A1(n3026), .A2(n2784), .ZN(n2785) );
NOR2_X1 U3156 ( .A1(n2786), .A2(n2785), .ZN(n2788) );
NOR2_X1 U3157 ( .A1(ID_pipeline_reg_out_46), .A2(ID_pipeline_reg_out_30), .ZN(n2787) );
NOR2_X1 U3158 ( .A1(n2788), .A2(n2787), .ZN(n2789) );
NOR2_X1 U3159 ( .A1(n2790), .A2(n2789), .ZN(n2811) );
NOR2_X1 U3160 ( .A1(n2815), .A2(n2812), .ZN(n2791) );
NOR2_X1 U3161 ( .A1(n2792), .A2(n2791), .ZN(n2793) );
NOR2_X1 U3162 ( .A1(n3080), .A2(n2793), .ZN(n2809) );
NAND2_X1 U3163 ( .A1(n2794), .A2(n3037), .ZN(n2797) );
NAND2_X1 U3164 ( .A1(n2871), .A2(n2795), .ZN(n2796) );
NAND2_X1 U3165 ( .A1(n2797), .A2(n2796), .ZN(n2805) );
NAND2_X1 U3166 ( .A1(ID_pipeline_reg_out_43), .A2(n2943), .ZN(n2799) );
NAND2_X1 U3167 ( .A1(ID_pipeline_reg_out_46), .A2(n2874), .ZN(n2798) );
NAND2_X1 U3168 ( .A1(n2799), .A2(n2798), .ZN(n2803) );
NAND2_X1 U3169 ( .A1(n2801), .A2(n2800), .ZN(n2802) );
NOR2_X1 U3170 ( .A1(n2803), .A2(n2802), .ZN(n2938) );
NOR2_X1 U3171 ( .A1(n2938), .A2(n3075), .ZN(n2804) );
NOR2_X1 U3172 ( .A1(n2805), .A2(n2804), .ZN(n2807) );
NOR2_X1 U3173 ( .A1(n2806), .A2(ID_pipeline_reg_out_26), .ZN(n3119) );
NOR2_X1 U3174 ( .A1(n2807), .A2(n2936), .ZN(n2808) );
NOR2_X1 U3175 ( .A1(n2809), .A2(n2808), .ZN(n2810) );
NAND2_X1 U3176 ( .A1(n2811), .A2(n2810), .ZN(n2817) );
NOR2_X1 U3177 ( .A1(n3473), .A2(n2812), .ZN(n2813) );
NAND2_X1 U3178 ( .A1(n2814), .A2(n2813), .ZN(n2967) );
NOR2_X1 U3179 ( .A1(n2967), .A2(n2815), .ZN(n2816) );
NOR2_X1 U3180 ( .A1(n2817), .A2(n2816), .ZN(n2818) );
NOR2_X1 U3181 ( .A1(rst), .A2(n2818), .ZN(EX_stage_inst_N33) );
NAND2_X1 U3182 ( .A1(ID_pipeline_reg_out_31), .A2(ID_pipeline_reg_out_47), .ZN(n2820) );
NAND2_X1 U3183 ( .A1(n3022), .A2(n2820), .ZN(n2819) );
NAND2_X1 U3184 ( .A1(n3024), .A2(n2819), .ZN(n2822) );
NOR2_X1 U3185 ( .A1(n3026), .A2(n2820), .ZN(n2821) );
NOR2_X1 U3186 ( .A1(n2822), .A2(n2821), .ZN(n2824) );
NOR2_X1 U3187 ( .A1(ID_pipeline_reg_out_31), .A2(ID_pipeline_reg_out_47), .ZN(n2823) );
NOR2_X1 U3188 ( .A1(n2824), .A2(n2823), .ZN(n2837) );
NAND2_X1 U3189 ( .A1(n2826), .A2(n2825), .ZN(n2827) );
NOR2_X1 U3190 ( .A1(n2828), .A2(n2827), .ZN(n2830) );
NAND2_X1 U3191 ( .A1(ID_pipeline_reg_out_44), .A2(n2943), .ZN(n2829) );
NAND2_X1 U3192 ( .A1(n2830), .A2(n2829), .ZN(n2980) );
NAND2_X1 U3193 ( .A1(n3115), .A2(n2980), .ZN(n2832) );
NAND2_X1 U3194 ( .A1(n3037), .A2(n2993), .ZN(n2831) );
NAND2_X1 U3195 ( .A1(n2832), .A2(n2831), .ZN(n2834) );
AND2_X1 U3196 ( .A1(n2981), .A2(n2871), .ZN(n2833) );
NOR2_X1 U3197 ( .A1(n2834), .A2(n2833), .ZN(n2835) );
NOR2_X1 U3198 ( .A1(n2936), .A2(n2835), .ZN(n2836) );
NOR2_X1 U3199 ( .A1(n2837), .A2(n2836), .ZN(n2845) );
AND2_X1 U3200 ( .A1(n2838), .A2(ID_pipeline_reg_out_46), .ZN(n2842) );
XOR2_X1 U3201 ( .A(n3093), .B(ID_pipeline_reg_out_31), .Z(n2862) );
XOR2_X1 U3202 ( .A(n2862), .B(ID_pipeline_reg_out_47), .Z(n2863) );
XOR2_X1 U3203 ( .A(n2864), .B(n2863), .Z(n2843) );
NAND2_X1 U3204 ( .A1(n3098), .A2(n2843), .ZN(n2844) );
NAND2_X1 U3205 ( .A1(n2845), .A2(n2844), .ZN(n2848) );
NOR2_X1 U3206 ( .A1(n2967), .A2(n2846), .ZN(n2847) );
NOR2_X1 U3207 ( .A1(n2848), .A2(n2847), .ZN(n2849) );
NOR2_X1 U3208 ( .A1(rst), .A2(n2849), .ZN(n2852) );
NAND2_X1 U3209 ( .A1(n2854), .A2(n3471), .ZN(n3069) );
NOR2_X1 U3210 ( .A1(n2850), .A2(n3069), .ZN(n2851) );
NOR2_X1 U3211 ( .A1(n2852), .A2(n2851), .ZN(n2855) );
NAND2_X1 U3212 ( .A1(n2854), .A2(n2853), .ZN(n3073) );
NAND2_X1 U3213 ( .A1(n2855), .A2(n3073), .ZN(EX_stage_inst_N34) );
NAND2_X1 U3214 ( .A1(ID_pipeline_reg_out_32), .A2(ID_pipeline_reg_out_48), .ZN(n2857) );
NAND2_X1 U3215 ( .A1(n3022), .A2(n2857), .ZN(n2856) );
NAND2_X1 U3216 ( .A1(n3024), .A2(n2856), .ZN(n2859) );
NOR2_X1 U3217 ( .A1(n3026), .A2(n2857), .ZN(n2858) );
NOR2_X1 U3218 ( .A1(n2859), .A2(n2858), .ZN(n2861) );
NOR2_X1 U3219 ( .A1(ID_pipeline_reg_out_32), .A2(ID_pipeline_reg_out_48), .ZN(n2860) );
NOR2_X1 U3220 ( .A1(n2861), .A2(n2860), .ZN(n2870) );
AND2_X1 U3221 ( .A1(n2862), .A2(ID_pipeline_reg_out_47), .ZN(n2866) );
AND2_X1 U3222 ( .A1(n2864), .A2(n2863), .ZN(n2865) );
XOR2_X1 U3223 ( .A(n3093), .B(ID_pipeline_reg_out_32), .Z(n2900) );
XOR2_X1 U3224 ( .A(n2900), .B(ID_pipeline_reg_out_48), .Z(n2901) );
XOR2_X1 U3225 ( .A(n2902), .B(n2901), .Z(n2867) );
NAND2_X1 U3226 ( .A1(n3098), .A2(n2867), .ZN(n2868) );
NAND2_X1 U3227 ( .A1(n2907), .A2(n2868), .ZN(n2869) );
NOR2_X1 U3228 ( .A1(n2870), .A2(n2869), .ZN(n2889) );
NAND2_X1 U3229 ( .A1(n3037), .A2(n3033), .ZN(n2873) );
NAND2_X1 U3230 ( .A1(n2871), .A2(n3032), .ZN(n2872) );
NAND2_X1 U3231 ( .A1(n2873), .A2(n2872), .ZN(n2882) );
NAND2_X1 U3232 ( .A1(ID_pipeline_reg_out_47), .A2(n3108), .ZN(n2876) );
NAND2_X1 U3233 ( .A1(ID_pipeline_reg_out_48), .A2(n2874), .ZN(n2875) );
NAND2_X1 U3234 ( .A1(n2876), .A2(n2875), .ZN(n2880) );
NAND2_X1 U3235 ( .A1(n2878), .A2(n2877), .ZN(n2879) );
NOR2_X1 U3236 ( .A1(n2880), .A2(n2879), .ZN(n3038) );
NOR2_X1 U3237 ( .A1(n3038), .A2(n3075), .ZN(n2881) );
NOR2_X1 U3238 ( .A1(n2882), .A2(n2881), .ZN(n2883) );
NOR2_X1 U3239 ( .A1(n2883), .A2(n2936), .ZN(n2887) );
NAND2_X1 U3240 ( .A1(n2884), .A2(n3471), .ZN(n2925) );
NOR2_X1 U3241 ( .A1(n2885), .A2(n2925), .ZN(n2886) );
NOR2_X1 U3242 ( .A1(n2887), .A2(n2886), .ZN(n2888) );
NAND2_X1 U3243 ( .A1(n2889), .A2(n2888), .ZN(n2892) );
NOR2_X1 U3244 ( .A1(n2967), .A2(n2890), .ZN(n2891) );
NOR2_X1 U3245 ( .A1(n2892), .A2(n2891), .ZN(n2893) );
NOR2_X1 U3246 ( .A1(rst), .A2(n2893), .ZN(EX_stage_inst_N35) );
NAND2_X1 U3247 ( .A1(ID_pipeline_reg_out_33), .A2(ID_pipeline_reg_out_49), .ZN(n2895) );
NAND2_X1 U3248 ( .A1(n3022), .A2(n2895), .ZN(n2894) );
NAND2_X1 U3249 ( .A1(n3024), .A2(n2894), .ZN(n2897) );
NOR2_X1 U3250 ( .A1(n3026), .A2(n2895), .ZN(n2896) );
NOR2_X1 U3251 ( .A1(n2897), .A2(n2896), .ZN(n2899) );
NOR2_X1 U3252 ( .A1(ID_pipeline_reg_out_33), .A2(ID_pipeline_reg_out_49), .ZN(n2898) );
NOR2_X1 U3253 ( .A1(n2899), .A2(n2898), .ZN(n2909) );
AND2_X1 U3254 ( .A1(n2900), .A2(ID_pipeline_reg_out_48), .ZN(n2904) );
AND2_X1 U3255 ( .A1(n2902), .A2(n2901), .ZN(n2903) );
XOR2_X1 U3256 ( .A(n3093), .B(ID_pipeline_reg_out_33), .Z(n2959) );
XOR2_X1 U3257 ( .A(n2959), .B(ID_pipeline_reg_out_49), .Z(n2960) );
XOR2_X1 U3258 ( .A(n2961), .B(n2960), .Z(n2905) );
NAND2_X1 U3259 ( .A1(n3098), .A2(n2905), .ZN(n2906) );
NAND2_X1 U3260 ( .A1(n2907), .A2(n2906), .ZN(n2908) );
NOR2_X1 U3261 ( .A1(n2909), .A2(n2908), .ZN(n2930) );
NAND2_X1 U3262 ( .A1(n2911), .A2(n2910), .ZN(n2915) );
NAND2_X1 U3263 ( .A1(n2913), .A2(n2912), .ZN(n2914) );
NOR2_X1 U3264 ( .A1(n2915), .A2(n2914), .ZN(n3105) );
NAND2_X1 U3265 ( .A1(n3105), .A2(n3476), .ZN(n2918) );
NAND2_X1 U3266 ( .A1(n2916), .A2(ID_pipeline_reg_out_24), .ZN(n2917) );
NAND2_X1 U3267 ( .A1(n2918), .A2(n2917), .ZN(n2919) );
NAND2_X1 U3268 ( .A1(n3471), .A2(n2919), .ZN(n2923) );
NAND2_X1 U3269 ( .A1(n2920), .A2(n3476), .ZN(n2921) );
NAND2_X1 U3270 ( .A1(ID_pipeline_reg_out_25), .A2(n2921), .ZN(n2922) );
NAND2_X1 U3271 ( .A1(n2923), .A2(n2922), .ZN(n2924) );
NOR2_X1 U3272 ( .A1(n2936), .A2(n2924), .ZN(n2928) );
NOR2_X1 U3273 ( .A1(n2926), .A2(n2925), .ZN(n2927) );
NOR2_X1 U3274 ( .A1(n2928), .A2(n2927), .ZN(n2929) );
NAND2_X1 U3275 ( .A1(n2930), .A2(n2929), .ZN(n2933) );
NOR2_X1 U3276 ( .A1(n2967), .A2(n2931), .ZN(n2932) );
NOR2_X1 U3277 ( .A1(n2933), .A2(n2932), .ZN(n2934) );
NOR2_X1 U3278 ( .A1(rst), .A2(n2934), .ZN(EX_stage_inst_N36) );
NOR2_X1 U3279 ( .A1(n2935), .A2(n3471), .ZN(n2937) );
NOR2_X1 U3280 ( .A1(n2937), .A2(n2936), .ZN(n2940) );
NAND2_X1 U3281 ( .A1(n3037), .A2(n2938), .ZN(n2939) );
NAND2_X1 U3282 ( .A1(n2940), .A2(n2939), .ZN(n2950) );
NOR2_X1 U3283 ( .A1(ID_pipeline_reg_out_48), .A2(n3041), .ZN(n2942) );
NOR2_X1 U3284 ( .A1(ID_pipeline_reg_out_50), .A2(n3042), .ZN(n2941) );
NOR2_X1 U3285 ( .A1(n2942), .A2(n2941), .ZN(n2945) );
NAND2_X1 U3286 ( .A1(n2943), .A2(n3490), .ZN(n2944) );
NAND2_X1 U3287 ( .A1(n2945), .A2(n2944), .ZN(n2947) );
NOR2_X1 U3288 ( .A1(ID_pipeline_reg_out_49), .A2(n3045), .ZN(n2946) );
NOR2_X1 U3289 ( .A1(n2947), .A2(n2946), .ZN(n2948) );
NOR2_X1 U3290 ( .A1(n2948), .A2(n3075), .ZN(n2949) );
NOR2_X1 U3291 ( .A1(n2950), .A2(n2949), .ZN(n2958) );
NAND2_X1 U3292 ( .A1(ID_pipeline_reg_out_34), .A2(ID_pipeline_reg_out_50), .ZN(n2952) );
NAND2_X1 U3293 ( .A1(n3022), .A2(n2952), .ZN(n2951) );
NAND2_X1 U3294 ( .A1(n3024), .A2(n2951), .ZN(n2954) );
NOR2_X1 U3295 ( .A1(n3026), .A2(n2952), .ZN(n2953) );
NOR2_X1 U3296 ( .A1(n2954), .A2(n2953), .ZN(n2956) );
NOR2_X1 U3297 ( .A1(ID_pipeline_reg_out_34), .A2(ID_pipeline_reg_out_50), .ZN(n2955) );
NOR2_X1 U3298 ( .A1(n2956), .A2(n2955), .ZN(n2957) );
NOR2_X1 U3299 ( .A1(n2958), .A2(n2957), .ZN(n2966) );
AND2_X1 U3300 ( .A1(n2959), .A2(ID_pipeline_reg_out_49), .ZN(n2963) );
OR2_X1 U3301 ( .A1(n2963), .A2(n2962), .ZN(n3008) );
XOR2_X1 U3302 ( .A(n3093), .B(ID_pipeline_reg_out_34), .Z(n3006) );
XOR2_X1 U3303 ( .A(n3006), .B(ID_pipeline_reg_out_50), .Z(n3007) );
XOR2_X1 U3304 ( .A(n3008), .B(n3007), .Z(n2964) );
NAND2_X1 U3305 ( .A1(n3098), .A2(n2964), .ZN(n2965) );
NAND2_X1 U3306 ( .A1(n2966), .A2(n2965), .ZN(n2970) );
OR2_X1 U3307 ( .A1(n2967), .A2(ID_pipeline_reg_out_24), .ZN(n3123) );
NOR2_X1 U3308 ( .A1(n3123), .A2(n2968), .ZN(n2969) );
NOR2_X1 U3309 ( .A1(n2970), .A2(n2969), .ZN(n2971) );
NOR2_X1 U3310 ( .A1(rst), .A2(n2971), .ZN(n2974) );
NOR2_X1 U3311 ( .A1(n2972), .A2(n3069), .ZN(n2973) );
NOR2_X1 U3312 ( .A1(n2974), .A2(n2973), .ZN(n2975) );
NAND2_X1 U3313 ( .A1(n2975), .A2(n3073), .ZN(EX_stage_inst_N37) );
NOR2_X1 U3314 ( .A1(ID_pipeline_reg_out_35), .A2(n2976), .ZN(n2977) );
NOR2_X1 U3315 ( .A1(n2978), .A2(n2977), .ZN(n2979) );
NOR2_X1 U3316 ( .A1(n3483), .A2(n2979), .ZN(n3005) );
NOR2_X1 U3317 ( .A1(n3104), .A2(n2980), .ZN(n2983) );
NAND2_X1 U3318 ( .A1(ID_pipeline_reg_out_24), .A2(ID_pipeline_reg_out_25), .ZN(n3031) );
NOR2_X1 U3319 ( .A1(n2981), .A2(n3031), .ZN(n2982) );
NOR2_X1 U3320 ( .A1(n2983), .A2(n2982), .ZN(n2992) );
NOR2_X1 U3321 ( .A1(ID_pipeline_reg_out_49), .A2(n3041), .ZN(n2985) );
NOR2_X1 U3322 ( .A1(ID_pipeline_reg_out_51), .A2(n3042), .ZN(n2984) );
NOR2_X1 U3323 ( .A1(n2985), .A2(n2984), .ZN(n2989) );
NOR2_X1 U3324 ( .A1(ID_pipeline_reg_out_50), .A2(n3045), .ZN(n2987) );
NOR2_X1 U3325 ( .A1(ID_pipeline_reg_out_48), .A2(n3046), .ZN(n2986) );
NOR2_X1 U3326 ( .A1(n2987), .A2(n2986), .ZN(n2988) );
NAND2_X1 U3327 ( .A1(n2989), .A2(n2988), .ZN(n2990) );
NAND2_X1 U3328 ( .A1(n3115), .A2(n2990), .ZN(n2991) );
NAND2_X1 U3329 ( .A1(n2992), .A2(n2991), .ZN(n2995) );
NOR2_X1 U3330 ( .A1(n3034), .A2(n2993), .ZN(n2994) );
NOR2_X1 U3331 ( .A1(n2995), .A2(n2994), .ZN(n2996) );
NAND2_X1 U3332 ( .A1(n3119), .A2(n2996), .ZN(n3003) );
NAND2_X1 U3333 ( .A1(n3022), .A2(n3483), .ZN(n3000) );
NAND2_X1 U3334 ( .A1(n3483), .A2(n3473), .ZN(n2997) );
NAND2_X1 U3335 ( .A1(n2998), .A2(n2997), .ZN(n2999) );
NAND2_X1 U3336 ( .A1(n3000), .A2(n2999), .ZN(n3001) );
NAND2_X1 U3337 ( .A1(ID_pipeline_reg_out_35), .A2(n3001), .ZN(n3002) );
NAND2_X1 U3338 ( .A1(n3003), .A2(n3002), .ZN(n3004) );
NOR2_X1 U3339 ( .A1(n3005), .A2(n3004), .ZN(n3013) );
AND2_X1 U3340 ( .A1(n3006), .A2(ID_pipeline_reg_out_50), .ZN(n3010) );
OR2_X1 U3341 ( .A1(n3010), .A2(n3009), .ZN(n3059) );
XOR2_X1 U3342 ( .A(n3093), .B(ID_pipeline_reg_out_35), .Z(n3057) );
XOR2_X1 U3343 ( .A(n3057), .B(ID_pipeline_reg_out_51), .Z(n3058) );
XOR2_X1 U3344 ( .A(n3059), .B(n3058), .Z(n3011) );
NAND2_X1 U3345 ( .A1(n3098), .A2(n3011), .ZN(n3012) );
NAND2_X1 U3346 ( .A1(n3013), .A2(n3012), .ZN(n3016) );
NOR2_X1 U3347 ( .A1(n3123), .A2(n3014), .ZN(n3015) );
NOR2_X1 U3348 ( .A1(n3016), .A2(n3015), .ZN(n3017) );
NOR2_X1 U3349 ( .A1(rst), .A2(n3017), .ZN(n3020) );
NOR2_X1 U3350 ( .A1(n3018), .A2(n3069), .ZN(n3019) );
NOR2_X1 U3351 ( .A1(n3020), .A2(n3019), .ZN(n3021) );
NAND2_X1 U3352 ( .A1(n3021), .A2(n3073), .ZN(EX_stage_inst_N38) );
NAND2_X1 U3353 ( .A1(ID_pipeline_reg_out_36), .A2(ID_pipeline_reg_out_52), .ZN(n3025) );
NAND2_X1 U3354 ( .A1(n3022), .A2(n3025), .ZN(n3023) );
NAND2_X1 U3355 ( .A1(n3024), .A2(n3023), .ZN(n3028) );
NOR2_X1 U3356 ( .A1(n3026), .A2(n3025), .ZN(n3027) );
NOR2_X1 U3357 ( .A1(n3028), .A2(n3027), .ZN(n3030) );
NOR2_X1 U3358 ( .A1(ID_pipeline_reg_out_36), .A2(ID_pipeline_reg_out_52), .ZN(n3029) );
NOR2_X1 U3359 ( .A1(n3030), .A2(n3029), .ZN(n3056) );
NOR2_X1 U3360 ( .A1(n3032), .A2(n3031), .ZN(n3036) );
NOR2_X1 U3361 ( .A1(n3034), .A2(n3033), .ZN(n3035) );
NOR2_X1 U3362 ( .A1(n3036), .A2(n3035), .ZN(n3040) );
NAND2_X1 U3363 ( .A1(n3038), .A2(n3037), .ZN(n3039) );
NAND2_X1 U3364 ( .A1(n3040), .A2(n3039), .ZN(n3054) );
NOR2_X1 U3365 ( .A1(ID_pipeline_reg_out_50), .A2(n3041), .ZN(n3044) );
NOR2_X1 U3366 ( .A1(ID_pipeline_reg_out_52), .A2(n3042), .ZN(n3043) );
NOR2_X1 U3367 ( .A1(n3044), .A2(n3043), .ZN(n3050) );
NOR2_X1 U3368 ( .A1(ID_pipeline_reg_out_51), .A2(n3045), .ZN(n3048) );
NOR2_X1 U3369 ( .A1(ID_pipeline_reg_out_49), .A2(n3046), .ZN(n3047) );
NOR2_X1 U3370 ( .A1(n3048), .A2(n3047), .ZN(n3049) );
NAND2_X1 U3371 ( .A1(n3050), .A2(n3049), .ZN(n3051) );
NAND2_X1 U3372 ( .A1(n3115), .A2(n3051), .ZN(n3052) );
NAND2_X1 U3373 ( .A1(n3119), .A2(n3052), .ZN(n3053) );
NOR2_X1 U3374 ( .A1(n3054), .A2(n3053), .ZN(n3055) );
NOR2_X1 U3375 ( .A1(n3056), .A2(n3055), .ZN(n3064) );
AND2_X1 U3376 ( .A1(n3057), .A2(ID_pipeline_reg_out_51), .ZN(n3061) );
AND2_X1 U3377 ( .A1(n3059), .A2(n3058), .ZN(n3060) );
XOR2_X1 U3378 ( .A(n3093), .B(ID_pipeline_reg_out_36), .Z(n3088) );
XOR2_X1 U3379 ( .A(n3088), .B(ID_pipeline_reg_out_52), .Z(n3089) );
XOR2_X1 U3380 ( .A(n3090), .B(n3089), .Z(n3062) );
NAND2_X1 U3381 ( .A1(n3098), .A2(n3062), .ZN(n3063) );
NAND2_X1 U3382 ( .A1(n3064), .A2(n3063), .ZN(n3067) );
NOR2_X1 U3383 ( .A1(n3123), .A2(n3065), .ZN(n3066) );
NOR2_X1 U3384 ( .A1(n3067), .A2(n3066), .ZN(n3068) );
NOR2_X1 U3385 ( .A1(rst), .A2(n3068), .ZN(n3072) );
NOR2_X1 U3386 ( .A1(n3070), .A2(n3069), .ZN(n3071) );
NOR2_X1 U3387 ( .A1(n3072), .A2(n3071), .ZN(n3074) );
NAND2_X1 U3388 ( .A1(n3074), .A2(n3073), .ZN(EX_stage_inst_N39) );
NOR2_X1 U3389 ( .A1(n3076), .A2(n3075), .ZN(n3077) );
NOR2_X1 U3390 ( .A1(n3078), .A2(n3077), .ZN(n3079) );
NOR2_X1 U3391 ( .A1(n3080), .A2(n3079), .ZN(n3102) );
AND2_X1 U3392 ( .A1(ID_pipeline_reg_out_53), .A2(ID_pipeline_reg_out_37), .ZN(n3081) );
NOR2_X1 U3393 ( .A1(ID_pipeline_reg_out_54), .A2(n3081), .ZN(n3082) );
NOR2_X1 U3394 ( .A1(n3082), .A2(n3488), .ZN(n3084) );
AND2_X1 U3395 ( .A1(n3082), .A2(ID_pipeline_reg_out_55), .ZN(n3083) );
NOR2_X1 U3396 ( .A1(n3084), .A2(n3083), .ZN(n3087) );
NOR2_X1 U3397 ( .A1(ID_pipeline_reg_out_53), .A2(ID_pipeline_reg_out_37), .ZN(n3085) );
NOR2_X1 U3398 ( .A1(n3085), .A2(n3098), .ZN(n3086) );
NAND2_X1 U3399 ( .A1(n3087), .A2(n3086), .ZN(n3100) );
AND2_X1 U3400 ( .A1(n3088), .A2(ID_pipeline_reg_out_52), .ZN(n3092) );
AND2_X1 U3401 ( .A1(n3090), .A2(n3089), .ZN(n3091) );
XOR2_X1 U3402 ( .A(n3093), .B(ID_pipeline_reg_out_37), .Z(n3094) );
XOR2_X1 U3403 ( .A(n3094), .B(ID_pipeline_reg_out_53), .Z(n3095) );
XOR2_X1 U3404 ( .A(n3096), .B(n3095), .Z(n3097) );
NAND2_X1 U3405 ( .A1(n3098), .A2(n3097), .ZN(n3099) );
NAND2_X1 U3406 ( .A1(n3100), .A2(n3099), .ZN(n3101) );
NOR2_X1 U3407 ( .A1(n3102), .A2(n3101), .ZN(n3121) );
NOR2_X1 U3408 ( .A1(n3471), .A2(n3103), .ZN(n3107) );
NOR2_X1 U3409 ( .A1(n3105), .A2(n3104), .ZN(n3106) );
NOR2_X1 U3410 ( .A1(n3107), .A2(n3106), .ZN(n3117) );
AND2_X1 U3411 ( .A1(n3108), .A2(ID_pipeline_reg_out_52), .ZN(n3111) );
NAND2_X1 U3412 ( .A1(n3122), .A2(n3109), .ZN(n3110) );
NOR2_X1 U3413 ( .A1(n3111), .A2(n3110), .ZN(n3113) );
NAND2_X1 U3414 ( .A1(n3113), .A2(n3112), .ZN(n3114) );
NAND2_X1 U3415 ( .A1(n3115), .A2(n3114), .ZN(n3116) );
NAND2_X1 U3416 ( .A1(n3117), .A2(n3116), .ZN(n3118) );
NAND2_X1 U3417 ( .A1(n3119), .A2(n3118), .ZN(n3120) );
NAND2_X1 U3418 ( .A1(n3121), .A2(n3120), .ZN(n3125) );
NOR2_X1 U3419 ( .A1(n3123), .A2(n3122), .ZN(n3124) );
NOR2_X1 U3420 ( .A1(n3125), .A2(n3124), .ZN(n3126) );
NOR2_X1 U3421 ( .A1(rst), .A2(n3126), .ZN(EX_stage_inst_N40) );
AND2_X1 U3423 ( .A1(reg_write_dest_0), .A2(reg_write_en), .ZN(n3202) );
NOR2_X1 U3424 ( .A1(n3475), .A2(n3484), .ZN(n3187) );
NAND2_X1 U3425 ( .A1(n3202), .A2(n3187), .ZN(n3427) );
NAND2_X1 U3426 ( .A1(register_file_inst_reg_array_111), .A2(n3427), .ZN(n3130) );
INV_X1 U3427 ( .A(n3427), .ZN(n3430) );
NAND2_X1 U3428 ( .A1(MEM_pipeline_reg_out_20), .A2(MEM_pipeline_reg_out_0), .ZN(n3128) );
NAND2_X1 U3429 ( .A1(MEM_pipeline_reg_out_36), .A2(n3477), .ZN(n3127) );
NAND2_X1 U3430 ( .A1(n3128), .A2(n3127), .ZN(n3467) );
NAND2_X1 U3431 ( .A1(n3430), .A2(n3467), .ZN(n3129) );
NAND2_X1 U3432 ( .A1(n3130), .A2(n3129), .ZN(n1735) );
NOR2_X1 U3433 ( .A1(pc_1_), .A2(n3131), .ZN(n3150) );
NAND2_X1 U3434 ( .A1(n3167), .A2(n3143), .ZN(n3132) );
NOR2_X1 U3435 ( .A1(n3150), .A2(n3132), .ZN(n3134) );
NAND2_X1 U3436 ( .A1(reg_read_addr_1_0), .A2(n3176), .ZN(n3133) );
NAND2_X1 U3437 ( .A1(n3134), .A2(n3133), .ZN(n1721) );
NOR2_X1 U3438 ( .A1(pc_2_), .A2(n3153), .ZN(n3136) );
NAND2_X1 U3439 ( .A1(n3167), .A2(n3173), .ZN(n3135) );
NOR2_X1 U3440 ( .A1(n3136), .A2(n3135), .ZN(n3138) );
NAND2_X1 U3441 ( .A1(reg_read_addr_1_1), .A2(n3176), .ZN(n3137) );
NAND2_X1 U3442 ( .A1(n3138), .A2(n3137), .ZN(n1720) );
NOR2_X1 U3443 ( .A1(n3163), .A2(n3479), .ZN(n3139) );
NOR2_X1 U3444 ( .A1(n3140), .A2(n3139), .ZN(n3142) );
NAND2_X1 U3445 ( .A1(n3142), .A2(n3141), .ZN(n1719) );
INV_X1 U3446 ( .A(n3143), .ZN(n3158) );
AND2_X1 U3447 ( .A1(pc_0_), .A2(n3158), .ZN(n3147) );
NOR2_X1 U3448 ( .A1(n3144), .A2(pc_0_), .ZN(n3165) );
NAND2_X1 U3449 ( .A1(n3165), .A2(n3481), .ZN(n3145) );
NAND2_X1 U3450 ( .A1(n3167), .A2(n3145), .ZN(n3146) );
NOR2_X1 U3451 ( .A1(n3147), .A2(n3146), .ZN(n3149) );
NAND2_X1 U3452 ( .A1(ID_stage_inst_instruction_reg_9), .A2(n3176), .ZN(n3148) );
NAND2_X1 U3453 ( .A1(n3149), .A2(n3148), .ZN(n1718) );
NAND2_X1 U3454 ( .A1(ID_stage_inst_instruction_reg_10), .A2(n3176), .ZN(n3152) );
NAND2_X1 U3455 ( .A1(n3150), .A2(n3481), .ZN(n3151) );
NAND2_X1 U3456 ( .A1(n3152), .A2(n3151), .ZN(n3155) );
NOR2_X1 U3457 ( .A1(pc_0_), .A2(n3153), .ZN(n3154) );
NOR2_X1 U3458 ( .A1(n3155), .A2(n3154), .ZN(n3156) );
NAND2_X1 U3459 ( .A1(n3156), .A2(n3167), .ZN(n1717) );
NOR2_X1 U3460 ( .A1(pc_2_), .A2(n3173), .ZN(n3160) );
AND2_X1 U3461 ( .A1(n3165), .A2(pc_2_), .ZN(n3157) );
NOR2_X1 U3462 ( .A1(n3158), .A2(n3157), .ZN(n3172) );
NAND2_X1 U3463 ( .A1(n3172), .A2(n3167), .ZN(n3159) );
NOR2_X1 U3464 ( .A1(n3160), .A2(n3159), .ZN(n3162) );
NAND2_X1 U3465 ( .A1(ID_stage_inst_instruction_reg_11), .A2(n3176), .ZN(n3161) );
NAND2_X1 U3466 ( .A1(n3162), .A2(n3161), .ZN(n1716) );
NOR2_X1 U3467 ( .A1(n3163), .A2(n3487), .ZN(n3168) );
NAND2_X1 U3468 ( .A1(pc_1_), .A2(pc_2_), .ZN(n3164) );
NAND2_X1 U3469 ( .A1(n3165), .A2(n3164), .ZN(n3166) );
NAND2_X1 U3470 ( .A1(n3167), .A2(n3166), .ZN(n3178) );
NOR2_X1 U3471 ( .A1(n3168), .A2(n3178), .ZN(n3170) );
NAND2_X1 U3472 ( .A1(n3180), .A2(n3481), .ZN(n3169) );
NAND2_X1 U3473 ( .A1(n3170), .A2(n3169), .ZN(n1715) );
NAND2_X1 U3474 ( .A1(ID_stage_inst_instruction_reg_13), .A2(n3176), .ZN(n3171) );
NAND2_X1 U3475 ( .A1(n3172), .A2(n3171), .ZN(n1714) );
OR2_X1 U3476 ( .A1(n3481), .A2(n3173), .ZN(n3175) );
NAND2_X1 U3477 ( .A1(ID_stage_inst_instruction_reg_14), .A2(n3176), .ZN(n3174) );
NAND2_X1 U3478 ( .A1(n3175), .A2(n3174), .ZN(n1713) );
AND2_X1 U3479 ( .A1(n3176), .A2(ID_stage_inst_instruction_reg_15), .ZN(n3177) );
NOR2_X1 U3480 ( .A1(n3178), .A2(n3177), .ZN(n3182) );
NAND2_X1 U3481 ( .A1(pc_1_), .A2(n3481), .ZN(n3179) );
NAND2_X1 U3482 ( .A1(n3180), .A2(n3179), .ZN(n3181) );
NAND2_X1 U3483 ( .A1(n3182), .A2(n3181), .ZN(n1712) );
NAND2_X1 U3484 ( .A1(register_file_inst_reg_array_96), .A2(n3427), .ZN(n3186) );
NAND2_X1 U3485 ( .A1(MEM_pipeline_reg_out_0), .A2(MEM_pipeline_reg_out_5), .ZN(n3184) );
NAND2_X1 U3486 ( .A1(MEM_pipeline_reg_out_21), .A2(n3477), .ZN(n3183) );
NAND2_X1 U3487 ( .A1(n3184), .A2(n3183), .ZN(n3203) );
NAND2_X1 U3488 ( .A1(n3430), .A2(n3203), .ZN(n3185) );
NAND2_X1 U3489 ( .A1(n3186), .A2(n3185), .ZN(n1711) );
NOR2_X1 U3490 ( .A1(reg_write_dest_0), .A2(n3516), .ZN(n3198) );
NAND2_X1 U3491 ( .A1(n3187), .A2(n3198), .ZN(n3446) );
NAND2_X1 U3492 ( .A1(register_file_inst_reg_array_80), .A2(n3446), .ZN(n3189) );
NAND2_X1 U3493 ( .A1(n3447), .A2(n3203), .ZN(n3188) );
NAND2_X1 U3494 ( .A1(n3189), .A2(n3188), .ZN(n1710) );
NOR2_X1 U3495 ( .A1(reg_write_dest_1), .A2(n3475), .ZN(n3192) );
NAND2_X1 U3496 ( .A1(n3202), .A2(n3192), .ZN(n3450) );
NAND2_X1 U3497 ( .A1(register_file_inst_reg_array_64), .A2(n3450), .ZN(n3191) );
INV_X1 U3498 ( .A(n3450), .ZN(n3451) );
NAND2_X1 U3499 ( .A1(n3451), .A2(n3203), .ZN(n3190) );
NAND2_X1 U3500 ( .A1(n3191), .A2(n3190), .ZN(n1709) );
NAND2_X1 U3501 ( .A1(n3198), .A2(n3192), .ZN(n3454) );
NAND2_X1 U3502 ( .A1(register_file_inst_reg_array_48), .A2(n3454), .ZN(n3194) );
INV_X1 U3503 ( .A(n3454), .ZN(n3455) );
NAND2_X1 U3504 ( .A1(n3455), .A2(n3203), .ZN(n3193) );
NAND2_X1 U3505 ( .A1(n3194), .A2(n3193), .ZN(n1708) );
NOR2_X1 U3506 ( .A1(reg_write_dest_2), .A2(n3484), .ZN(n3197) );
NAND2_X1 U3507 ( .A1(n3202), .A2(n3197), .ZN(n3458) );
NAND2_X1 U3508 ( .A1(register_file_inst_reg_array_32), .A2(n3458), .ZN(n3196) );
INV_X1 U3509 ( .A(n3458), .ZN(n3459) );
NAND2_X1 U3510 ( .A1(n3459), .A2(n3203), .ZN(n3195) );
NAND2_X1 U3511 ( .A1(n3196), .A2(n3195), .ZN(n1707) );
NAND2_X1 U3512 ( .A1(n3198), .A2(n3197), .ZN(n3462) );
NAND2_X1 U3513 ( .A1(register_file_inst_reg_array_16), .A2(n3462), .ZN(n3200) );
INV_X1 U3514 ( .A(n3462), .ZN(n3463) );
NAND2_X1 U3515 ( .A1(n3463), .A2(n3203), .ZN(n3199) );
NAND2_X1 U3516 ( .A1(n3200), .A2(n3199), .ZN(n1706) );
NOR2_X1 U3517 ( .A1(reg_write_dest_2), .A2(reg_write_dest_1), .ZN(n3201) );
NAND2_X1 U3518 ( .A1(n3202), .A2(n3201), .ZN(n3466) );
NAND2_X1 U3519 ( .A1(register_file_inst_reg_array_0), .A2(n3466), .ZN(n3205) );
INV_X1 U3520 ( .A(n3466), .ZN(n3468) );
NAND2_X1 U3521 ( .A1(n3468), .A2(n3203), .ZN(n3204) );
NAND2_X1 U3522 ( .A1(n3205), .A2(n3204), .ZN(n1705) );
NAND2_X1 U3523 ( .A1(register_file_inst_reg_array_97), .A2(n3427), .ZN(n3209) );
NAND2_X1 U3524 ( .A1(MEM_pipeline_reg_out_0), .A2(MEM_pipeline_reg_out_6), .ZN(n3207) );
NAND2_X1 U3525 ( .A1(MEM_pipeline_reg_out_22), .A2(n3477), .ZN(n3206) );
NAND2_X1 U3526 ( .A1(n3207), .A2(n3206), .ZN(n3220) );
NAND2_X1 U3527 ( .A1(n3430), .A2(n3220), .ZN(n3208) );
NAND2_X1 U3528 ( .A1(n3209), .A2(n3208), .ZN(n1704) );
NAND2_X1 U3529 ( .A1(register_file_inst_reg_array_81), .A2(n3446), .ZN(n3211) );
NAND2_X1 U3530 ( .A1(n3447), .A2(n3220), .ZN(n3210) );
NAND2_X1 U3531 ( .A1(n3211), .A2(n3210), .ZN(n1703) );
NAND2_X1 U3532 ( .A1(register_file_inst_reg_array_65), .A2(n3450), .ZN(n3213) );
NAND2_X1 U3533 ( .A1(n3451), .A2(n3220), .ZN(n3212) );
NAND2_X1 U3534 ( .A1(n3213), .A2(n3212), .ZN(n1702) );
NAND2_X1 U3535 ( .A1(register_file_inst_reg_array_49), .A2(n3454), .ZN(n3215) );
NAND2_X1 U3536 ( .A1(n3455), .A2(n3220), .ZN(n3214) );
NAND2_X1 U3537 ( .A1(n3215), .A2(n3214), .ZN(n1701) );
NAND2_X1 U3538 ( .A1(register_file_inst_reg_array_33), .A2(n3458), .ZN(n3217) );
NAND2_X1 U3539 ( .A1(n3459), .A2(n3220), .ZN(n3216) );
NAND2_X1 U3540 ( .A1(n3217), .A2(n3216), .ZN(n1700) );
NAND2_X1 U3541 ( .A1(register_file_inst_reg_array_17), .A2(n3462), .ZN(n3219) );
NAND2_X1 U3542 ( .A1(n3463), .A2(n3220), .ZN(n3218) );
NAND2_X1 U3543 ( .A1(n3219), .A2(n3218), .ZN(n1699) );
NAND2_X1 U3544 ( .A1(register_file_inst_reg_array_1), .A2(n3466), .ZN(n3222) );
NAND2_X1 U3545 ( .A1(n3468), .A2(n3220), .ZN(n3221) );
NAND2_X1 U3546 ( .A1(n3222), .A2(n3221), .ZN(n1698) );
NAND2_X1 U3547 ( .A1(register_file_inst_reg_array_98), .A2(n3427), .ZN(n3226) );
NAND2_X1 U3548 ( .A1(MEM_pipeline_reg_out_0), .A2(MEM_pipeline_reg_out_7), .ZN(n3224) );
NAND2_X1 U3549 ( .A1(MEM_pipeline_reg_out_23), .A2(n3477), .ZN(n3223) );
NAND2_X1 U3550 ( .A1(n3224), .A2(n3223), .ZN(n3237) );
NAND2_X1 U3551 ( .A1(n3430), .A2(n3237), .ZN(n3225) );
NAND2_X1 U3552 ( .A1(n3226), .A2(n3225), .ZN(n1697) );
NAND2_X1 U3553 ( .A1(register_file_inst_reg_array_82), .A2(n3446), .ZN(n3228) );
NAND2_X1 U3554 ( .A1(n3447), .A2(n3237), .ZN(n3227) );
NAND2_X1 U3555 ( .A1(n3228), .A2(n3227), .ZN(n1696) );
NAND2_X1 U3556 ( .A1(register_file_inst_reg_array_66), .A2(n3450), .ZN(n3230) );
NAND2_X1 U3557 ( .A1(n3451), .A2(n3237), .ZN(n3229) );
NAND2_X1 U3558 ( .A1(n3230), .A2(n3229), .ZN(n1695) );
NAND2_X1 U3559 ( .A1(register_file_inst_reg_array_50), .A2(n3454), .ZN(n3232) );
NAND2_X1 U3560 ( .A1(n3455), .A2(n3237), .ZN(n3231) );
NAND2_X1 U3561 ( .A1(n3232), .A2(n3231), .ZN(n1694) );
NAND2_X1 U3562 ( .A1(register_file_inst_reg_array_34), .A2(n3458), .ZN(n3234) );
NAND2_X1 U3563 ( .A1(n3459), .A2(n3237), .ZN(n3233) );
NAND2_X1 U3564 ( .A1(n3234), .A2(n3233), .ZN(n1693) );
NAND2_X1 U3565 ( .A1(register_file_inst_reg_array_18), .A2(n3462), .ZN(n3236) );
NAND2_X1 U3566 ( .A1(n3463), .A2(n3237), .ZN(n3235) );
NAND2_X1 U3567 ( .A1(n3236), .A2(n3235), .ZN(n1692) );
NAND2_X1 U3568 ( .A1(register_file_inst_reg_array_2), .A2(n3466), .ZN(n3239) );
NAND2_X1 U3569 ( .A1(n3468), .A2(n3237), .ZN(n3238) );
NAND2_X1 U3570 ( .A1(n3239), .A2(n3238), .ZN(n1691) );
NAND2_X1 U3571 ( .A1(register_file_inst_reg_array_99), .A2(n3427), .ZN(n3243) );
NAND2_X1 U3572 ( .A1(MEM_pipeline_reg_out_0), .A2(MEM_pipeline_reg_out_8), .ZN(n3241) );
NAND2_X1 U3573 ( .A1(MEM_pipeline_reg_out_24), .A2(n3477), .ZN(n3240) );
NAND2_X1 U3574 ( .A1(n3241), .A2(n3240), .ZN(n3254) );
NAND2_X1 U3575 ( .A1(n3430), .A2(n3254), .ZN(n3242) );
NAND2_X1 U3576 ( .A1(n3243), .A2(n3242), .ZN(n1690) );
NAND2_X1 U3577 ( .A1(register_file_inst_reg_array_83), .A2(n3446), .ZN(n3245) );
NAND2_X1 U3578 ( .A1(n3447), .A2(n3254), .ZN(n3244) );
NAND2_X1 U3579 ( .A1(n3245), .A2(n3244), .ZN(n1689) );
NAND2_X1 U3580 ( .A1(register_file_inst_reg_array_67), .A2(n3450), .ZN(n3247) );
NAND2_X1 U3581 ( .A1(n3451), .A2(n3254), .ZN(n3246) );
NAND2_X1 U3582 ( .A1(n3247), .A2(n3246), .ZN(n1688) );
NAND2_X1 U3583 ( .A1(register_file_inst_reg_array_51), .A2(n3454), .ZN(n3249) );
NAND2_X1 U3584 ( .A1(n3455), .A2(n3254), .ZN(n3248) );
NAND2_X1 U3585 ( .A1(n3249), .A2(n3248), .ZN(n1687) );
NAND2_X1 U3586 ( .A1(register_file_inst_reg_array_35), .A2(n3458), .ZN(n3251) );
NAND2_X1 U3587 ( .A1(n3459), .A2(n3254), .ZN(n3250) );
NAND2_X1 U3588 ( .A1(n3251), .A2(n3250), .ZN(n1686) );
NAND2_X1 U3589 ( .A1(register_file_inst_reg_array_19), .A2(n3462), .ZN(n3253) );
NAND2_X1 U3590 ( .A1(n3463), .A2(n3254), .ZN(n3252) );
NAND2_X1 U3591 ( .A1(n3253), .A2(n3252), .ZN(n1685) );
NAND2_X1 U3592 ( .A1(register_file_inst_reg_array_3), .A2(n3466), .ZN(n3256) );
NAND2_X1 U3593 ( .A1(n3468), .A2(n3254), .ZN(n3255) );
NAND2_X1 U3594 ( .A1(n3256), .A2(n3255), .ZN(n1684) );
NAND2_X1 U3595 ( .A1(register_file_inst_reg_array_100), .A2(n3427), .ZN(n3260) );
NAND2_X1 U3596 ( .A1(MEM_pipeline_reg_out_0), .A2(MEM_pipeline_reg_out_9), .ZN(n3258) );
NAND2_X1 U3597 ( .A1(MEM_pipeline_reg_out_25), .A2(n3477), .ZN(n3257) );
NAND2_X1 U3598 ( .A1(n3258), .A2(n3257), .ZN(n3271) );
NAND2_X1 U3599 ( .A1(n3430), .A2(n3271), .ZN(n3259) );
NAND2_X1 U3600 ( .A1(n3260), .A2(n3259), .ZN(n1683) );
NAND2_X1 U3601 ( .A1(register_file_inst_reg_array_84), .A2(n3446), .ZN(n3262) );
NAND2_X1 U3602 ( .A1(n3447), .A2(n3271), .ZN(n3261) );
NAND2_X1 U3603 ( .A1(n3262), .A2(n3261), .ZN(n1682) );
NAND2_X1 U3604 ( .A1(register_file_inst_reg_array_68), .A2(n3450), .ZN(n3264) );
NAND2_X1 U3605 ( .A1(n3451), .A2(n3271), .ZN(n3263) );
NAND2_X1 U3606 ( .A1(n3264), .A2(n3263), .ZN(n1681) );
NAND2_X1 U3607 ( .A1(register_file_inst_reg_array_52), .A2(n3454), .ZN(n3266) );
NAND2_X1 U3608 ( .A1(n3455), .A2(n3271), .ZN(n3265) );
NAND2_X1 U3609 ( .A1(n3266), .A2(n3265), .ZN(n1680) );
NAND2_X1 U3610 ( .A1(register_file_inst_reg_array_36), .A2(n3458), .ZN(n3268) );
NAND2_X1 U3611 ( .A1(n3459), .A2(n3271), .ZN(n3267) );
NAND2_X1 U3612 ( .A1(n3268), .A2(n3267), .ZN(n1679) );
NAND2_X1 U3613 ( .A1(register_file_inst_reg_array_20), .A2(n3462), .ZN(n3270) );
NAND2_X1 U3614 ( .A1(n3463), .A2(n3271), .ZN(n3269) );
NAND2_X1 U3615 ( .A1(n3270), .A2(n3269), .ZN(n1678) );
NAND2_X1 U3616 ( .A1(register_file_inst_reg_array_4), .A2(n3466), .ZN(n3273) );
NAND2_X1 U3617 ( .A1(n3468), .A2(n3271), .ZN(n3272) );
NAND2_X1 U3618 ( .A1(n3273), .A2(n3272), .ZN(n1677) );
NAND2_X1 U3619 ( .A1(register_file_inst_reg_array_101), .A2(n3427), .ZN(n3277) );
NAND2_X1 U3620 ( .A1(MEM_pipeline_reg_out_0), .A2(MEM_pipeline_reg_out_10), .ZN(n3275) );
NAND2_X1 U3621 ( .A1(MEM_pipeline_reg_out_26), .A2(n3477), .ZN(n3274) );
NAND2_X1 U3622 ( .A1(n3275), .A2(n3274), .ZN(n3288) );
NAND2_X1 U3623 ( .A1(n3430), .A2(n3288), .ZN(n3276) );
NAND2_X1 U3624 ( .A1(n3277), .A2(n3276), .ZN(n1676) );
NAND2_X1 U3625 ( .A1(register_file_inst_reg_array_85), .A2(n3446), .ZN(n3279) );
NAND2_X1 U3626 ( .A1(n3447), .A2(n3288), .ZN(n3278) );
NAND2_X1 U3627 ( .A1(n3279), .A2(n3278), .ZN(n1675) );
NAND2_X1 U3628 ( .A1(register_file_inst_reg_array_69), .A2(n3450), .ZN(n3281) );
NAND2_X1 U3629 ( .A1(n3451), .A2(n3288), .ZN(n3280) );
NAND2_X1 U3630 ( .A1(n3281), .A2(n3280), .ZN(n1674) );
NAND2_X1 U3631 ( .A1(register_file_inst_reg_array_53), .A2(n3454), .ZN(n3283) );
NAND2_X1 U3632 ( .A1(n3455), .A2(n3288), .ZN(n3282) );
NAND2_X1 U3633 ( .A1(n3283), .A2(n3282), .ZN(n1673) );
NAND2_X1 U3634 ( .A1(register_file_inst_reg_array_37), .A2(n3458), .ZN(n3285) );
NAND2_X1 U3635 ( .A1(n3459), .A2(n3288), .ZN(n3284) );
NAND2_X1 U3636 ( .A1(n3285), .A2(n3284), .ZN(n1672) );
NAND2_X1 U3637 ( .A1(register_file_inst_reg_array_21), .A2(n3462), .ZN(n3287) );
NAND2_X1 U3638 ( .A1(n3463), .A2(n3288), .ZN(n3286) );
NAND2_X1 U3639 ( .A1(n3287), .A2(n3286), .ZN(n1671) );
NAND2_X1 U3640 ( .A1(register_file_inst_reg_array_5), .A2(n3466), .ZN(n3290) );
NAND2_X1 U3641 ( .A1(n3468), .A2(n3288), .ZN(n3289) );
NAND2_X1 U3642 ( .A1(n3290), .A2(n3289), .ZN(n1670) );
NAND2_X1 U3643 ( .A1(register_file_inst_reg_array_102), .A2(n3427), .ZN(n3294) );
NAND2_X1 U3644 ( .A1(MEM_pipeline_reg_out_0), .A2(MEM_pipeline_reg_out_11), .ZN(n3292) );
NAND2_X1 U3645 ( .A1(MEM_pipeline_reg_out_27), .A2(n3477), .ZN(n3291) );
NAND2_X1 U3646 ( .A1(n3292), .A2(n3291), .ZN(n3305) );
NAND2_X1 U3647 ( .A1(n3430), .A2(n3305), .ZN(n3293) );
NAND2_X1 U3648 ( .A1(n3294), .A2(n3293), .ZN(n1669) );
NAND2_X1 U3649 ( .A1(register_file_inst_reg_array_86), .A2(n3446), .ZN(n3296) );
NAND2_X1 U3650 ( .A1(n3447), .A2(n3305), .ZN(n3295) );
NAND2_X1 U3651 ( .A1(n3296), .A2(n3295), .ZN(n1668) );
NAND2_X1 U3652 ( .A1(register_file_inst_reg_array_70), .A2(n3450), .ZN(n3298) );
NAND2_X1 U3653 ( .A1(n3451), .A2(n3305), .ZN(n3297) );
NAND2_X1 U3654 ( .A1(n3298), .A2(n3297), .ZN(n1667) );
NAND2_X1 U3655 ( .A1(register_file_inst_reg_array_54), .A2(n3454), .ZN(n3300) );
NAND2_X1 U3656 ( .A1(n3455), .A2(n3305), .ZN(n3299) );
NAND2_X1 U3657 ( .A1(n3300), .A2(n3299), .ZN(n1666) );
NAND2_X1 U3658 ( .A1(register_file_inst_reg_array_38), .A2(n3458), .ZN(n3302) );
NAND2_X1 U3659 ( .A1(n3459), .A2(n3305), .ZN(n3301) );
NAND2_X1 U3660 ( .A1(n3302), .A2(n3301), .ZN(n1665) );
NAND2_X1 U3661 ( .A1(register_file_inst_reg_array_22), .A2(n3462), .ZN(n3304) );
NAND2_X1 U3662 ( .A1(n3463), .A2(n3305), .ZN(n3303) );
NAND2_X1 U3663 ( .A1(n3304), .A2(n3303), .ZN(n1664) );
NAND2_X1 U3664 ( .A1(register_file_inst_reg_array_6), .A2(n3466), .ZN(n3307) );
NAND2_X1 U3665 ( .A1(n3468), .A2(n3305), .ZN(n3306) );
NAND2_X1 U3666 ( .A1(n3307), .A2(n3306), .ZN(n1663) );
NAND2_X1 U3667 ( .A1(register_file_inst_reg_array_103), .A2(n3427), .ZN(n3311) );
NAND2_X1 U3668 ( .A1(MEM_pipeline_reg_out_0), .A2(MEM_pipeline_reg_out_12), .ZN(n3309) );
NAND2_X1 U3669 ( .A1(MEM_pipeline_reg_out_28), .A2(n3477), .ZN(n3308) );
NAND2_X1 U3670 ( .A1(n3309), .A2(n3308), .ZN(n3322) );
NAND2_X1 U3671 ( .A1(n3430), .A2(n3322), .ZN(n3310) );
NAND2_X1 U3672 ( .A1(n3311), .A2(n3310), .ZN(n1662) );
NAND2_X1 U3673 ( .A1(register_file_inst_reg_array_87), .A2(n3446), .ZN(n3313) );
NAND2_X1 U3674 ( .A1(n3447), .A2(n3322), .ZN(n3312) );
NAND2_X1 U3675 ( .A1(n3313), .A2(n3312), .ZN(n1661) );
NAND2_X1 U3676 ( .A1(register_file_inst_reg_array_71), .A2(n3450), .ZN(n3315) );
NAND2_X1 U3677 ( .A1(n3451), .A2(n3322), .ZN(n3314) );
NAND2_X1 U3678 ( .A1(n3315), .A2(n3314), .ZN(n1660) );
NAND2_X1 U3679 ( .A1(register_file_inst_reg_array_55), .A2(n3454), .ZN(n3317) );
NAND2_X1 U3680 ( .A1(n3455), .A2(n3322), .ZN(n3316) );
NAND2_X1 U3681 ( .A1(n3317), .A2(n3316), .ZN(n1659) );
NAND2_X1 U3682 ( .A1(register_file_inst_reg_array_39), .A2(n3458), .ZN(n3319) );
NAND2_X1 U3683 ( .A1(n3459), .A2(n3322), .ZN(n3318) );
NAND2_X1 U3684 ( .A1(n3319), .A2(n3318), .ZN(n1658) );
NAND2_X1 U3685 ( .A1(register_file_inst_reg_array_23), .A2(n3462), .ZN(n3321) );
NAND2_X1 U3686 ( .A1(n3463), .A2(n3322), .ZN(n3320) );
NAND2_X1 U3687 ( .A1(n3321), .A2(n3320), .ZN(n1657) );
NAND2_X1 U3688 ( .A1(register_file_inst_reg_array_7), .A2(n3466), .ZN(n3324) );
NAND2_X1 U3689 ( .A1(n3468), .A2(n3322), .ZN(n3323) );
NAND2_X1 U3690 ( .A1(n3324), .A2(n3323), .ZN(n1656) );
NAND2_X1 U3691 ( .A1(register_file_inst_reg_array_104), .A2(n3427), .ZN(n3328) );
NAND2_X1 U3692 ( .A1(MEM_pipeline_reg_out_0), .A2(MEM_pipeline_reg_out_13), .ZN(n3326) );
NAND2_X1 U3693 ( .A1(MEM_pipeline_reg_out_29), .A2(n3477), .ZN(n3325) );
NAND2_X1 U3694 ( .A1(n3326), .A2(n3325), .ZN(n3339) );
NAND2_X1 U3695 ( .A1(n3430), .A2(n3339), .ZN(n3327) );
NAND2_X1 U3696 ( .A1(n3328), .A2(n3327), .ZN(n1655) );
NAND2_X1 U3697 ( .A1(register_file_inst_reg_array_88), .A2(n3446), .ZN(n3330) );
NAND2_X1 U3698 ( .A1(n3447), .A2(n3339), .ZN(n3329) );
NAND2_X1 U3699 ( .A1(n3330), .A2(n3329), .ZN(n1654) );
NAND2_X1 U3700 ( .A1(register_file_inst_reg_array_72), .A2(n3450), .ZN(n3332) );
NAND2_X1 U3701 ( .A1(n3451), .A2(n3339), .ZN(n3331) );
NAND2_X1 U3702 ( .A1(n3332), .A2(n3331), .ZN(n1653) );
NAND2_X1 U3703 ( .A1(register_file_inst_reg_array_56), .A2(n3454), .ZN(n3334) );
NAND2_X1 U3704 ( .A1(n3455), .A2(n3339), .ZN(n3333) );
NAND2_X1 U3705 ( .A1(n3334), .A2(n3333), .ZN(n1652) );
NAND2_X1 U3706 ( .A1(register_file_inst_reg_array_40), .A2(n3458), .ZN(n3336) );
NAND2_X1 U3707 ( .A1(n3459), .A2(n3339), .ZN(n3335) );
NAND2_X1 U3708 ( .A1(n3336), .A2(n3335), .ZN(n1651) );
NAND2_X1 U3709 ( .A1(register_file_inst_reg_array_24), .A2(n3462), .ZN(n3338) );
NAND2_X1 U3710 ( .A1(n3463), .A2(n3339), .ZN(n3337) );
NAND2_X1 U3711 ( .A1(n3338), .A2(n3337), .ZN(n1650) );
NAND2_X1 U3712 ( .A1(register_file_inst_reg_array_8), .A2(n3466), .ZN(n3341) );
NAND2_X1 U3713 ( .A1(n3468), .A2(n3339), .ZN(n3340) );
NAND2_X1 U3714 ( .A1(n3341), .A2(n3340), .ZN(n1649) );
NAND2_X1 U3715 ( .A1(register_file_inst_reg_array_105), .A2(n3427), .ZN(n3345) );
NAND2_X1 U3716 ( .A1(MEM_pipeline_reg_out_0), .A2(MEM_pipeline_reg_out_14), .ZN(n3343) );
NAND2_X1 U3717 ( .A1(MEM_pipeline_reg_out_30), .A2(n3477), .ZN(n3342) );
NAND2_X1 U3718 ( .A1(n3343), .A2(n3342), .ZN(n3356) );
NAND2_X1 U3719 ( .A1(n3430), .A2(n3356), .ZN(n3344) );
NAND2_X1 U3720 ( .A1(n3345), .A2(n3344), .ZN(n1648) );
NAND2_X1 U3721 ( .A1(register_file_inst_reg_array_89), .A2(n3446), .ZN(n3347) );
NAND2_X1 U3722 ( .A1(n3447), .A2(n3356), .ZN(n3346) );
NAND2_X1 U3723 ( .A1(n3347), .A2(n3346), .ZN(n1647) );
NAND2_X1 U3724 ( .A1(register_file_inst_reg_array_73), .A2(n3450), .ZN(n3349) );
NAND2_X1 U3725 ( .A1(n3451), .A2(n3356), .ZN(n3348) );
NAND2_X1 U3726 ( .A1(n3349), .A2(n3348), .ZN(n1646) );
NAND2_X1 U3727 ( .A1(register_file_inst_reg_array_57), .A2(n3454), .ZN(n3351) );
NAND2_X1 U3728 ( .A1(n3455), .A2(n3356), .ZN(n3350) );
NAND2_X1 U3729 ( .A1(n3351), .A2(n3350), .ZN(n1645) );
NAND2_X1 U3730 ( .A1(register_file_inst_reg_array_41), .A2(n3458), .ZN(n3353) );
NAND2_X1 U3731 ( .A1(n3459), .A2(n3356), .ZN(n3352) );
NAND2_X1 U3732 ( .A1(n3353), .A2(n3352), .ZN(n1644) );
NAND2_X1 U3733 ( .A1(register_file_inst_reg_array_25), .A2(n3462), .ZN(n3355) );
NAND2_X1 U3734 ( .A1(n3463), .A2(n3356), .ZN(n3354) );
NAND2_X1 U3735 ( .A1(n3355), .A2(n3354), .ZN(n1643) );
NAND2_X1 U3736 ( .A1(register_file_inst_reg_array_9), .A2(n3466), .ZN(n3358) );
NAND2_X1 U3737 ( .A1(n3468), .A2(n3356), .ZN(n3357) );
NAND2_X1 U3738 ( .A1(n3358), .A2(n3357), .ZN(n1642) );
NAND2_X1 U3739 ( .A1(register_file_inst_reg_array_106), .A2(n3427), .ZN(n3362) );
NAND2_X1 U3740 ( .A1(MEM_pipeline_reg_out_0), .A2(MEM_pipeline_reg_out_15), .ZN(n3360) );
NAND2_X1 U3741 ( .A1(MEM_pipeline_reg_out_31), .A2(n3477), .ZN(n3359) );
NAND2_X1 U3742 ( .A1(n3360), .A2(n3359), .ZN(n3373) );
NAND2_X1 U3743 ( .A1(n3430), .A2(n3373), .ZN(n3361) );
NAND2_X1 U3744 ( .A1(n3362), .A2(n3361), .ZN(n1641) );
NAND2_X1 U3745 ( .A1(register_file_inst_reg_array_90), .A2(n3446), .ZN(n3364) );
NAND2_X1 U3746 ( .A1(n3447), .A2(n3373), .ZN(n3363) );
NAND2_X1 U3747 ( .A1(n3364), .A2(n3363), .ZN(n1640) );
NAND2_X1 U3748 ( .A1(register_file_inst_reg_array_74), .A2(n3450), .ZN(n3366) );
NAND2_X1 U3749 ( .A1(n3451), .A2(n3373), .ZN(n3365) );
NAND2_X1 U3750 ( .A1(n3366), .A2(n3365), .ZN(n1639) );
NAND2_X1 U3751 ( .A1(register_file_inst_reg_array_58), .A2(n3454), .ZN(n3368) );
NAND2_X1 U3752 ( .A1(n3455), .A2(n3373), .ZN(n3367) );
NAND2_X1 U3753 ( .A1(n3368), .A2(n3367), .ZN(n1638) );
NAND2_X1 U3754 ( .A1(register_file_inst_reg_array_42), .A2(n3458), .ZN(n3370) );
NAND2_X1 U3755 ( .A1(n3459), .A2(n3373), .ZN(n3369) );
NAND2_X1 U3756 ( .A1(n3370), .A2(n3369), .ZN(n1637) );
NAND2_X1 U3757 ( .A1(register_file_inst_reg_array_26), .A2(n3462), .ZN(n3372) );
NAND2_X1 U3758 ( .A1(n3463), .A2(n3373), .ZN(n3371) );
NAND2_X1 U3759 ( .A1(n3372), .A2(n3371), .ZN(n1636) );
NAND2_X1 U3760 ( .A1(register_file_inst_reg_array_10), .A2(n3466), .ZN(n3375) );
NAND2_X1 U3761 ( .A1(n3468), .A2(n3373), .ZN(n3374) );
NAND2_X1 U3762 ( .A1(n3375), .A2(n3374), .ZN(n1635) );
NAND2_X1 U3763 ( .A1(register_file_inst_reg_array_107), .A2(n3427), .ZN(n3379) );
NAND2_X1 U3764 ( .A1(MEM_pipeline_reg_out_0), .A2(MEM_pipeline_reg_out_16), .ZN(n3377) );
NAND2_X1 U3765 ( .A1(MEM_pipeline_reg_out_32), .A2(n3477), .ZN(n3376) );
NAND2_X1 U3766 ( .A1(n3377), .A2(n3376), .ZN(n3390) );
NAND2_X1 U3767 ( .A1(n3430), .A2(n3390), .ZN(n3378) );
NAND2_X1 U3768 ( .A1(n3379), .A2(n3378), .ZN(n1634) );
NAND2_X1 U3769 ( .A1(register_file_inst_reg_array_91), .A2(n3446), .ZN(n3381) );
NAND2_X1 U3770 ( .A1(n3447), .A2(n3390), .ZN(n3380) );
NAND2_X1 U3771 ( .A1(n3381), .A2(n3380), .ZN(n1633) );
NAND2_X1 U3772 ( .A1(register_file_inst_reg_array_75), .A2(n3450), .ZN(n3383) );
NAND2_X1 U3773 ( .A1(n3451), .A2(n3390), .ZN(n3382) );
NAND2_X1 U3774 ( .A1(n3383), .A2(n3382), .ZN(n1632) );
NAND2_X1 U3775 ( .A1(register_file_inst_reg_array_59), .A2(n3454), .ZN(n3385) );
NAND2_X1 U3776 ( .A1(n3455), .A2(n3390), .ZN(n3384) );
NAND2_X1 U3777 ( .A1(n3385), .A2(n3384), .ZN(n1631) );
NAND2_X1 U3778 ( .A1(register_file_inst_reg_array_43), .A2(n3458), .ZN(n3387) );
NAND2_X1 U3779 ( .A1(n3459), .A2(n3390), .ZN(n3386) );
NAND2_X1 U3780 ( .A1(n3387), .A2(n3386), .ZN(n1630) );
NAND2_X1 U3781 ( .A1(register_file_inst_reg_array_27), .A2(n3462), .ZN(n3389) );
NAND2_X1 U3782 ( .A1(n3463), .A2(n3390), .ZN(n3388) );
NAND2_X1 U3783 ( .A1(n3389), .A2(n3388), .ZN(n1629) );
NAND2_X1 U3784 ( .A1(register_file_inst_reg_array_11), .A2(n3466), .ZN(n3392) );
NAND2_X1 U3785 ( .A1(n3468), .A2(n3390), .ZN(n3391) );
NAND2_X1 U3786 ( .A1(n3392), .A2(n3391), .ZN(n1628) );
NAND2_X1 U3787 ( .A1(register_file_inst_reg_array_108), .A2(n3427), .ZN(n3396) );
NAND2_X1 U3788 ( .A1(MEM_pipeline_reg_out_0), .A2(MEM_pipeline_reg_out_17), .ZN(n3394) );
NAND2_X1 U3789 ( .A1(MEM_pipeline_reg_out_33), .A2(n3477), .ZN(n3393) );
NAND2_X1 U3790 ( .A1(n3394), .A2(n3393), .ZN(n3407) );
NAND2_X1 U3791 ( .A1(n3430), .A2(n3407), .ZN(n3395) );
NAND2_X1 U3792 ( .A1(n3396), .A2(n3395), .ZN(n1627) );
NAND2_X1 U3793 ( .A1(register_file_inst_reg_array_92), .A2(n3446), .ZN(n3398) );
NAND2_X1 U3794 ( .A1(n3447), .A2(n3407), .ZN(n3397) );
NAND2_X1 U3795 ( .A1(n3398), .A2(n3397), .ZN(n1626) );
NAND2_X1 U3796 ( .A1(register_file_inst_reg_array_76), .A2(n3450), .ZN(n3400) );
NAND2_X1 U3797 ( .A1(n3451), .A2(n3407), .ZN(n3399) );
NAND2_X1 U3798 ( .A1(n3400), .A2(n3399), .ZN(n1625) );
NAND2_X1 U3799 ( .A1(register_file_inst_reg_array_60), .A2(n3454), .ZN(n3402) );
NAND2_X1 U3800 ( .A1(n3455), .A2(n3407), .ZN(n3401) );
NAND2_X1 U3801 ( .A1(n3402), .A2(n3401), .ZN(n1624) );
NAND2_X1 U3802 ( .A1(register_file_inst_reg_array_44), .A2(n3458), .ZN(n3404) );
NAND2_X1 U3803 ( .A1(n3459), .A2(n3407), .ZN(n3403) );
NAND2_X1 U3804 ( .A1(n3404), .A2(n3403), .ZN(n1623) );
NAND2_X1 U3805 ( .A1(register_file_inst_reg_array_28), .A2(n3462), .ZN(n3406) );
NAND2_X1 U3806 ( .A1(n3463), .A2(n3407), .ZN(n3405) );
NAND2_X1 U3807 ( .A1(n3406), .A2(n3405), .ZN(n1622) );
NAND2_X1 U3808 ( .A1(register_file_inst_reg_array_12), .A2(n3466), .ZN(n3409) );
NAND2_X1 U3809 ( .A1(n3468), .A2(n3407), .ZN(n3408) );
NAND2_X1 U3810 ( .A1(n3409), .A2(n3408), .ZN(n1621) );
NAND2_X1 U3811 ( .A1(register_file_inst_reg_array_109), .A2(n3427), .ZN(n3413) );
NAND2_X1 U3812 ( .A1(MEM_pipeline_reg_out_0), .A2(MEM_pipeline_reg_out_18), .ZN(n3411) );
NAND2_X1 U3813 ( .A1(MEM_pipeline_reg_out_34), .A2(n3477), .ZN(n3410) );
NAND2_X1 U3814 ( .A1(n3411), .A2(n3410), .ZN(n3424) );
NAND2_X1 U3815 ( .A1(n3430), .A2(n3424), .ZN(n3412) );
NAND2_X1 U3816 ( .A1(n3413), .A2(n3412), .ZN(n1620) );
NAND2_X1 U3817 ( .A1(register_file_inst_reg_array_93), .A2(n3446), .ZN(n3415) );
NAND2_X1 U3818 ( .A1(n3447), .A2(n3424), .ZN(n3414) );
NAND2_X1 U3819 ( .A1(n3415), .A2(n3414), .ZN(n1619) );
NAND2_X1 U3820 ( .A1(register_file_inst_reg_array_77), .A2(n3450), .ZN(n3417) );
NAND2_X1 U3821 ( .A1(n3451), .A2(n3424), .ZN(n3416) );
NAND2_X1 U3822 ( .A1(n3417), .A2(n3416), .ZN(n1618) );
NAND2_X1 U3823 ( .A1(register_file_inst_reg_array_61), .A2(n3454), .ZN(n3419) );
NAND2_X1 U3824 ( .A1(n3455), .A2(n3424), .ZN(n3418) );
NAND2_X1 U3825 ( .A1(n3419), .A2(n3418), .ZN(n1617) );
NAND2_X1 U3826 ( .A1(register_file_inst_reg_array_45), .A2(n3458), .ZN(n3421) );
NAND2_X1 U3827 ( .A1(n3459), .A2(n3424), .ZN(n3420) );
NAND2_X1 U3828 ( .A1(n3421), .A2(n3420), .ZN(n1616) );
NAND2_X1 U3829 ( .A1(register_file_inst_reg_array_29), .A2(n3462), .ZN(n3423) );
NAND2_X1 U3830 ( .A1(n3463), .A2(n3424), .ZN(n3422) );
NAND2_X1 U3831 ( .A1(n3423), .A2(n3422), .ZN(n1615) );
NAND2_X1 U3832 ( .A1(register_file_inst_reg_array_13), .A2(n3466), .ZN(n3426) );
NAND2_X1 U3833 ( .A1(n3468), .A2(n3424), .ZN(n3425) );
NAND2_X1 U3834 ( .A1(n3426), .A2(n3425), .ZN(n1614) );
NAND2_X1 U3835 ( .A1(register_file_inst_reg_array_110), .A2(n3427), .ZN(n3432) );
NAND2_X1 U3836 ( .A1(MEM_pipeline_reg_out_0), .A2(MEM_pipeline_reg_out_19), .ZN(n3429) );
NAND2_X1 U3837 ( .A1(MEM_pipeline_reg_out_35), .A2(n3477), .ZN(n3428) );
NAND2_X1 U3838 ( .A1(n3429), .A2(n3428), .ZN(n3443) );
NAND2_X1 U3839 ( .A1(n3430), .A2(n3443), .ZN(n3431) );
NAND2_X1 U3840 ( .A1(n3432), .A2(n3431), .ZN(n1613) );
NAND2_X1 U3841 ( .A1(register_file_inst_reg_array_94), .A2(n3446), .ZN(n3434) );
NAND2_X1 U3842 ( .A1(n3447), .A2(n3443), .ZN(n3433) );
NAND2_X1 U3843 ( .A1(n3434), .A2(n3433), .ZN(n1612) );
NAND2_X1 U3844 ( .A1(register_file_inst_reg_array_78), .A2(n3450), .ZN(n3436) );
NAND2_X1 U3845 ( .A1(n3451), .A2(n3443), .ZN(n3435) );
NAND2_X1 U3846 ( .A1(n3436), .A2(n3435), .ZN(n1611) );
NAND2_X1 U3847 ( .A1(register_file_inst_reg_array_62), .A2(n3454), .ZN(n3438) );
NAND2_X1 U3848 ( .A1(n3455), .A2(n3443), .ZN(n3437) );
NAND2_X1 U3849 ( .A1(n3438), .A2(n3437), .ZN(n1610) );
NAND2_X1 U3850 ( .A1(register_file_inst_reg_array_46), .A2(n3458), .ZN(n3440) );
NAND2_X1 U3851 ( .A1(n3459), .A2(n3443), .ZN(n3439) );
NAND2_X1 U3852 ( .A1(n3440), .A2(n3439), .ZN(n1609) );
NAND2_X1 U3853 ( .A1(register_file_inst_reg_array_30), .A2(n3462), .ZN(n3442) );
NAND2_X1 U3854 ( .A1(n3463), .A2(n3443), .ZN(n3441) );
NAND2_X1 U3855 ( .A1(n3442), .A2(n3441), .ZN(n1608) );
NAND2_X1 U3856 ( .A1(register_file_inst_reg_array_14), .A2(n3466), .ZN(n3445) );
NAND2_X1 U3857 ( .A1(n3468), .A2(n3443), .ZN(n3444) );
NAND2_X1 U3858 ( .A1(n3445), .A2(n3444), .ZN(n1607) );
NAND2_X1 U3859 ( .A1(register_file_inst_reg_array_95), .A2(n3446), .ZN(n3449) );
NAND2_X1 U3860 ( .A1(n3447), .A2(n3467), .ZN(n3448) );
NAND2_X1 U3861 ( .A1(n3449), .A2(n3448), .ZN(n1606) );
NAND2_X1 U3862 ( .A1(register_file_inst_reg_array_79), .A2(n3450), .ZN(n3453) );
NAND2_X1 U3863 ( .A1(n3451), .A2(n3467), .ZN(n3452) );
NAND2_X1 U3864 ( .A1(n3453), .A2(n3452), .ZN(n1605) );
NAND2_X1 U3865 ( .A1(register_file_inst_reg_array_63), .A2(n3454), .ZN(n3457) );
NAND2_X1 U3866 ( .A1(n3455), .A2(n3467), .ZN(n3456) );
NAND2_X1 U3867 ( .A1(n3457), .A2(n3456), .ZN(n1604) );
NAND2_X1 U3868 ( .A1(register_file_inst_reg_array_47), .A2(n3458), .ZN(n3461) );
NAND2_X1 U3869 ( .A1(n3459), .A2(n3467), .ZN(n3460) );
NAND2_X1 U3870 ( .A1(n3461), .A2(n3460), .ZN(n1603) );
NAND2_X1 U3871 ( .A1(register_file_inst_reg_array_31), .A2(n3462), .ZN(n3465) );
NAND2_X1 U3872 ( .A1(n3463), .A2(n3467), .ZN(n3464) );
NAND2_X1 U3873 ( .A1(n3465), .A2(n3464), .ZN(n1602) );
NAND2_X1 U3874 ( .A1(register_file_inst_reg_array_15), .A2(n3466), .ZN(n3470) );
NAND2_X1 U3875 ( .A1(n3468), .A2(n3467), .ZN(n3469) );
NAND2_X1 U3876 ( .A1(n3470), .A2(n3469), .ZN(n1601) );
BUF_X1 MEM_stage_inst_dmem_U8713 ( .A(clk), .Z(MEM_stage_inst_dmem_n21637) );
BUF_X1 MEM_stage_inst_dmem_U265 ( .A(clk), .Z(MEM_stage_inst_dmem_n21636) );
BUF_X1 MEM_stage_inst_dmem_U263 ( .A(clk), .Z(MEM_stage_inst_dmem_n21635) );
BUF_X1 MEM_stage_inst_dmem_U244 ( .A(clk), .Z(MEM_stage_inst_dmem_n21634) );
BUF_X1 MEM_stage_inst_dmem_U243 ( .A(MEM_stage_inst_dmem_n21618), .Z(MEM_stage_inst_dmem_n21633) );
BUF_X1 MEM_stage_inst_dmem_U242 ( .A(MEM_stage_inst_dmem_n21634), .Z(MEM_stage_inst_dmem_n21632) );
BUF_X1 MEM_stage_inst_dmem_U241 ( .A(MEM_stage_inst_dmem_n21634), .Z(MEM_stage_inst_dmem_n21631) );
BUF_X1 MEM_stage_inst_dmem_U240 ( .A(MEM_stage_inst_dmem_n21634), .Z(MEM_stage_inst_dmem_n21630) );
BUF_X1 MEM_stage_inst_dmem_U239 ( .A(MEM_stage_inst_dmem_n21634), .Z(MEM_stage_inst_dmem_n21629) );
BUF_X1 MEM_stage_inst_dmem_U238 ( .A(MEM_stage_inst_dmem_n21634), .Z(MEM_stage_inst_dmem_n21628) );
BUF_X1 MEM_stage_inst_dmem_U237 ( .A(MEM_stage_inst_dmem_n21635), .Z(MEM_stage_inst_dmem_n21627) );
BUF_X1 MEM_stage_inst_dmem_U236 ( .A(MEM_stage_inst_dmem_n21635), .Z(MEM_stage_inst_dmem_n21626) );
BUF_X1 MEM_stage_inst_dmem_U235 ( .A(MEM_stage_inst_dmem_n21635), .Z(MEM_stage_inst_dmem_n21625) );
BUF_X1 MEM_stage_inst_dmem_U234 ( .A(MEM_stage_inst_dmem_n21635), .Z(MEM_stage_inst_dmem_n21624) );
BUF_X1 MEM_stage_inst_dmem_U233 ( .A(MEM_stage_inst_dmem_n21635), .Z(MEM_stage_inst_dmem_n21623) );
BUF_X1 MEM_stage_inst_dmem_U232 ( .A(MEM_stage_inst_dmem_n21636), .Z(MEM_stage_inst_dmem_n21622) );
BUF_X1 MEM_stage_inst_dmem_U231 ( .A(MEM_stage_inst_dmem_n21636), .Z(MEM_stage_inst_dmem_n21621) );
BUF_X1 MEM_stage_inst_dmem_U230 ( .A(MEM_stage_inst_dmem_n21636), .Z(MEM_stage_inst_dmem_n21620) );
BUF_X1 MEM_stage_inst_dmem_U229 ( .A(MEM_stage_inst_dmem_n21636), .Z(MEM_stage_inst_dmem_n21619) );
BUF_X1 MEM_stage_inst_dmem_U228 ( .A(MEM_stage_inst_dmem_n21636), .Z(MEM_stage_inst_dmem_n21618) );
BUF_X1 MEM_stage_inst_dmem_U227 ( .A(MEM_stage_inst_dmem_n21637), .Z(MEM_stage_inst_dmem_n21617) );
BUF_X1 MEM_stage_inst_dmem_U226 ( .A(MEM_stage_inst_dmem_n21637), .Z(MEM_stage_inst_dmem_n21616) );
BUF_X1 MEM_stage_inst_dmem_U225 ( .A(MEM_stage_inst_dmem_n21637), .Z(MEM_stage_inst_dmem_n21615) );
BUF_X1 MEM_stage_inst_dmem_U224 ( .A(MEM_stage_inst_dmem_n21637), .Z(MEM_stage_inst_dmem_n21614) );
BUF_X1 MEM_stage_inst_dmem_U223 ( .A(MEM_stage_inst_dmem_n21637), .Z(MEM_stage_inst_dmem_n21613) );
BUF_X1 MEM_stage_inst_dmem_U222 ( .A(MEM_stage_inst_dmem_n21613), .Z(MEM_stage_inst_dmem_n21612) );
BUF_X1 MEM_stage_inst_dmem_U221 ( .A(MEM_stage_inst_dmem_n21613), .Z(MEM_stage_inst_dmem_n21611) );
BUF_X1 MEM_stage_inst_dmem_U220 ( .A(MEM_stage_inst_dmem_n21613), .Z(MEM_stage_inst_dmem_n21610) );
BUF_X1 MEM_stage_inst_dmem_U219 ( .A(MEM_stage_inst_dmem_n21613), .Z(MEM_stage_inst_dmem_n21609) );
BUF_X1 MEM_stage_inst_dmem_U218 ( .A(MEM_stage_inst_dmem_n21613), .Z(MEM_stage_inst_dmem_n21608) );
BUF_X1 MEM_stage_inst_dmem_U217 ( .A(MEM_stage_inst_dmem_n21614), .Z(MEM_stage_inst_dmem_n21607) );
BUF_X1 MEM_stage_inst_dmem_U216 ( .A(MEM_stage_inst_dmem_n21614), .Z(MEM_stage_inst_dmem_n21606) );
BUF_X1 MEM_stage_inst_dmem_U215 ( .A(MEM_stage_inst_dmem_n21614), .Z(MEM_stage_inst_dmem_n21605) );
BUF_X1 MEM_stage_inst_dmem_U214 ( .A(MEM_stage_inst_dmem_n21614), .Z(MEM_stage_inst_dmem_n21604) );
BUF_X1 MEM_stage_inst_dmem_U213 ( .A(MEM_stage_inst_dmem_n21614), .Z(MEM_stage_inst_dmem_n21603) );
BUF_X1 MEM_stage_inst_dmem_U212 ( .A(MEM_stage_inst_dmem_n21615), .Z(MEM_stage_inst_dmem_n21602) );
BUF_X1 MEM_stage_inst_dmem_U211 ( .A(MEM_stage_inst_dmem_n21615), .Z(MEM_stage_inst_dmem_n21601) );
BUF_X1 MEM_stage_inst_dmem_U210 ( .A(MEM_stage_inst_dmem_n21615), .Z(MEM_stage_inst_dmem_n21600) );
BUF_X1 MEM_stage_inst_dmem_U209 ( .A(MEM_stage_inst_dmem_n21615), .Z(MEM_stage_inst_dmem_n21599) );
BUF_X1 MEM_stage_inst_dmem_U208 ( .A(MEM_stage_inst_dmem_n21615), .Z(MEM_stage_inst_dmem_n21598) );
BUF_X1 MEM_stage_inst_dmem_U207 ( .A(MEM_stage_inst_dmem_n21616), .Z(MEM_stage_inst_dmem_n21597) );
BUF_X1 MEM_stage_inst_dmem_U206 ( .A(MEM_stage_inst_dmem_n21616), .Z(MEM_stage_inst_dmem_n21596) );
BUF_X1 MEM_stage_inst_dmem_U205 ( .A(MEM_stage_inst_dmem_n21616), .Z(MEM_stage_inst_dmem_n21595) );
BUF_X1 MEM_stage_inst_dmem_U204 ( .A(MEM_stage_inst_dmem_n21616), .Z(MEM_stage_inst_dmem_n21594) );
BUF_X1 MEM_stage_inst_dmem_U203 ( .A(MEM_stage_inst_dmem_n21616), .Z(MEM_stage_inst_dmem_n21593) );
BUF_X1 MEM_stage_inst_dmem_U202 ( .A(MEM_stage_inst_dmem_n21617), .Z(MEM_stage_inst_dmem_n21592) );
BUF_X1 MEM_stage_inst_dmem_U201 ( .A(MEM_stage_inst_dmem_n21617), .Z(MEM_stage_inst_dmem_n21591) );
BUF_X1 MEM_stage_inst_dmem_U200 ( .A(MEM_stage_inst_dmem_n21617), .Z(MEM_stage_inst_dmem_n21590) );
BUF_X1 MEM_stage_inst_dmem_U199 ( .A(MEM_stage_inst_dmem_n21617), .Z(MEM_stage_inst_dmem_n21589) );
BUF_X1 MEM_stage_inst_dmem_U198 ( .A(MEM_stage_inst_dmem_n21617), .Z(MEM_stage_inst_dmem_n21588) );
BUF_X1 MEM_stage_inst_dmem_U197 ( .A(MEM_stage_inst_dmem_n21618), .Z(MEM_stage_inst_dmem_n21587) );
BUF_X1 MEM_stage_inst_dmem_U196 ( .A(MEM_stage_inst_dmem_n21618), .Z(MEM_stage_inst_dmem_n21586) );
BUF_X1 MEM_stage_inst_dmem_U195 ( .A(MEM_stage_inst_dmem_n21618), .Z(MEM_stage_inst_dmem_n21585) );
BUF_X1 MEM_stage_inst_dmem_U194 ( .A(MEM_stage_inst_dmem_n21618), .Z(MEM_stage_inst_dmem_n21584) );
BUF_X1 MEM_stage_inst_dmem_U193 ( .A(MEM_stage_inst_dmem_n21618), .Z(MEM_stage_inst_dmem_n21583) );
BUF_X1 MEM_stage_inst_dmem_U192 ( .A(MEM_stage_inst_dmem_n21619), .Z(MEM_stage_inst_dmem_n21582) );
BUF_X1 MEM_stage_inst_dmem_U191 ( .A(MEM_stage_inst_dmem_n21619), .Z(MEM_stage_inst_dmem_n21581) );
BUF_X1 MEM_stage_inst_dmem_U190 ( .A(MEM_stage_inst_dmem_n21619), .Z(MEM_stage_inst_dmem_n21580) );
BUF_X1 MEM_stage_inst_dmem_U189 ( .A(MEM_stage_inst_dmem_n21619), .Z(MEM_stage_inst_dmem_n21579) );
BUF_X1 MEM_stage_inst_dmem_U188 ( .A(MEM_stage_inst_dmem_n21619), .Z(MEM_stage_inst_dmem_n21578) );
BUF_X1 MEM_stage_inst_dmem_U187 ( .A(MEM_stage_inst_dmem_n21620), .Z(MEM_stage_inst_dmem_n21577) );
BUF_X1 MEM_stage_inst_dmem_U186 ( .A(MEM_stage_inst_dmem_n21620), .Z(MEM_stage_inst_dmem_n21576) );
BUF_X1 MEM_stage_inst_dmem_U185 ( .A(MEM_stage_inst_dmem_n21620), .Z(MEM_stage_inst_dmem_n21575) );
BUF_X1 MEM_stage_inst_dmem_U184 ( .A(MEM_stage_inst_dmem_n21620), .Z(MEM_stage_inst_dmem_n21574) );
BUF_X1 MEM_stage_inst_dmem_U183 ( .A(MEM_stage_inst_dmem_n21620), .Z(MEM_stage_inst_dmem_n21573) );
BUF_X1 MEM_stage_inst_dmem_U182 ( .A(MEM_stage_inst_dmem_n21621), .Z(MEM_stage_inst_dmem_n21572) );
BUF_X1 MEM_stage_inst_dmem_U181 ( .A(MEM_stage_inst_dmem_n21621), .Z(MEM_stage_inst_dmem_n21571) );
BUF_X1 MEM_stage_inst_dmem_U180 ( .A(MEM_stage_inst_dmem_n21621), .Z(MEM_stage_inst_dmem_n21570) );
BUF_X1 MEM_stage_inst_dmem_U179 ( .A(MEM_stage_inst_dmem_n21621), .Z(MEM_stage_inst_dmem_n21569) );
BUF_X1 MEM_stage_inst_dmem_U178 ( .A(MEM_stage_inst_dmem_n21621), .Z(MEM_stage_inst_dmem_n21568) );
BUF_X1 MEM_stage_inst_dmem_U177 ( .A(MEM_stage_inst_dmem_n21622), .Z(MEM_stage_inst_dmem_n21567) );
BUF_X1 MEM_stage_inst_dmem_U176 ( .A(MEM_stage_inst_dmem_n21622), .Z(MEM_stage_inst_dmem_n21566) );
BUF_X1 MEM_stage_inst_dmem_U175 ( .A(MEM_stage_inst_dmem_n21622), .Z(MEM_stage_inst_dmem_n21565) );
BUF_X1 MEM_stage_inst_dmem_U174 ( .A(MEM_stage_inst_dmem_n21622), .Z(MEM_stage_inst_dmem_n21564) );
BUF_X1 MEM_stage_inst_dmem_U173 ( .A(MEM_stage_inst_dmem_n21622), .Z(MEM_stage_inst_dmem_n21563) );
BUF_X1 MEM_stage_inst_dmem_U172 ( .A(MEM_stage_inst_dmem_n21623), .Z(MEM_stage_inst_dmem_n21562) );
BUF_X1 MEM_stage_inst_dmem_U171 ( .A(MEM_stage_inst_dmem_n21623), .Z(MEM_stage_inst_dmem_n21561) );
BUF_X1 MEM_stage_inst_dmem_U170 ( .A(MEM_stage_inst_dmem_n21623), .Z(MEM_stage_inst_dmem_n21560) );
BUF_X1 MEM_stage_inst_dmem_U169 ( .A(MEM_stage_inst_dmem_n21623), .Z(MEM_stage_inst_dmem_n21559) );
BUF_X1 MEM_stage_inst_dmem_U168 ( .A(MEM_stage_inst_dmem_n21623), .Z(MEM_stage_inst_dmem_n21558) );
BUF_X1 MEM_stage_inst_dmem_U167 ( .A(MEM_stage_inst_dmem_n21624), .Z(MEM_stage_inst_dmem_n21557) );
BUF_X1 MEM_stage_inst_dmem_U166 ( .A(MEM_stage_inst_dmem_n21624), .Z(MEM_stage_inst_dmem_n21556) );
BUF_X1 MEM_stage_inst_dmem_U165 ( .A(MEM_stage_inst_dmem_n21624), .Z(MEM_stage_inst_dmem_n21555) );
BUF_X1 MEM_stage_inst_dmem_U164 ( .A(MEM_stage_inst_dmem_n21624), .Z(MEM_stage_inst_dmem_n21554) );
BUF_X1 MEM_stage_inst_dmem_U163 ( .A(MEM_stage_inst_dmem_n21624), .Z(MEM_stage_inst_dmem_n21553) );
BUF_X1 MEM_stage_inst_dmem_U162 ( .A(MEM_stage_inst_dmem_n21625), .Z(MEM_stage_inst_dmem_n21552) );
BUF_X1 MEM_stage_inst_dmem_U161 ( .A(MEM_stage_inst_dmem_n21625), .Z(MEM_stage_inst_dmem_n21551) );
BUF_X1 MEM_stage_inst_dmem_U160 ( .A(MEM_stage_inst_dmem_n21625), .Z(MEM_stage_inst_dmem_n21550) );
BUF_X1 MEM_stage_inst_dmem_U159 ( .A(MEM_stage_inst_dmem_n21625), .Z(MEM_stage_inst_dmem_n21549) );
BUF_X1 MEM_stage_inst_dmem_U158 ( .A(MEM_stage_inst_dmem_n21625), .Z(MEM_stage_inst_dmem_n21548) );
BUF_X1 MEM_stage_inst_dmem_U157 ( .A(MEM_stage_inst_dmem_n21626), .Z(MEM_stage_inst_dmem_n21547) );
BUF_X1 MEM_stage_inst_dmem_U156 ( .A(MEM_stage_inst_dmem_n21626), .Z(MEM_stage_inst_dmem_n21546) );
BUF_X1 MEM_stage_inst_dmem_U155 ( .A(MEM_stage_inst_dmem_n21626), .Z(MEM_stage_inst_dmem_n21545) );
BUF_X1 MEM_stage_inst_dmem_U154 ( .A(MEM_stage_inst_dmem_n21626), .Z(MEM_stage_inst_dmem_n21544) );
BUF_X1 MEM_stage_inst_dmem_U153 ( .A(MEM_stage_inst_dmem_n21626), .Z(MEM_stage_inst_dmem_n21543) );
BUF_X1 MEM_stage_inst_dmem_U152 ( .A(MEM_stage_inst_dmem_n21627), .Z(MEM_stage_inst_dmem_n21542) );
BUF_X1 MEM_stage_inst_dmem_U151 ( .A(MEM_stage_inst_dmem_n21627), .Z(MEM_stage_inst_dmem_n21541) );
BUF_X1 MEM_stage_inst_dmem_U150 ( .A(MEM_stage_inst_dmem_n21627), .Z(MEM_stage_inst_dmem_n21540) );
BUF_X1 MEM_stage_inst_dmem_U149 ( .A(MEM_stage_inst_dmem_n21627), .Z(MEM_stage_inst_dmem_n21539) );
BUF_X1 MEM_stage_inst_dmem_U148 ( .A(MEM_stage_inst_dmem_n21627), .Z(MEM_stage_inst_dmem_n21538) );
BUF_X1 MEM_stage_inst_dmem_U147 ( .A(MEM_stage_inst_dmem_n21628), .Z(MEM_stage_inst_dmem_n21537) );
BUF_X1 MEM_stage_inst_dmem_U146 ( .A(MEM_stage_inst_dmem_n21628), .Z(MEM_stage_inst_dmem_n21536) );
BUF_X1 MEM_stage_inst_dmem_U145 ( .A(MEM_stage_inst_dmem_n21628), .Z(MEM_stage_inst_dmem_n21535) );
BUF_X1 MEM_stage_inst_dmem_U144 ( .A(MEM_stage_inst_dmem_n21628), .Z(MEM_stage_inst_dmem_n21534) );
BUF_X1 MEM_stage_inst_dmem_U143 ( .A(MEM_stage_inst_dmem_n21628), .Z(MEM_stage_inst_dmem_n21533) );
BUF_X1 MEM_stage_inst_dmem_U142 ( .A(MEM_stage_inst_dmem_n21629), .Z(MEM_stage_inst_dmem_n21532) );
BUF_X1 MEM_stage_inst_dmem_U141 ( .A(MEM_stage_inst_dmem_n21629), .Z(MEM_stage_inst_dmem_n21531) );
BUF_X1 MEM_stage_inst_dmem_U140 ( .A(MEM_stage_inst_dmem_n21629), .Z(MEM_stage_inst_dmem_n21530) );
BUF_X1 MEM_stage_inst_dmem_U136 ( .A(MEM_stage_inst_dmem_n21629), .Z(MEM_stage_inst_dmem_n21529) );
BUF_X1 MEM_stage_inst_dmem_U121 ( .A(MEM_stage_inst_dmem_n21629), .Z(MEM_stage_inst_dmem_n21528) );
BUF_X1 MEM_stage_inst_dmem_U120 ( .A(MEM_stage_inst_dmem_n21630), .Z(MEM_stage_inst_dmem_n21527) );
BUF_X1 MEM_stage_inst_dmem_U119 ( .A(MEM_stage_inst_dmem_n21630), .Z(MEM_stage_inst_dmem_n21526) );
BUF_X1 MEM_stage_inst_dmem_U117 ( .A(MEM_stage_inst_dmem_n21630), .Z(MEM_stage_inst_dmem_n21525) );
BUF_X1 MEM_stage_inst_dmem_U115 ( .A(MEM_stage_inst_dmem_n21630), .Z(MEM_stage_inst_dmem_n21524) );
BUF_X1 MEM_stage_inst_dmem_U114 ( .A(MEM_stage_inst_dmem_n21630), .Z(MEM_stage_inst_dmem_n21523) );
BUF_X1 MEM_stage_inst_dmem_U113 ( .A(MEM_stage_inst_dmem_n21631), .Z(MEM_stage_inst_dmem_n21522) );
BUF_X1 MEM_stage_inst_dmem_U112 ( .A(MEM_stage_inst_dmem_n21631), .Z(MEM_stage_inst_dmem_n21521) );
BUF_X1 MEM_stage_inst_dmem_U111 ( .A(MEM_stage_inst_dmem_n21631), .Z(MEM_stage_inst_dmem_n21520) );
BUF_X1 MEM_stage_inst_dmem_U110 ( .A(MEM_stage_inst_dmem_n21631), .Z(MEM_stage_inst_dmem_n21519) );
BUF_X1 MEM_stage_inst_dmem_U109 ( .A(MEM_stage_inst_dmem_n21631), .Z(MEM_stage_inst_dmem_n21518) );
BUF_X1 MEM_stage_inst_dmem_U108 ( .A(MEM_stage_inst_dmem_n21632), .Z(MEM_stage_inst_dmem_n21517) );
BUF_X1 MEM_stage_inst_dmem_U107 ( .A(MEM_stage_inst_dmem_n21632), .Z(MEM_stage_inst_dmem_n21516) );
BUF_X1 MEM_stage_inst_dmem_U106 ( .A(MEM_stage_inst_dmem_n21632), .Z(MEM_stage_inst_dmem_n21515) );
BUF_X1 MEM_stage_inst_dmem_U105 ( .A(MEM_stage_inst_dmem_n21632), .Z(MEM_stage_inst_dmem_n21514) );
BUF_X1 MEM_stage_inst_dmem_U104 ( .A(MEM_stage_inst_dmem_n21632), .Z(MEM_stage_inst_dmem_n21513) );
BUF_X1 MEM_stage_inst_dmem_U103 ( .A(MEM_stage_inst_dmem_n21636), .Z(MEM_stage_inst_dmem_n21512) );
BUF_X1 MEM_stage_inst_dmem_U102 ( .A(MEM_stage_inst_dmem_n21633), .Z(MEM_stage_inst_dmem_n21511) );
BUF_X1 MEM_stage_inst_dmem_U101 ( .A(MEM_stage_inst_dmem_n21633), .Z(MEM_stage_inst_dmem_n21510) );
BUF_X1 MEM_stage_inst_dmem_U100 ( .A(MEM_stage_inst_dmem_n21633), .Z(MEM_stage_inst_dmem_n21509) );
BUF_X2 MEM_stage_inst_dmem_U99 ( .A(MEM_stage_inst_dmem_n20533), .Z(MEM_stage_inst_dmem_n21340) );
BUF_X1 MEM_stage_inst_dmem_U98 ( .A(MEM_stage_inst_dmem_n20536), .Z(MEM_stage_inst_dmem_n19260) );
INV_X8 MEM_stage_inst_dmem_U97 ( .A(MEM_stage_inst_dmem_n21507), .ZN(MEM_stage_inst_dmem_n21508) );
INV_X1 MEM_stage_inst_dmem_U27 ( .A(MEM_stage_inst_dmem_n19260), .ZN(MEM_stage_inst_dmem_n21507) );
BUF_X1 MEM_stage_inst_dmem_U19 ( .A(MEM_stage_inst_dmem_n20541), .Z(MEM_stage_inst_dmem_n19266) );
INV_X8 MEM_stage_inst_dmem_U15 ( .A(MEM_stage_inst_dmem_n21505), .ZN(MEM_stage_inst_dmem_n21506) );
INV_X1 MEM_stage_inst_dmem_U2 ( .A(MEM_stage_inst_dmem_n19266), .ZN(MEM_stage_inst_dmem_n21505) );
INV_X8 MEM_stage_inst_dmem_U11 ( .A(MEM_stage_inst_dmem_n5), .ZN(MEM_stage_inst_dmem_n6) );
NAND2_X1 MEM_stage_inst_dmem_U21512 ( .A1(MEM_stage_inst_dmem_n21503), .A2(MEM_stage_inst_dmem_n21502), .ZN(MEM_stage_inst_dmem_n8763) );
NAND2_X1 MEM_stage_inst_dmem_U21511 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n21500), .ZN(MEM_stage_inst_dmem_n21502) );
NAND2_X1 MEM_stage_inst_dmem_U21510 ( .A1(MEM_stage_inst_dmem_ram_3584), .A2(MEM_stage_inst_dmem_n21499), .ZN(MEM_stage_inst_dmem_n21503) );
NAND2_X1 MEM_stage_inst_dmem_U21509 ( .A1(MEM_stage_inst_dmem_n21498), .A2(MEM_stage_inst_dmem_n21497), .ZN(MEM_stage_inst_dmem_n8764) );
NAND2_X1 MEM_stage_inst_dmem_U21508 ( .A1(MEM_stage_inst_dmem_n109), .A2(MEM_stage_inst_dmem_n21500), .ZN(MEM_stage_inst_dmem_n21497) );
NAND2_X1 MEM_stage_inst_dmem_U21507 ( .A1(MEM_stage_inst_dmem_ram_3585), .A2(MEM_stage_inst_dmem_n21499), .ZN(MEM_stage_inst_dmem_n21498) );
NAND2_X1 MEM_stage_inst_dmem_U21506 ( .A1(MEM_stage_inst_dmem_n21496), .A2(MEM_stage_inst_dmem_n21495), .ZN(MEM_stage_inst_dmem_n8765) );
NAND2_X1 MEM_stage_inst_dmem_U21505 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n21500), .ZN(MEM_stage_inst_dmem_n21495) );
NAND2_X1 MEM_stage_inst_dmem_U21504 ( .A1(MEM_stage_inst_dmem_ram_3586), .A2(MEM_stage_inst_dmem_n21499), .ZN(MEM_stage_inst_dmem_n21496) );
NAND2_X1 MEM_stage_inst_dmem_U21503 ( .A1(MEM_stage_inst_dmem_n21494), .A2(MEM_stage_inst_dmem_n21493), .ZN(MEM_stage_inst_dmem_n8766) );
NAND2_X1 MEM_stage_inst_dmem_U21502 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n21500), .ZN(MEM_stage_inst_dmem_n21493) );
NAND2_X1 MEM_stage_inst_dmem_U21501 ( .A1(MEM_stage_inst_dmem_ram_3587), .A2(MEM_stage_inst_dmem_n21499), .ZN(MEM_stage_inst_dmem_n21494) );
NAND2_X1 MEM_stage_inst_dmem_U21500 ( .A1(MEM_stage_inst_dmem_n21492), .A2(MEM_stage_inst_dmem_n21491), .ZN(MEM_stage_inst_dmem_n8767) );
NAND2_X1 MEM_stage_inst_dmem_U21499 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n21500), .ZN(MEM_stage_inst_dmem_n21491) );
NAND2_X1 MEM_stage_inst_dmem_U21498 ( .A1(MEM_stage_inst_dmem_ram_3588), .A2(MEM_stage_inst_dmem_n21499), .ZN(MEM_stage_inst_dmem_n21492) );
NAND2_X1 MEM_stage_inst_dmem_U21497 ( .A1(MEM_stage_inst_dmem_n21490), .A2(MEM_stage_inst_dmem_n21489), .ZN(MEM_stage_inst_dmem_n8768) );
NAND2_X1 MEM_stage_inst_dmem_U21496 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n21500), .ZN(MEM_stage_inst_dmem_n21489) );
NAND2_X1 MEM_stage_inst_dmem_U21495 ( .A1(MEM_stage_inst_dmem_ram_3589), .A2(MEM_stage_inst_dmem_n21499), .ZN(MEM_stage_inst_dmem_n21490) );
NAND2_X1 MEM_stage_inst_dmem_U21494 ( .A1(MEM_stage_inst_dmem_n21488), .A2(MEM_stage_inst_dmem_n21487), .ZN(MEM_stage_inst_dmem_n8769) );
NAND2_X1 MEM_stage_inst_dmem_U21493 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n21500), .ZN(MEM_stage_inst_dmem_n21487) );
NAND2_X1 MEM_stage_inst_dmem_U21492 ( .A1(MEM_stage_inst_dmem_ram_3590), .A2(MEM_stage_inst_dmem_n21499), .ZN(MEM_stage_inst_dmem_n21488) );
NAND2_X1 MEM_stage_inst_dmem_U21491 ( .A1(MEM_stage_inst_dmem_n21486), .A2(MEM_stage_inst_dmem_n21485), .ZN(MEM_stage_inst_dmem_n8770) );
NAND2_X1 MEM_stage_inst_dmem_U21490 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n21500), .ZN(MEM_stage_inst_dmem_n21485) );
NAND2_X1 MEM_stage_inst_dmem_U21489 ( .A1(MEM_stage_inst_dmem_ram_3591), .A2(MEM_stage_inst_dmem_n21499), .ZN(MEM_stage_inst_dmem_n21486) );
NAND2_X1 MEM_stage_inst_dmem_U21488 ( .A1(MEM_stage_inst_dmem_n21484), .A2(MEM_stage_inst_dmem_n21483), .ZN(MEM_stage_inst_dmem_n8771) );
NAND2_X1 MEM_stage_inst_dmem_U21487 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n21500), .ZN(MEM_stage_inst_dmem_n21483) );
NAND2_X1 MEM_stage_inst_dmem_U21486 ( .A1(MEM_stage_inst_dmem_ram_3592), .A2(MEM_stage_inst_dmem_n21499), .ZN(MEM_stage_inst_dmem_n21484) );
NAND2_X1 MEM_stage_inst_dmem_U21485 ( .A1(MEM_stage_inst_dmem_n21482), .A2(MEM_stage_inst_dmem_n21481), .ZN(MEM_stage_inst_dmem_n8772) );
NAND2_X1 MEM_stage_inst_dmem_U21484 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n21500), .ZN(MEM_stage_inst_dmem_n21481) );
NAND2_X1 MEM_stage_inst_dmem_U21483 ( .A1(MEM_stage_inst_dmem_ram_3593), .A2(MEM_stage_inst_dmem_n21499), .ZN(MEM_stage_inst_dmem_n21482) );
NAND2_X1 MEM_stage_inst_dmem_U21482 ( .A1(MEM_stage_inst_dmem_n21480), .A2(MEM_stage_inst_dmem_n21479), .ZN(MEM_stage_inst_dmem_n8773) );
NAND2_X1 MEM_stage_inst_dmem_U21481 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n21500), .ZN(MEM_stage_inst_dmem_n21479) );
NAND2_X1 MEM_stage_inst_dmem_U21480 ( .A1(MEM_stage_inst_dmem_ram_3594), .A2(MEM_stage_inst_dmem_n21499), .ZN(MEM_stage_inst_dmem_n21480) );
NAND2_X1 MEM_stage_inst_dmem_U21479 ( .A1(MEM_stage_inst_dmem_n21478), .A2(MEM_stage_inst_dmem_n21477), .ZN(MEM_stage_inst_dmem_n8774) );
NAND2_X1 MEM_stage_inst_dmem_U21478 ( .A1(MEM_stage_inst_dmem_n14705), .A2(MEM_stage_inst_dmem_n21500), .ZN(MEM_stage_inst_dmem_n21477) );
NAND2_X1 MEM_stage_inst_dmem_U21477 ( .A1(MEM_stage_inst_dmem_ram_3595), .A2(MEM_stage_inst_dmem_n21499), .ZN(MEM_stage_inst_dmem_n21478) );
NAND2_X1 MEM_stage_inst_dmem_U21476 ( .A1(MEM_stage_inst_dmem_n21476), .A2(MEM_stage_inst_dmem_n21475), .ZN(MEM_stage_inst_dmem_n8775) );
NAND2_X1 MEM_stage_inst_dmem_U21475 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n21500), .ZN(MEM_stage_inst_dmem_n21475) );
NAND2_X1 MEM_stage_inst_dmem_U21474 ( .A1(MEM_stage_inst_dmem_ram_3596), .A2(MEM_stage_inst_dmem_n21499), .ZN(MEM_stage_inst_dmem_n21476) );
NAND2_X1 MEM_stage_inst_dmem_U21473 ( .A1(MEM_stage_inst_dmem_n21473), .A2(MEM_stage_inst_dmem_n21472), .ZN(MEM_stage_inst_dmem_n8776) );
NAND2_X1 MEM_stage_inst_dmem_U21472 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n21500), .ZN(MEM_stage_inst_dmem_n21472) );
NAND2_X1 MEM_stage_inst_dmem_U21471 ( .A1(MEM_stage_inst_dmem_ram_3597), .A2(MEM_stage_inst_dmem_n21499), .ZN(MEM_stage_inst_dmem_n21473) );
NAND2_X1 MEM_stage_inst_dmem_U21470 ( .A1(MEM_stage_inst_dmem_n21470), .A2(MEM_stage_inst_dmem_n21469), .ZN(MEM_stage_inst_dmem_n8777) );
NAND2_X1 MEM_stage_inst_dmem_U21469 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n21500), .ZN(MEM_stage_inst_dmem_n21469) );
NAND2_X1 MEM_stage_inst_dmem_U21468 ( .A1(MEM_stage_inst_dmem_ram_3598), .A2(MEM_stage_inst_dmem_n21499), .ZN(MEM_stage_inst_dmem_n21470) );
NAND2_X1 MEM_stage_inst_dmem_U21467 ( .A1(MEM_stage_inst_dmem_n21467), .A2(MEM_stage_inst_dmem_n21466), .ZN(MEM_stage_inst_dmem_n8778) );
NAND2_X1 MEM_stage_inst_dmem_U21466 ( .A1(MEM_stage_inst_dmem_n20506), .A2(MEM_stage_inst_dmem_n21500), .ZN(MEM_stage_inst_dmem_n21466) );
NAND2_X1 MEM_stage_inst_dmem_U21465 ( .A1(MEM_stage_inst_dmem_ram_3599), .A2(MEM_stage_inst_dmem_n21499), .ZN(MEM_stage_inst_dmem_n21467) );
NAND2_X1 MEM_stage_inst_dmem_U21464 ( .A1(MEM_stage_inst_dmem_n21465), .A2(MEM_stage_inst_dmem_n21464), .ZN(MEM_stage_inst_dmem_n21499) );
NAND2_X1 MEM_stage_inst_dmem_U21463 ( .A1(MEM_stage_inst_dmem_n21463), .A2(MEM_stage_inst_dmem_n21462), .ZN(MEM_stage_inst_dmem_n8779) );
NAND2_X1 MEM_stage_inst_dmem_U21462 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n21461), .ZN(MEM_stage_inst_dmem_n21462) );
NAND2_X1 MEM_stage_inst_dmem_U21461 ( .A1(MEM_stage_inst_dmem_ram_3600), .A2(MEM_stage_inst_dmem_n21460), .ZN(MEM_stage_inst_dmem_n21463) );
NAND2_X1 MEM_stage_inst_dmem_U21460 ( .A1(MEM_stage_inst_dmem_n21459), .A2(MEM_stage_inst_dmem_n21458), .ZN(MEM_stage_inst_dmem_n8780) );
NAND2_X1 MEM_stage_inst_dmem_U21459 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n21461), .ZN(MEM_stage_inst_dmem_n21458) );
NAND2_X1 MEM_stage_inst_dmem_U21458 ( .A1(MEM_stage_inst_dmem_ram_3601), .A2(MEM_stage_inst_dmem_n21460), .ZN(MEM_stage_inst_dmem_n21459) );
NAND2_X1 MEM_stage_inst_dmem_U21457 ( .A1(MEM_stage_inst_dmem_n21457), .A2(MEM_stage_inst_dmem_n21456), .ZN(MEM_stage_inst_dmem_n8781) );
NAND2_X1 MEM_stage_inst_dmem_U21456 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n21461), .ZN(MEM_stage_inst_dmem_n21456) );
NAND2_X1 MEM_stage_inst_dmem_U21455 ( .A1(MEM_stage_inst_dmem_ram_3602), .A2(MEM_stage_inst_dmem_n21460), .ZN(MEM_stage_inst_dmem_n21457) );
NAND2_X1 MEM_stage_inst_dmem_U21454 ( .A1(MEM_stage_inst_dmem_n21455), .A2(MEM_stage_inst_dmem_n21454), .ZN(MEM_stage_inst_dmem_n8782) );
NAND2_X1 MEM_stage_inst_dmem_U21453 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n21461), .ZN(MEM_stage_inst_dmem_n21454) );
NAND2_X1 MEM_stage_inst_dmem_U21452 ( .A1(MEM_stage_inst_dmem_ram_3603), .A2(MEM_stage_inst_dmem_n21460), .ZN(MEM_stage_inst_dmem_n21455) );
NAND2_X1 MEM_stage_inst_dmem_U21451 ( .A1(MEM_stage_inst_dmem_n21453), .A2(MEM_stage_inst_dmem_n21452), .ZN(MEM_stage_inst_dmem_n8783) );
NAND2_X1 MEM_stage_inst_dmem_U21450 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n21461), .ZN(MEM_stage_inst_dmem_n21452) );
NAND2_X1 MEM_stage_inst_dmem_U21449 ( .A1(MEM_stage_inst_dmem_ram_3604), .A2(MEM_stage_inst_dmem_n21460), .ZN(MEM_stage_inst_dmem_n21453) );
NAND2_X1 MEM_stage_inst_dmem_U21448 ( .A1(MEM_stage_inst_dmem_n21451), .A2(MEM_stage_inst_dmem_n21450), .ZN(MEM_stage_inst_dmem_n8784) );
NAND2_X1 MEM_stage_inst_dmem_U21447 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n21461), .ZN(MEM_stage_inst_dmem_n21450) );
NAND2_X1 MEM_stage_inst_dmem_U21446 ( .A1(MEM_stage_inst_dmem_ram_3605), .A2(MEM_stage_inst_dmem_n21460), .ZN(MEM_stage_inst_dmem_n21451) );
NAND2_X1 MEM_stage_inst_dmem_U21445 ( .A1(MEM_stage_inst_dmem_n21449), .A2(MEM_stage_inst_dmem_n21448), .ZN(MEM_stage_inst_dmem_n8785) );
NAND2_X1 MEM_stage_inst_dmem_U21444 ( .A1(MEM_stage_inst_dmem_n14717), .A2(MEM_stage_inst_dmem_n21461), .ZN(MEM_stage_inst_dmem_n21448) );
NAND2_X1 MEM_stage_inst_dmem_U21443 ( .A1(MEM_stage_inst_dmem_ram_3606), .A2(MEM_stage_inst_dmem_n21460), .ZN(MEM_stage_inst_dmem_n21449) );
NAND2_X1 MEM_stage_inst_dmem_U21442 ( .A1(MEM_stage_inst_dmem_n21447), .A2(MEM_stage_inst_dmem_n21446), .ZN(MEM_stage_inst_dmem_n8786) );
NAND2_X1 MEM_stage_inst_dmem_U21441 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n21461), .ZN(MEM_stage_inst_dmem_n21446) );
NAND2_X1 MEM_stage_inst_dmem_U21440 ( .A1(MEM_stage_inst_dmem_ram_3607), .A2(MEM_stage_inst_dmem_n21460), .ZN(MEM_stage_inst_dmem_n21447) );
NAND2_X1 MEM_stage_inst_dmem_U21439 ( .A1(MEM_stage_inst_dmem_n21445), .A2(MEM_stage_inst_dmem_n21444), .ZN(MEM_stage_inst_dmem_n8787) );
NAND2_X1 MEM_stage_inst_dmem_U21438 ( .A1(MEM_stage_inst_dmem_n18013), .A2(MEM_stage_inst_dmem_n21461), .ZN(MEM_stage_inst_dmem_n21444) );
NAND2_X1 MEM_stage_inst_dmem_U21437 ( .A1(MEM_stage_inst_dmem_ram_3608), .A2(MEM_stage_inst_dmem_n21460), .ZN(MEM_stage_inst_dmem_n21445) );
NAND2_X1 MEM_stage_inst_dmem_U21436 ( .A1(MEM_stage_inst_dmem_n21443), .A2(MEM_stage_inst_dmem_n21442), .ZN(MEM_stage_inst_dmem_n8788) );
NAND2_X1 MEM_stage_inst_dmem_U21435 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n21461), .ZN(MEM_stage_inst_dmem_n21442) );
NAND2_X1 MEM_stage_inst_dmem_U21434 ( .A1(MEM_stage_inst_dmem_ram_3609), .A2(MEM_stage_inst_dmem_n21460), .ZN(MEM_stage_inst_dmem_n21443) );
NAND2_X1 MEM_stage_inst_dmem_U21433 ( .A1(MEM_stage_inst_dmem_n21441), .A2(MEM_stage_inst_dmem_n21440), .ZN(MEM_stage_inst_dmem_n8789) );
NAND2_X1 MEM_stage_inst_dmem_U21432 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n21461), .ZN(MEM_stage_inst_dmem_n21440) );
NAND2_X1 MEM_stage_inst_dmem_U21431 ( .A1(MEM_stage_inst_dmem_ram_3610), .A2(MEM_stage_inst_dmem_n21460), .ZN(MEM_stage_inst_dmem_n21441) );
NAND2_X1 MEM_stage_inst_dmem_U21430 ( .A1(MEM_stage_inst_dmem_n21439), .A2(MEM_stage_inst_dmem_n21438), .ZN(MEM_stage_inst_dmem_n8790) );
NAND2_X1 MEM_stage_inst_dmem_U21429 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n21461), .ZN(MEM_stage_inst_dmem_n21438) );
NAND2_X1 MEM_stage_inst_dmem_U21428 ( .A1(MEM_stage_inst_dmem_ram_3611), .A2(MEM_stage_inst_dmem_n21460), .ZN(MEM_stage_inst_dmem_n21439) );
NAND2_X1 MEM_stage_inst_dmem_U21427 ( .A1(MEM_stage_inst_dmem_n21437), .A2(MEM_stage_inst_dmem_n21436), .ZN(MEM_stage_inst_dmem_n8791) );
NAND2_X1 MEM_stage_inst_dmem_U21426 ( .A1(MEM_stage_inst_dmem_n14702), .A2(MEM_stage_inst_dmem_n21461), .ZN(MEM_stage_inst_dmem_n21436) );
NAND2_X1 MEM_stage_inst_dmem_U21425 ( .A1(MEM_stage_inst_dmem_ram_3612), .A2(MEM_stage_inst_dmem_n21460), .ZN(MEM_stage_inst_dmem_n21437) );
NAND2_X1 MEM_stage_inst_dmem_U21424 ( .A1(MEM_stage_inst_dmem_n21435), .A2(MEM_stage_inst_dmem_n21434), .ZN(MEM_stage_inst_dmem_n8792) );
NAND2_X1 MEM_stage_inst_dmem_U21423 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n21461), .ZN(MEM_stage_inst_dmem_n21434) );
NAND2_X1 MEM_stage_inst_dmem_U21422 ( .A1(MEM_stage_inst_dmem_ram_3613), .A2(MEM_stage_inst_dmem_n21460), .ZN(MEM_stage_inst_dmem_n21435) );
NAND2_X1 MEM_stage_inst_dmem_U21421 ( .A1(MEM_stage_inst_dmem_n21433), .A2(MEM_stage_inst_dmem_n21432), .ZN(MEM_stage_inst_dmem_n8793) );
NAND2_X1 MEM_stage_inst_dmem_U21420 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n21461), .ZN(MEM_stage_inst_dmem_n21432) );
NAND2_X1 MEM_stage_inst_dmem_U21419 ( .A1(MEM_stage_inst_dmem_ram_3614), .A2(MEM_stage_inst_dmem_n21460), .ZN(MEM_stage_inst_dmem_n21433) );
NAND2_X1 MEM_stage_inst_dmem_U21418 ( .A1(MEM_stage_inst_dmem_n21431), .A2(MEM_stage_inst_dmem_n21430), .ZN(MEM_stage_inst_dmem_n8794) );
NAND2_X1 MEM_stage_inst_dmem_U21417 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n21461), .ZN(MEM_stage_inst_dmem_n21430) );
INV_X1 MEM_stage_inst_dmem_U21416 ( .A(MEM_stage_inst_dmem_n21460), .ZN(MEM_stage_inst_dmem_n21461) );
NAND2_X1 MEM_stage_inst_dmem_U21415 ( .A1(MEM_stage_inst_dmem_ram_3615), .A2(MEM_stage_inst_dmem_n21460), .ZN(MEM_stage_inst_dmem_n21431) );
NAND2_X1 MEM_stage_inst_dmem_U21414 ( .A1(MEM_stage_inst_dmem_n21429), .A2(MEM_stage_inst_dmem_n21464), .ZN(MEM_stage_inst_dmem_n21460) );
NAND2_X1 MEM_stage_inst_dmem_U21413 ( .A1(MEM_stage_inst_dmem_n21428), .A2(MEM_stage_inst_dmem_n21427), .ZN(MEM_stage_inst_dmem_n8795) );
NAND2_X1 MEM_stage_inst_dmem_U21412 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n21426), .ZN(MEM_stage_inst_dmem_n21427) );
NAND2_X1 MEM_stage_inst_dmem_U21411 ( .A1(MEM_stage_inst_dmem_ram_3616), .A2(MEM_stage_inst_dmem_n21425), .ZN(MEM_stage_inst_dmem_n21428) );
NAND2_X1 MEM_stage_inst_dmem_U21410 ( .A1(MEM_stage_inst_dmem_n21424), .A2(MEM_stage_inst_dmem_n21423), .ZN(MEM_stage_inst_dmem_n8796) );
NAND2_X1 MEM_stage_inst_dmem_U21409 ( .A1(MEM_stage_inst_dmem_n109), .A2(MEM_stage_inst_dmem_n21426), .ZN(MEM_stage_inst_dmem_n21423) );
NAND2_X1 MEM_stage_inst_dmem_U21408 ( .A1(MEM_stage_inst_dmem_ram_3617), .A2(MEM_stage_inst_dmem_n21425), .ZN(MEM_stage_inst_dmem_n21424) );
NAND2_X1 MEM_stage_inst_dmem_U21407 ( .A1(MEM_stage_inst_dmem_n21422), .A2(MEM_stage_inst_dmem_n21421), .ZN(MEM_stage_inst_dmem_n8797) );
NAND2_X1 MEM_stage_inst_dmem_U21406 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n21426), .ZN(MEM_stage_inst_dmem_n21421) );
NAND2_X1 MEM_stage_inst_dmem_U21405 ( .A1(MEM_stage_inst_dmem_ram_3618), .A2(MEM_stage_inst_dmem_n21425), .ZN(MEM_stage_inst_dmem_n21422) );
NAND2_X1 MEM_stage_inst_dmem_U21404 ( .A1(MEM_stage_inst_dmem_n21420), .A2(MEM_stage_inst_dmem_n21419), .ZN(MEM_stage_inst_dmem_n8798) );
NAND2_X1 MEM_stage_inst_dmem_U21403 ( .A1(MEM_stage_inst_dmem_n13064), .A2(MEM_stage_inst_dmem_n21426), .ZN(MEM_stage_inst_dmem_n21419) );
NAND2_X1 MEM_stage_inst_dmem_U21402 ( .A1(MEM_stage_inst_dmem_ram_3619), .A2(MEM_stage_inst_dmem_n21425), .ZN(MEM_stage_inst_dmem_n21420) );
NAND2_X1 MEM_stage_inst_dmem_U21401 ( .A1(MEM_stage_inst_dmem_n21418), .A2(MEM_stage_inst_dmem_n21417), .ZN(MEM_stage_inst_dmem_n8799) );
NAND2_X1 MEM_stage_inst_dmem_U21400 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n21426), .ZN(MEM_stage_inst_dmem_n21417) );
NAND2_X1 MEM_stage_inst_dmem_U21399 ( .A1(MEM_stage_inst_dmem_ram_3620), .A2(MEM_stage_inst_dmem_n21425), .ZN(MEM_stage_inst_dmem_n21418) );
NAND2_X1 MEM_stage_inst_dmem_U21398 ( .A1(MEM_stage_inst_dmem_n21416), .A2(MEM_stage_inst_dmem_n21415), .ZN(MEM_stage_inst_dmem_n8800) );
NAND2_X1 MEM_stage_inst_dmem_U21397 ( .A1(MEM_stage_inst_dmem_n13059), .A2(MEM_stage_inst_dmem_n21426), .ZN(MEM_stage_inst_dmem_n21415) );
NAND2_X1 MEM_stage_inst_dmem_U21396 ( .A1(MEM_stage_inst_dmem_ram_3621), .A2(MEM_stage_inst_dmem_n21425), .ZN(MEM_stage_inst_dmem_n21416) );
NAND2_X1 MEM_stage_inst_dmem_U21395 ( .A1(MEM_stage_inst_dmem_n21414), .A2(MEM_stage_inst_dmem_n21413), .ZN(MEM_stage_inst_dmem_n8801) );
NAND2_X1 MEM_stage_inst_dmem_U21394 ( .A1(MEM_stage_inst_dmem_n13056), .A2(MEM_stage_inst_dmem_n21426), .ZN(MEM_stage_inst_dmem_n21413) );
NAND2_X1 MEM_stage_inst_dmem_U21393 ( .A1(MEM_stage_inst_dmem_ram_3622), .A2(MEM_stage_inst_dmem_n21425), .ZN(MEM_stage_inst_dmem_n21414) );
NAND2_X1 MEM_stage_inst_dmem_U21392 ( .A1(MEM_stage_inst_dmem_n21412), .A2(MEM_stage_inst_dmem_n21411), .ZN(MEM_stage_inst_dmem_n8802) );
NAND2_X1 MEM_stage_inst_dmem_U21391 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n21426), .ZN(MEM_stage_inst_dmem_n21411) );
NAND2_X1 MEM_stage_inst_dmem_U21390 ( .A1(MEM_stage_inst_dmem_ram_3623), .A2(MEM_stage_inst_dmem_n21425), .ZN(MEM_stage_inst_dmem_n21412) );
NAND2_X1 MEM_stage_inst_dmem_U21389 ( .A1(MEM_stage_inst_dmem_n21410), .A2(MEM_stage_inst_dmem_n21409), .ZN(MEM_stage_inst_dmem_n8803) );
NAND2_X1 MEM_stage_inst_dmem_U21388 ( .A1(MEM_stage_inst_dmem_n111), .A2(MEM_stage_inst_dmem_n21426), .ZN(MEM_stage_inst_dmem_n21409) );
NAND2_X1 MEM_stage_inst_dmem_U21387 ( .A1(MEM_stage_inst_dmem_ram_3624), .A2(MEM_stage_inst_dmem_n21425), .ZN(MEM_stage_inst_dmem_n21410) );
NAND2_X1 MEM_stage_inst_dmem_U21386 ( .A1(MEM_stage_inst_dmem_n21408), .A2(MEM_stage_inst_dmem_n21407), .ZN(MEM_stage_inst_dmem_n8804) );
NAND2_X1 MEM_stage_inst_dmem_U21385 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n21426), .ZN(MEM_stage_inst_dmem_n21407) );
NAND2_X1 MEM_stage_inst_dmem_U21384 ( .A1(MEM_stage_inst_dmem_ram_3625), .A2(MEM_stage_inst_dmem_n21425), .ZN(MEM_stage_inst_dmem_n21408) );
NAND2_X1 MEM_stage_inst_dmem_U21383 ( .A1(MEM_stage_inst_dmem_n21406), .A2(MEM_stage_inst_dmem_n21405), .ZN(MEM_stage_inst_dmem_n8805) );
NAND2_X1 MEM_stage_inst_dmem_U21382 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n21426), .ZN(MEM_stage_inst_dmem_n21405) );
NAND2_X1 MEM_stage_inst_dmem_U21381 ( .A1(MEM_stage_inst_dmem_ram_3626), .A2(MEM_stage_inst_dmem_n21425), .ZN(MEM_stage_inst_dmem_n21406) );
NAND2_X1 MEM_stage_inst_dmem_U21380 ( .A1(MEM_stage_inst_dmem_n21404), .A2(MEM_stage_inst_dmem_n21403), .ZN(MEM_stage_inst_dmem_n8806) );
NAND2_X1 MEM_stage_inst_dmem_U21379 ( .A1(MEM_stage_inst_dmem_n13044), .A2(MEM_stage_inst_dmem_n21426), .ZN(MEM_stage_inst_dmem_n21403) );
NAND2_X1 MEM_stage_inst_dmem_U21378 ( .A1(MEM_stage_inst_dmem_ram_3627), .A2(MEM_stage_inst_dmem_n21425), .ZN(MEM_stage_inst_dmem_n21404) );
NAND2_X1 MEM_stage_inst_dmem_U21377 ( .A1(MEM_stage_inst_dmem_n21402), .A2(MEM_stage_inst_dmem_n21401), .ZN(MEM_stage_inst_dmem_n8807) );
NAND2_X1 MEM_stage_inst_dmem_U21376 ( .A1(MEM_stage_inst_dmem_n21474), .A2(MEM_stage_inst_dmem_n21426), .ZN(MEM_stage_inst_dmem_n21401) );
NAND2_X1 MEM_stage_inst_dmem_U21375 ( .A1(MEM_stage_inst_dmem_ram_3628), .A2(MEM_stage_inst_dmem_n21425), .ZN(MEM_stage_inst_dmem_n21402) );
NAND2_X1 MEM_stage_inst_dmem_U21374 ( .A1(MEM_stage_inst_dmem_n21400), .A2(MEM_stage_inst_dmem_n21399), .ZN(MEM_stage_inst_dmem_n8808) );
NAND2_X1 MEM_stage_inst_dmem_U21373 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n21426), .ZN(MEM_stage_inst_dmem_n21399) );
NAND2_X1 MEM_stage_inst_dmem_U21372 ( .A1(MEM_stage_inst_dmem_ram_3629), .A2(MEM_stage_inst_dmem_n21425), .ZN(MEM_stage_inst_dmem_n21400) );
NAND2_X1 MEM_stage_inst_dmem_U21371 ( .A1(MEM_stage_inst_dmem_n21398), .A2(MEM_stage_inst_dmem_n21397), .ZN(MEM_stage_inst_dmem_n8809) );
NAND2_X1 MEM_stage_inst_dmem_U21370 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n21426), .ZN(MEM_stage_inst_dmem_n21397) );
NAND2_X1 MEM_stage_inst_dmem_U21369 ( .A1(MEM_stage_inst_dmem_ram_3630), .A2(MEM_stage_inst_dmem_n21425), .ZN(MEM_stage_inst_dmem_n21398) );
NAND2_X1 MEM_stage_inst_dmem_U21368 ( .A1(MEM_stage_inst_dmem_n21396), .A2(MEM_stage_inst_dmem_n21395), .ZN(MEM_stage_inst_dmem_n8810) );
NAND2_X1 MEM_stage_inst_dmem_U21367 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n21426), .ZN(MEM_stage_inst_dmem_n21395) );
INV_X1 MEM_stage_inst_dmem_U21366 ( .A(MEM_stage_inst_dmem_n21425), .ZN(MEM_stage_inst_dmem_n21426) );
NAND2_X1 MEM_stage_inst_dmem_U21365 ( .A1(MEM_stage_inst_dmem_ram_3631), .A2(MEM_stage_inst_dmem_n21425), .ZN(MEM_stage_inst_dmem_n21396) );
NAND2_X1 MEM_stage_inst_dmem_U21364 ( .A1(MEM_stage_inst_dmem_n21394), .A2(MEM_stage_inst_dmem_n21464), .ZN(MEM_stage_inst_dmem_n21425) );
NAND2_X1 MEM_stage_inst_dmem_U21363 ( .A1(MEM_stage_inst_dmem_n21393), .A2(MEM_stage_inst_dmem_n21392), .ZN(MEM_stage_inst_dmem_n8811) );
NAND2_X1 MEM_stage_inst_dmem_U21362 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n21391), .ZN(MEM_stage_inst_dmem_n21392) );
NAND2_X1 MEM_stage_inst_dmem_U21361 ( .A1(MEM_stage_inst_dmem_ram_3632), .A2(MEM_stage_inst_dmem_n21390), .ZN(MEM_stage_inst_dmem_n21393) );
NAND2_X1 MEM_stage_inst_dmem_U21360 ( .A1(MEM_stage_inst_dmem_n21389), .A2(MEM_stage_inst_dmem_n21388), .ZN(MEM_stage_inst_dmem_n8812) );
NAND2_X1 MEM_stage_inst_dmem_U21359 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n21391), .ZN(MEM_stage_inst_dmem_n21388) );
NAND2_X1 MEM_stage_inst_dmem_U21358 ( .A1(MEM_stage_inst_dmem_ram_3633), .A2(MEM_stage_inst_dmem_n21390), .ZN(MEM_stage_inst_dmem_n21389) );
NAND2_X1 MEM_stage_inst_dmem_U21357 ( .A1(MEM_stage_inst_dmem_n21387), .A2(MEM_stage_inst_dmem_n21386), .ZN(MEM_stage_inst_dmem_n8813) );
NAND2_X1 MEM_stage_inst_dmem_U21356 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n21391), .ZN(MEM_stage_inst_dmem_n21386) );
NAND2_X1 MEM_stage_inst_dmem_U21355 ( .A1(MEM_stage_inst_dmem_ram_3634), .A2(MEM_stage_inst_dmem_n21390), .ZN(MEM_stage_inst_dmem_n21387) );
NAND2_X1 MEM_stage_inst_dmem_U21354 ( .A1(MEM_stage_inst_dmem_n21385), .A2(MEM_stage_inst_dmem_n21384), .ZN(MEM_stage_inst_dmem_n8814) );
NAND2_X1 MEM_stage_inst_dmem_U21353 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n21391), .ZN(MEM_stage_inst_dmem_n21384) );
NAND2_X1 MEM_stage_inst_dmem_U21352 ( .A1(MEM_stage_inst_dmem_ram_3635), .A2(MEM_stage_inst_dmem_n21390), .ZN(MEM_stage_inst_dmem_n21385) );
NAND2_X1 MEM_stage_inst_dmem_U21351 ( .A1(MEM_stage_inst_dmem_n21383), .A2(MEM_stage_inst_dmem_n21382), .ZN(MEM_stage_inst_dmem_n8815) );
NAND2_X1 MEM_stage_inst_dmem_U21350 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n21391), .ZN(MEM_stage_inst_dmem_n21382) );
NAND2_X1 MEM_stage_inst_dmem_U21349 ( .A1(MEM_stage_inst_dmem_ram_3636), .A2(MEM_stage_inst_dmem_n21390), .ZN(MEM_stage_inst_dmem_n21383) );
NAND2_X1 MEM_stage_inst_dmem_U21348 ( .A1(MEM_stage_inst_dmem_n21381), .A2(MEM_stage_inst_dmem_n21380), .ZN(MEM_stage_inst_dmem_n8816) );
NAND2_X1 MEM_stage_inst_dmem_U21347 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n21391), .ZN(MEM_stage_inst_dmem_n21380) );
NAND2_X1 MEM_stage_inst_dmem_U21346 ( .A1(MEM_stage_inst_dmem_ram_3637), .A2(MEM_stage_inst_dmem_n21390), .ZN(MEM_stage_inst_dmem_n21381) );
NAND2_X1 MEM_stage_inst_dmem_U21345 ( .A1(MEM_stage_inst_dmem_n21379), .A2(MEM_stage_inst_dmem_n21378), .ZN(MEM_stage_inst_dmem_n8817) );
NAND2_X1 MEM_stage_inst_dmem_U21344 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n21391), .ZN(MEM_stage_inst_dmem_n21378) );
NAND2_X1 MEM_stage_inst_dmem_U21343 ( .A1(MEM_stage_inst_dmem_ram_3638), .A2(MEM_stage_inst_dmem_n21390), .ZN(MEM_stage_inst_dmem_n21379) );
NAND2_X1 MEM_stage_inst_dmem_U21342 ( .A1(MEM_stage_inst_dmem_n21377), .A2(MEM_stage_inst_dmem_n21376), .ZN(MEM_stage_inst_dmem_n8818) );
NAND2_X1 MEM_stage_inst_dmem_U21341 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n21391), .ZN(MEM_stage_inst_dmem_n21376) );
NAND2_X1 MEM_stage_inst_dmem_U21340 ( .A1(MEM_stage_inst_dmem_ram_3639), .A2(MEM_stage_inst_dmem_n21390), .ZN(MEM_stage_inst_dmem_n21377) );
NAND2_X1 MEM_stage_inst_dmem_U21339 ( .A1(MEM_stage_inst_dmem_n21375), .A2(MEM_stage_inst_dmem_n21374), .ZN(MEM_stage_inst_dmem_n8819) );
NAND2_X1 MEM_stage_inst_dmem_U21338 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n21391), .ZN(MEM_stage_inst_dmem_n21374) );
NAND2_X1 MEM_stage_inst_dmem_U21337 ( .A1(MEM_stage_inst_dmem_ram_3640), .A2(MEM_stage_inst_dmem_n21390), .ZN(MEM_stage_inst_dmem_n21375) );
NAND2_X1 MEM_stage_inst_dmem_U21336 ( .A1(MEM_stage_inst_dmem_n21373), .A2(MEM_stage_inst_dmem_n21372), .ZN(MEM_stage_inst_dmem_n8820) );
NAND2_X1 MEM_stage_inst_dmem_U21335 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n21391), .ZN(MEM_stage_inst_dmem_n21372) );
NAND2_X1 MEM_stage_inst_dmem_U21334 ( .A1(MEM_stage_inst_dmem_ram_3641), .A2(MEM_stage_inst_dmem_n21390), .ZN(MEM_stage_inst_dmem_n21373) );
NAND2_X1 MEM_stage_inst_dmem_U21333 ( .A1(MEM_stage_inst_dmem_n21371), .A2(MEM_stage_inst_dmem_n21370), .ZN(MEM_stage_inst_dmem_n8821) );
NAND2_X1 MEM_stage_inst_dmem_U21332 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n21391), .ZN(MEM_stage_inst_dmem_n21370) );
NAND2_X1 MEM_stage_inst_dmem_U21331 ( .A1(MEM_stage_inst_dmem_ram_3642), .A2(MEM_stage_inst_dmem_n21390), .ZN(MEM_stage_inst_dmem_n21371) );
NAND2_X1 MEM_stage_inst_dmem_U21330 ( .A1(MEM_stage_inst_dmem_n21369), .A2(MEM_stage_inst_dmem_n21368), .ZN(MEM_stage_inst_dmem_n8822) );
NAND2_X1 MEM_stage_inst_dmem_U21329 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n21391), .ZN(MEM_stage_inst_dmem_n21368) );
NAND2_X1 MEM_stage_inst_dmem_U21328 ( .A1(MEM_stage_inst_dmem_ram_3643), .A2(MEM_stage_inst_dmem_n21390), .ZN(MEM_stage_inst_dmem_n21369) );
NAND2_X1 MEM_stage_inst_dmem_U21327 ( .A1(MEM_stage_inst_dmem_n21367), .A2(MEM_stage_inst_dmem_n21366), .ZN(MEM_stage_inst_dmem_n8823) );
NAND2_X1 MEM_stage_inst_dmem_U21326 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n21391), .ZN(MEM_stage_inst_dmem_n21366) );
NAND2_X1 MEM_stage_inst_dmem_U21325 ( .A1(MEM_stage_inst_dmem_ram_3644), .A2(MEM_stage_inst_dmem_n21390), .ZN(MEM_stage_inst_dmem_n21367) );
NAND2_X1 MEM_stage_inst_dmem_U21324 ( .A1(MEM_stage_inst_dmem_n21365), .A2(MEM_stage_inst_dmem_n21364), .ZN(MEM_stage_inst_dmem_n8824) );
NAND2_X1 MEM_stage_inst_dmem_U21323 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n21391), .ZN(MEM_stage_inst_dmem_n21364) );
NAND2_X1 MEM_stage_inst_dmem_U21322 ( .A1(MEM_stage_inst_dmem_ram_3645), .A2(MEM_stage_inst_dmem_n21390), .ZN(MEM_stage_inst_dmem_n21365) );
NAND2_X1 MEM_stage_inst_dmem_U21321 ( .A1(MEM_stage_inst_dmem_n21363), .A2(MEM_stage_inst_dmem_n21362), .ZN(MEM_stage_inst_dmem_n8825) );
NAND2_X1 MEM_stage_inst_dmem_U21320 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n21391), .ZN(MEM_stage_inst_dmem_n21362) );
NAND2_X1 MEM_stage_inst_dmem_U21319 ( .A1(MEM_stage_inst_dmem_ram_3646), .A2(MEM_stage_inst_dmem_n21390), .ZN(MEM_stage_inst_dmem_n21363) );
NAND2_X1 MEM_stage_inst_dmem_U21318 ( .A1(MEM_stage_inst_dmem_n21361), .A2(MEM_stage_inst_dmem_n21360), .ZN(MEM_stage_inst_dmem_n8826) );
NAND2_X1 MEM_stage_inst_dmem_U21317 ( .A1(MEM_stage_inst_dmem_n15110), .A2(MEM_stage_inst_dmem_n21391), .ZN(MEM_stage_inst_dmem_n21360) );
NAND2_X1 MEM_stage_inst_dmem_U21316 ( .A1(MEM_stage_inst_dmem_ram_3647), .A2(MEM_stage_inst_dmem_n21390), .ZN(MEM_stage_inst_dmem_n21361) );
NAND2_X1 MEM_stage_inst_dmem_U21315 ( .A1(MEM_stage_inst_dmem_n21359), .A2(MEM_stage_inst_dmem_n21464), .ZN(MEM_stage_inst_dmem_n21390) );
NAND2_X1 MEM_stage_inst_dmem_U21314 ( .A1(MEM_stage_inst_dmem_n21358), .A2(MEM_stage_inst_dmem_n21357), .ZN(MEM_stage_inst_dmem_n8827) );
NAND2_X1 MEM_stage_inst_dmem_U21313 ( .A1(EX_pipeline_reg_out_5), .A2(MEM_stage_inst_dmem_n21356), .ZN(MEM_stage_inst_dmem_n21357) );
NAND2_X1 MEM_stage_inst_dmem_U21312 ( .A1(MEM_stage_inst_dmem_ram_3648), .A2(MEM_stage_inst_dmem_n21355), .ZN(MEM_stage_inst_dmem_n21358) );
NAND2_X1 MEM_stage_inst_dmem_U21311 ( .A1(MEM_stage_inst_dmem_n21354), .A2(MEM_stage_inst_dmem_n21353), .ZN(MEM_stage_inst_dmem_n8828) );
NAND2_X1 MEM_stage_inst_dmem_U21310 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n21356), .ZN(MEM_stage_inst_dmem_n21353) );
NAND2_X1 MEM_stage_inst_dmem_U21309 ( .A1(MEM_stage_inst_dmem_ram_3649), .A2(MEM_stage_inst_dmem_n21355), .ZN(MEM_stage_inst_dmem_n21354) );
NAND2_X1 MEM_stage_inst_dmem_U21308 ( .A1(MEM_stage_inst_dmem_n21351), .A2(MEM_stage_inst_dmem_n21350), .ZN(MEM_stage_inst_dmem_n8829) );
NAND2_X1 MEM_stage_inst_dmem_U21307 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n21356), .ZN(MEM_stage_inst_dmem_n21350) );
NAND2_X1 MEM_stage_inst_dmem_U21306 ( .A1(MEM_stage_inst_dmem_ram_3650), .A2(MEM_stage_inst_dmem_n21355), .ZN(MEM_stage_inst_dmem_n21351) );
NAND2_X1 MEM_stage_inst_dmem_U21305 ( .A1(MEM_stage_inst_dmem_n21349), .A2(MEM_stage_inst_dmem_n21348), .ZN(MEM_stage_inst_dmem_n8830) );
NAND2_X1 MEM_stage_inst_dmem_U21304 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n21356), .ZN(MEM_stage_inst_dmem_n21348) );
NAND2_X1 MEM_stage_inst_dmem_U21303 ( .A1(MEM_stage_inst_dmem_ram_3651), .A2(MEM_stage_inst_dmem_n21355), .ZN(MEM_stage_inst_dmem_n21349) );
NAND2_X1 MEM_stage_inst_dmem_U21302 ( .A1(MEM_stage_inst_dmem_n21347), .A2(MEM_stage_inst_dmem_n21346), .ZN(MEM_stage_inst_dmem_n8831) );
NAND2_X1 MEM_stage_inst_dmem_U21301 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n21356), .ZN(MEM_stage_inst_dmem_n21346) );
NAND2_X1 MEM_stage_inst_dmem_U21300 ( .A1(MEM_stage_inst_dmem_ram_3652), .A2(MEM_stage_inst_dmem_n21355), .ZN(MEM_stage_inst_dmem_n21347) );
NAND2_X1 MEM_stage_inst_dmem_U21299 ( .A1(MEM_stage_inst_dmem_n21344), .A2(MEM_stage_inst_dmem_n21343), .ZN(MEM_stage_inst_dmem_n8832) );
NAND2_X1 MEM_stage_inst_dmem_U21298 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n21356), .ZN(MEM_stage_inst_dmem_n21343) );
NAND2_X1 MEM_stage_inst_dmem_U21297 ( .A1(MEM_stage_inst_dmem_ram_3653), .A2(MEM_stage_inst_dmem_n21355), .ZN(MEM_stage_inst_dmem_n21344) );
NAND2_X1 MEM_stage_inst_dmem_U21296 ( .A1(MEM_stage_inst_dmem_n21342), .A2(MEM_stage_inst_dmem_n21341), .ZN(MEM_stage_inst_dmem_n8833) );
NAND2_X1 MEM_stage_inst_dmem_U21295 ( .A1(MEM_stage_inst_dmem_n21340), .A2(MEM_stage_inst_dmem_n21356), .ZN(MEM_stage_inst_dmem_n21341) );
NAND2_X1 MEM_stage_inst_dmem_U21294 ( .A1(MEM_stage_inst_dmem_ram_3654), .A2(MEM_stage_inst_dmem_n21355), .ZN(MEM_stage_inst_dmem_n21342) );
NAND2_X1 MEM_stage_inst_dmem_U21293 ( .A1(MEM_stage_inst_dmem_n21339), .A2(MEM_stage_inst_dmem_n21338), .ZN(MEM_stage_inst_dmem_n8834) );
NAND2_X1 MEM_stage_inst_dmem_U21292 ( .A1(MEM_stage_inst_dmem_n17), .A2(MEM_stage_inst_dmem_n21356), .ZN(MEM_stage_inst_dmem_n21338) );
NAND2_X1 MEM_stage_inst_dmem_U21291 ( .A1(MEM_stage_inst_dmem_ram_3655), .A2(MEM_stage_inst_dmem_n21355), .ZN(MEM_stage_inst_dmem_n21339) );
NAND2_X1 MEM_stage_inst_dmem_U21290 ( .A1(MEM_stage_inst_dmem_n21337), .A2(MEM_stage_inst_dmem_n21336), .ZN(MEM_stage_inst_dmem_n8835) );
NAND2_X1 MEM_stage_inst_dmem_U21289 ( .A1(MEM_stage_inst_dmem_n21335), .A2(MEM_stage_inst_dmem_n21356), .ZN(MEM_stage_inst_dmem_n21336) );
NAND2_X1 MEM_stage_inst_dmem_U21288 ( .A1(MEM_stage_inst_dmem_ram_3656), .A2(MEM_stage_inst_dmem_n21355), .ZN(MEM_stage_inst_dmem_n21337) );
NAND2_X1 MEM_stage_inst_dmem_U21287 ( .A1(MEM_stage_inst_dmem_n21334), .A2(MEM_stage_inst_dmem_n21333), .ZN(MEM_stage_inst_dmem_n8836) );
NAND2_X1 MEM_stage_inst_dmem_U21286 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n21356), .ZN(MEM_stage_inst_dmem_n21333) );
NAND2_X1 MEM_stage_inst_dmem_U21285 ( .A1(MEM_stage_inst_dmem_ram_3657), .A2(MEM_stage_inst_dmem_n21355), .ZN(MEM_stage_inst_dmem_n21334) );
NAND2_X1 MEM_stage_inst_dmem_U21284 ( .A1(MEM_stage_inst_dmem_n21332), .A2(MEM_stage_inst_dmem_n21331), .ZN(MEM_stage_inst_dmem_n8837) );
NAND2_X1 MEM_stage_inst_dmem_U21283 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n21356), .ZN(MEM_stage_inst_dmem_n21331) );
NAND2_X1 MEM_stage_inst_dmem_U21282 ( .A1(MEM_stage_inst_dmem_ram_3658), .A2(MEM_stage_inst_dmem_n21355), .ZN(MEM_stage_inst_dmem_n21332) );
NAND2_X1 MEM_stage_inst_dmem_U21281 ( .A1(MEM_stage_inst_dmem_n21330), .A2(MEM_stage_inst_dmem_n21329), .ZN(MEM_stage_inst_dmem_n8838) );
NAND2_X1 MEM_stage_inst_dmem_U21280 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n21356), .ZN(MEM_stage_inst_dmem_n21329) );
NAND2_X1 MEM_stage_inst_dmem_U21279 ( .A1(MEM_stage_inst_dmem_ram_3659), .A2(MEM_stage_inst_dmem_n21355), .ZN(MEM_stage_inst_dmem_n21330) );
NAND2_X1 MEM_stage_inst_dmem_U21278 ( .A1(MEM_stage_inst_dmem_n21328), .A2(MEM_stage_inst_dmem_n21327), .ZN(MEM_stage_inst_dmem_n8839) );
NAND2_X1 MEM_stage_inst_dmem_U21277 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n21356), .ZN(MEM_stage_inst_dmem_n21327) );
NAND2_X1 MEM_stage_inst_dmem_U21276 ( .A1(MEM_stage_inst_dmem_ram_3660), .A2(MEM_stage_inst_dmem_n21355), .ZN(MEM_stage_inst_dmem_n21328) );
NAND2_X1 MEM_stage_inst_dmem_U21275 ( .A1(MEM_stage_inst_dmem_n21326), .A2(MEM_stage_inst_dmem_n21325), .ZN(MEM_stage_inst_dmem_n8840) );
NAND2_X1 MEM_stage_inst_dmem_U21274 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n21356), .ZN(MEM_stage_inst_dmem_n21325) );
NAND2_X1 MEM_stage_inst_dmem_U21273 ( .A1(MEM_stage_inst_dmem_ram_3661), .A2(MEM_stage_inst_dmem_n21355), .ZN(MEM_stage_inst_dmem_n21326) );
NAND2_X1 MEM_stage_inst_dmem_U21272 ( .A1(MEM_stage_inst_dmem_n21324), .A2(MEM_stage_inst_dmem_n21323), .ZN(MEM_stage_inst_dmem_n8841) );
NAND2_X1 MEM_stage_inst_dmem_U21271 ( .A1(EX_pipeline_reg_out_19), .A2(MEM_stage_inst_dmem_n21356), .ZN(MEM_stage_inst_dmem_n21323) );
NAND2_X1 MEM_stage_inst_dmem_U21270 ( .A1(MEM_stage_inst_dmem_ram_3662), .A2(MEM_stage_inst_dmem_n21355), .ZN(MEM_stage_inst_dmem_n21324) );
NAND2_X1 MEM_stage_inst_dmem_U21269 ( .A1(MEM_stage_inst_dmem_n21322), .A2(MEM_stage_inst_dmem_n21321), .ZN(MEM_stage_inst_dmem_n8842) );
NAND2_X1 MEM_stage_inst_dmem_U21268 ( .A1(MEM_stage_inst_dmem_n21320), .A2(MEM_stage_inst_dmem_n21356), .ZN(MEM_stage_inst_dmem_n21321) );
INV_X1 MEM_stage_inst_dmem_U21267 ( .A(MEM_stage_inst_dmem_n21355), .ZN(MEM_stage_inst_dmem_n21356) );
NAND2_X1 MEM_stage_inst_dmem_U21266 ( .A1(MEM_stage_inst_dmem_ram_3663), .A2(MEM_stage_inst_dmem_n21355), .ZN(MEM_stage_inst_dmem_n21322) );
NAND2_X1 MEM_stage_inst_dmem_U21265 ( .A1(MEM_stage_inst_dmem_n21319), .A2(MEM_stage_inst_dmem_n21464), .ZN(MEM_stage_inst_dmem_n21355) );
NAND2_X1 MEM_stage_inst_dmem_U21264 ( .A1(MEM_stage_inst_dmem_n21318), .A2(MEM_stage_inst_dmem_n21317), .ZN(MEM_stage_inst_dmem_n8843) );
NAND2_X1 MEM_stage_inst_dmem_U21263 ( .A1(MEM_stage_inst_dmem_n14732), .A2(MEM_stage_inst_dmem_n21316), .ZN(MEM_stage_inst_dmem_n21317) );
NAND2_X1 MEM_stage_inst_dmem_U21262 ( .A1(MEM_stage_inst_dmem_ram_3664), .A2(MEM_stage_inst_dmem_n21315), .ZN(MEM_stage_inst_dmem_n21318) );
NAND2_X1 MEM_stage_inst_dmem_U21261 ( .A1(MEM_stage_inst_dmem_n21314), .A2(MEM_stage_inst_dmem_n21313), .ZN(MEM_stage_inst_dmem_n8844) );
NAND2_X1 MEM_stage_inst_dmem_U21260 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n21316), .ZN(MEM_stage_inst_dmem_n21313) );
NAND2_X1 MEM_stage_inst_dmem_U21259 ( .A1(MEM_stage_inst_dmem_ram_3665), .A2(MEM_stage_inst_dmem_n21315), .ZN(MEM_stage_inst_dmem_n21314) );
NAND2_X1 MEM_stage_inst_dmem_U21258 ( .A1(MEM_stage_inst_dmem_n21312), .A2(MEM_stage_inst_dmem_n21311), .ZN(MEM_stage_inst_dmem_n8845) );
NAND2_X1 MEM_stage_inst_dmem_U21257 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n21316), .ZN(MEM_stage_inst_dmem_n21311) );
NAND2_X1 MEM_stage_inst_dmem_U21256 ( .A1(MEM_stage_inst_dmem_ram_3666), .A2(MEM_stage_inst_dmem_n21315), .ZN(MEM_stage_inst_dmem_n21312) );
NAND2_X1 MEM_stage_inst_dmem_U21255 ( .A1(MEM_stage_inst_dmem_n21310), .A2(MEM_stage_inst_dmem_n21309), .ZN(MEM_stage_inst_dmem_n8846) );
NAND2_X1 MEM_stage_inst_dmem_U21254 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n21316), .ZN(MEM_stage_inst_dmem_n21309) );
NAND2_X1 MEM_stage_inst_dmem_U21253 ( .A1(MEM_stage_inst_dmem_ram_3667), .A2(MEM_stage_inst_dmem_n21315), .ZN(MEM_stage_inst_dmem_n21310) );
NAND2_X1 MEM_stage_inst_dmem_U21252 ( .A1(MEM_stage_inst_dmem_n21308), .A2(MEM_stage_inst_dmem_n21307), .ZN(MEM_stage_inst_dmem_n8847) );
NAND2_X1 MEM_stage_inst_dmem_U21251 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n21316), .ZN(MEM_stage_inst_dmem_n21307) );
NAND2_X1 MEM_stage_inst_dmem_U21250 ( .A1(MEM_stage_inst_dmem_ram_3668), .A2(MEM_stage_inst_dmem_n21315), .ZN(MEM_stage_inst_dmem_n21308) );
NAND2_X1 MEM_stage_inst_dmem_U21249 ( .A1(MEM_stage_inst_dmem_n21306), .A2(MEM_stage_inst_dmem_n21305), .ZN(MEM_stage_inst_dmem_n8848) );
NAND2_X1 MEM_stage_inst_dmem_U21248 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n21316), .ZN(MEM_stage_inst_dmem_n21305) );
NAND2_X1 MEM_stage_inst_dmem_U21247 ( .A1(MEM_stage_inst_dmem_ram_3669), .A2(MEM_stage_inst_dmem_n21315), .ZN(MEM_stage_inst_dmem_n21306) );
NAND2_X1 MEM_stage_inst_dmem_U21246 ( .A1(MEM_stage_inst_dmem_n21304), .A2(MEM_stage_inst_dmem_n21303), .ZN(MEM_stage_inst_dmem_n8849) );
NAND2_X1 MEM_stage_inst_dmem_U21245 ( .A1(MEM_stage_inst_dmem_n21340), .A2(MEM_stage_inst_dmem_n21316), .ZN(MEM_stage_inst_dmem_n21303) );
NAND2_X1 MEM_stage_inst_dmem_U21244 ( .A1(MEM_stage_inst_dmem_ram_3670), .A2(MEM_stage_inst_dmem_n21315), .ZN(MEM_stage_inst_dmem_n21304) );
NAND2_X1 MEM_stage_inst_dmem_U21243 ( .A1(MEM_stage_inst_dmem_n21302), .A2(MEM_stage_inst_dmem_n21301), .ZN(MEM_stage_inst_dmem_n8850) );
NAND2_X1 MEM_stage_inst_dmem_U21242 ( .A1(MEM_stage_inst_dmem_n18), .A2(MEM_stage_inst_dmem_n21316), .ZN(MEM_stage_inst_dmem_n21301) );
NAND2_X1 MEM_stage_inst_dmem_U21241 ( .A1(MEM_stage_inst_dmem_ram_3671), .A2(MEM_stage_inst_dmem_n21315), .ZN(MEM_stage_inst_dmem_n21302) );
NAND2_X1 MEM_stage_inst_dmem_U21240 ( .A1(MEM_stage_inst_dmem_n21300), .A2(MEM_stage_inst_dmem_n21299), .ZN(MEM_stage_inst_dmem_n8851) );
NAND2_X1 MEM_stage_inst_dmem_U21239 ( .A1(MEM_stage_inst_dmem_n21335), .A2(MEM_stage_inst_dmem_n21316), .ZN(MEM_stage_inst_dmem_n21299) );
NAND2_X1 MEM_stage_inst_dmem_U21238 ( .A1(MEM_stage_inst_dmem_ram_3672), .A2(MEM_stage_inst_dmem_n21315), .ZN(MEM_stage_inst_dmem_n21300) );
NAND2_X1 MEM_stage_inst_dmem_U21237 ( .A1(MEM_stage_inst_dmem_n21298), .A2(MEM_stage_inst_dmem_n21297), .ZN(MEM_stage_inst_dmem_n8852) );
NAND2_X1 MEM_stage_inst_dmem_U21236 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n21316), .ZN(MEM_stage_inst_dmem_n21297) );
NAND2_X1 MEM_stage_inst_dmem_U21235 ( .A1(MEM_stage_inst_dmem_ram_3673), .A2(MEM_stage_inst_dmem_n21315), .ZN(MEM_stage_inst_dmem_n21298) );
NAND2_X1 MEM_stage_inst_dmem_U21234 ( .A1(MEM_stage_inst_dmem_n21296), .A2(MEM_stage_inst_dmem_n21295), .ZN(MEM_stage_inst_dmem_n8853) );
NAND2_X1 MEM_stage_inst_dmem_U21233 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n21316), .ZN(MEM_stage_inst_dmem_n21295) );
NAND2_X1 MEM_stage_inst_dmem_U21232 ( .A1(MEM_stage_inst_dmem_ram_3674), .A2(MEM_stage_inst_dmem_n21315), .ZN(MEM_stage_inst_dmem_n21296) );
NAND2_X1 MEM_stage_inst_dmem_U21231 ( .A1(MEM_stage_inst_dmem_n21294), .A2(MEM_stage_inst_dmem_n21293), .ZN(MEM_stage_inst_dmem_n8854) );
NAND2_X1 MEM_stage_inst_dmem_U21230 ( .A1(MEM_stage_inst_dmem_n20904), .A2(MEM_stage_inst_dmem_n21316), .ZN(MEM_stage_inst_dmem_n21293) );
NAND2_X1 MEM_stage_inst_dmem_U21229 ( .A1(MEM_stage_inst_dmem_ram_3675), .A2(MEM_stage_inst_dmem_n21315), .ZN(MEM_stage_inst_dmem_n21294) );
NAND2_X1 MEM_stage_inst_dmem_U21228 ( .A1(MEM_stage_inst_dmem_n21292), .A2(MEM_stage_inst_dmem_n21291), .ZN(MEM_stage_inst_dmem_n8855) );
NAND2_X1 MEM_stage_inst_dmem_U21227 ( .A1(MEM_stage_inst_dmem_n21474), .A2(MEM_stage_inst_dmem_n21316), .ZN(MEM_stage_inst_dmem_n21291) );
NAND2_X1 MEM_stage_inst_dmem_U21226 ( .A1(MEM_stage_inst_dmem_ram_3676), .A2(MEM_stage_inst_dmem_n21315), .ZN(MEM_stage_inst_dmem_n21292) );
NAND2_X1 MEM_stage_inst_dmem_U21225 ( .A1(MEM_stage_inst_dmem_n21290), .A2(MEM_stage_inst_dmem_n21289), .ZN(MEM_stage_inst_dmem_n8856) );
NAND2_X1 MEM_stage_inst_dmem_U21224 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n21316), .ZN(MEM_stage_inst_dmem_n21289) );
NAND2_X1 MEM_stage_inst_dmem_U21223 ( .A1(MEM_stage_inst_dmem_ram_3677), .A2(MEM_stage_inst_dmem_n21315), .ZN(MEM_stage_inst_dmem_n21290) );
NAND2_X1 MEM_stage_inst_dmem_U21222 ( .A1(MEM_stage_inst_dmem_n21288), .A2(MEM_stage_inst_dmem_n21287), .ZN(MEM_stage_inst_dmem_n8857) );
NAND2_X1 MEM_stage_inst_dmem_U21221 ( .A1(MEM_stage_inst_dmem_n14696), .A2(MEM_stage_inst_dmem_n21316), .ZN(MEM_stage_inst_dmem_n21287) );
NAND2_X1 MEM_stage_inst_dmem_U21220 ( .A1(MEM_stage_inst_dmem_ram_3678), .A2(MEM_stage_inst_dmem_n21315), .ZN(MEM_stage_inst_dmem_n21288) );
NAND2_X1 MEM_stage_inst_dmem_U21219 ( .A1(MEM_stage_inst_dmem_n21286), .A2(MEM_stage_inst_dmem_n21285), .ZN(MEM_stage_inst_dmem_n8858) );
NAND2_X1 MEM_stage_inst_dmem_U21218 ( .A1(MEM_stage_inst_dmem_n21320), .A2(MEM_stage_inst_dmem_n21316), .ZN(MEM_stage_inst_dmem_n21285) );
INV_X1 MEM_stage_inst_dmem_U21217 ( .A(MEM_stage_inst_dmem_n21315), .ZN(MEM_stage_inst_dmem_n21316) );
NAND2_X1 MEM_stage_inst_dmem_U21216 ( .A1(MEM_stage_inst_dmem_ram_3679), .A2(MEM_stage_inst_dmem_n21315), .ZN(MEM_stage_inst_dmem_n21286) );
NAND2_X1 MEM_stage_inst_dmem_U21215 ( .A1(MEM_stage_inst_dmem_n21284), .A2(MEM_stage_inst_dmem_n21464), .ZN(MEM_stage_inst_dmem_n21315) );
NAND2_X1 MEM_stage_inst_dmem_U21214 ( .A1(MEM_stage_inst_dmem_n21283), .A2(MEM_stage_inst_dmem_n21282), .ZN(MEM_stage_inst_dmem_n8859) );
NAND2_X1 MEM_stage_inst_dmem_U21213 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n21281), .ZN(MEM_stage_inst_dmem_n21282) );
NAND2_X1 MEM_stage_inst_dmem_U21212 ( .A1(MEM_stage_inst_dmem_ram_3680), .A2(MEM_stage_inst_dmem_n21280), .ZN(MEM_stage_inst_dmem_n21283) );
NAND2_X1 MEM_stage_inst_dmem_U21211 ( .A1(MEM_stage_inst_dmem_n21279), .A2(MEM_stage_inst_dmem_n21278), .ZN(MEM_stage_inst_dmem_n8860) );
NAND2_X1 MEM_stage_inst_dmem_U21210 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n21281), .ZN(MEM_stage_inst_dmem_n21278) );
NAND2_X1 MEM_stage_inst_dmem_U21209 ( .A1(MEM_stage_inst_dmem_ram_3681), .A2(MEM_stage_inst_dmem_n21280), .ZN(MEM_stage_inst_dmem_n21279) );
NAND2_X1 MEM_stage_inst_dmem_U21208 ( .A1(MEM_stage_inst_dmem_n21277), .A2(MEM_stage_inst_dmem_n21276), .ZN(MEM_stage_inst_dmem_n8861) );
NAND2_X1 MEM_stage_inst_dmem_U21207 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n21281), .ZN(MEM_stage_inst_dmem_n21276) );
NAND2_X1 MEM_stage_inst_dmem_U21206 ( .A1(MEM_stage_inst_dmem_ram_3682), .A2(MEM_stage_inst_dmem_n21280), .ZN(MEM_stage_inst_dmem_n21277) );
NAND2_X1 MEM_stage_inst_dmem_U21205 ( .A1(MEM_stage_inst_dmem_n21275), .A2(MEM_stage_inst_dmem_n21274), .ZN(MEM_stage_inst_dmem_n8862) );
NAND2_X1 MEM_stage_inst_dmem_U21204 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n21281), .ZN(MEM_stage_inst_dmem_n21274) );
NAND2_X1 MEM_stage_inst_dmem_U21203 ( .A1(MEM_stage_inst_dmem_ram_3683), .A2(MEM_stage_inst_dmem_n21280), .ZN(MEM_stage_inst_dmem_n21275) );
NAND2_X1 MEM_stage_inst_dmem_U21202 ( .A1(MEM_stage_inst_dmem_n21273), .A2(MEM_stage_inst_dmem_n21272), .ZN(MEM_stage_inst_dmem_n8863) );
NAND2_X1 MEM_stage_inst_dmem_U21201 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n21281), .ZN(MEM_stage_inst_dmem_n21272) );
NAND2_X1 MEM_stage_inst_dmem_U21200 ( .A1(MEM_stage_inst_dmem_ram_3684), .A2(MEM_stage_inst_dmem_n21280), .ZN(MEM_stage_inst_dmem_n21273) );
NAND2_X1 MEM_stage_inst_dmem_U21199 ( .A1(MEM_stage_inst_dmem_n21271), .A2(MEM_stage_inst_dmem_n21270), .ZN(MEM_stage_inst_dmem_n8864) );
NAND2_X1 MEM_stage_inst_dmem_U21198 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n21281), .ZN(MEM_stage_inst_dmem_n21270) );
NAND2_X1 MEM_stage_inst_dmem_U21197 ( .A1(MEM_stage_inst_dmem_ram_3685), .A2(MEM_stage_inst_dmem_n21280), .ZN(MEM_stage_inst_dmem_n21271) );
NAND2_X1 MEM_stage_inst_dmem_U21196 ( .A1(MEM_stage_inst_dmem_n21269), .A2(MEM_stage_inst_dmem_n21268), .ZN(MEM_stage_inst_dmem_n8865) );
NAND2_X1 MEM_stage_inst_dmem_U21195 ( .A1(MEM_stage_inst_dmem_n21340), .A2(MEM_stage_inst_dmem_n21281), .ZN(MEM_stage_inst_dmem_n21268) );
NAND2_X1 MEM_stage_inst_dmem_U21194 ( .A1(MEM_stage_inst_dmem_ram_3686), .A2(MEM_stage_inst_dmem_n21280), .ZN(MEM_stage_inst_dmem_n21269) );
NAND2_X1 MEM_stage_inst_dmem_U21193 ( .A1(MEM_stage_inst_dmem_n21267), .A2(MEM_stage_inst_dmem_n21266), .ZN(MEM_stage_inst_dmem_n8866) );
NAND2_X1 MEM_stage_inst_dmem_U21192 ( .A1(MEM_stage_inst_dmem_n17), .A2(MEM_stage_inst_dmem_n21281), .ZN(MEM_stage_inst_dmem_n21266) );
NAND2_X1 MEM_stage_inst_dmem_U21191 ( .A1(MEM_stage_inst_dmem_ram_3687), .A2(MEM_stage_inst_dmem_n21280), .ZN(MEM_stage_inst_dmem_n21267) );
NAND2_X1 MEM_stage_inst_dmem_U21190 ( .A1(MEM_stage_inst_dmem_n21265), .A2(MEM_stage_inst_dmem_n21264), .ZN(MEM_stage_inst_dmem_n8867) );
NAND2_X1 MEM_stage_inst_dmem_U21189 ( .A1(MEM_stage_inst_dmem_n21335), .A2(MEM_stage_inst_dmem_n21281), .ZN(MEM_stage_inst_dmem_n21264) );
NAND2_X1 MEM_stage_inst_dmem_U21188 ( .A1(MEM_stage_inst_dmem_ram_3688), .A2(MEM_stage_inst_dmem_n21280), .ZN(MEM_stage_inst_dmem_n21265) );
NAND2_X1 MEM_stage_inst_dmem_U21187 ( .A1(MEM_stage_inst_dmem_n21263), .A2(MEM_stage_inst_dmem_n21262), .ZN(MEM_stage_inst_dmem_n8868) );
NAND2_X1 MEM_stage_inst_dmem_U21186 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n21281), .ZN(MEM_stage_inst_dmem_n21262) );
NAND2_X1 MEM_stage_inst_dmem_U21185 ( .A1(MEM_stage_inst_dmem_ram_3689), .A2(MEM_stage_inst_dmem_n21280), .ZN(MEM_stage_inst_dmem_n21263) );
NAND2_X1 MEM_stage_inst_dmem_U21184 ( .A1(MEM_stage_inst_dmem_n21261), .A2(MEM_stage_inst_dmem_n21260), .ZN(MEM_stage_inst_dmem_n8869) );
NAND2_X1 MEM_stage_inst_dmem_U21183 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n21281), .ZN(MEM_stage_inst_dmem_n21260) );
NAND2_X1 MEM_stage_inst_dmem_U21182 ( .A1(MEM_stage_inst_dmem_ram_3690), .A2(MEM_stage_inst_dmem_n21280), .ZN(MEM_stage_inst_dmem_n21261) );
NAND2_X1 MEM_stage_inst_dmem_U21181 ( .A1(MEM_stage_inst_dmem_n21259), .A2(MEM_stage_inst_dmem_n21258), .ZN(MEM_stage_inst_dmem_n8870) );
NAND2_X1 MEM_stage_inst_dmem_U21180 ( .A1(MEM_stage_inst_dmem_n13044), .A2(MEM_stage_inst_dmem_n21281), .ZN(MEM_stage_inst_dmem_n21258) );
NAND2_X1 MEM_stage_inst_dmem_U21179 ( .A1(MEM_stage_inst_dmem_ram_3691), .A2(MEM_stage_inst_dmem_n21280), .ZN(MEM_stage_inst_dmem_n21259) );
NAND2_X1 MEM_stage_inst_dmem_U21178 ( .A1(MEM_stage_inst_dmem_n21257), .A2(MEM_stage_inst_dmem_n21256), .ZN(MEM_stage_inst_dmem_n8871) );
NAND2_X1 MEM_stage_inst_dmem_U21177 ( .A1(MEM_stage_inst_dmem_n13041), .A2(MEM_stage_inst_dmem_n21281), .ZN(MEM_stage_inst_dmem_n21256) );
NAND2_X1 MEM_stage_inst_dmem_U21176 ( .A1(MEM_stage_inst_dmem_ram_3692), .A2(MEM_stage_inst_dmem_n21280), .ZN(MEM_stage_inst_dmem_n21257) );
NAND2_X1 MEM_stage_inst_dmem_U21175 ( .A1(MEM_stage_inst_dmem_n21255), .A2(MEM_stage_inst_dmem_n21254), .ZN(MEM_stage_inst_dmem_n8872) );
NAND2_X1 MEM_stage_inst_dmem_U21174 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n21281), .ZN(MEM_stage_inst_dmem_n21254) );
NAND2_X1 MEM_stage_inst_dmem_U21173 ( .A1(MEM_stage_inst_dmem_ram_3693), .A2(MEM_stage_inst_dmem_n21280), .ZN(MEM_stage_inst_dmem_n21255) );
NAND2_X1 MEM_stage_inst_dmem_U21172 ( .A1(MEM_stage_inst_dmem_n21253), .A2(MEM_stage_inst_dmem_n21252), .ZN(MEM_stage_inst_dmem_n8873) );
NAND2_X1 MEM_stage_inst_dmem_U21171 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n21281), .ZN(MEM_stage_inst_dmem_n21252) );
NAND2_X1 MEM_stage_inst_dmem_U21170 ( .A1(MEM_stage_inst_dmem_ram_3694), .A2(MEM_stage_inst_dmem_n21280), .ZN(MEM_stage_inst_dmem_n21253) );
NAND2_X1 MEM_stage_inst_dmem_U21169 ( .A1(MEM_stage_inst_dmem_n21251), .A2(MEM_stage_inst_dmem_n21250), .ZN(MEM_stage_inst_dmem_n8874) );
NAND2_X1 MEM_stage_inst_dmem_U21168 ( .A1(MEM_stage_inst_dmem_n21320), .A2(MEM_stage_inst_dmem_n21281), .ZN(MEM_stage_inst_dmem_n21250) );
INV_X1 MEM_stage_inst_dmem_U21167 ( .A(MEM_stage_inst_dmem_n21280), .ZN(MEM_stage_inst_dmem_n21281) );
NAND2_X1 MEM_stage_inst_dmem_U21166 ( .A1(MEM_stage_inst_dmem_ram_3695), .A2(MEM_stage_inst_dmem_n21280), .ZN(MEM_stage_inst_dmem_n21251) );
NAND2_X1 MEM_stage_inst_dmem_U21165 ( .A1(MEM_stage_inst_dmem_n21249), .A2(MEM_stage_inst_dmem_n21464), .ZN(MEM_stage_inst_dmem_n21280) );
NAND2_X1 MEM_stage_inst_dmem_U21164 ( .A1(MEM_stage_inst_dmem_n21248), .A2(MEM_stage_inst_dmem_n21247), .ZN(MEM_stage_inst_dmem_n8875) );
NAND2_X1 MEM_stage_inst_dmem_U21163 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n21246), .ZN(MEM_stage_inst_dmem_n21247) );
NAND2_X1 MEM_stage_inst_dmem_U21162 ( .A1(MEM_stage_inst_dmem_ram_3696), .A2(MEM_stage_inst_dmem_n21245), .ZN(MEM_stage_inst_dmem_n21248) );
NAND2_X1 MEM_stage_inst_dmem_U21161 ( .A1(MEM_stage_inst_dmem_n21244), .A2(MEM_stage_inst_dmem_n21243), .ZN(MEM_stage_inst_dmem_n8876) );
NAND2_X1 MEM_stage_inst_dmem_U21160 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n21246), .ZN(MEM_stage_inst_dmem_n21243) );
NAND2_X1 MEM_stage_inst_dmem_U21159 ( .A1(MEM_stage_inst_dmem_ram_3697), .A2(MEM_stage_inst_dmem_n21245), .ZN(MEM_stage_inst_dmem_n21244) );
NAND2_X1 MEM_stage_inst_dmem_U21158 ( .A1(MEM_stage_inst_dmem_n21242), .A2(MEM_stage_inst_dmem_n21241), .ZN(MEM_stage_inst_dmem_n8877) );
NAND2_X1 MEM_stage_inst_dmem_U21157 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n21246), .ZN(MEM_stage_inst_dmem_n21241) );
NAND2_X1 MEM_stage_inst_dmem_U21156 ( .A1(MEM_stage_inst_dmem_ram_3698), .A2(MEM_stage_inst_dmem_n21245), .ZN(MEM_stage_inst_dmem_n21242) );
NAND2_X1 MEM_stage_inst_dmem_U21155 ( .A1(MEM_stage_inst_dmem_n21240), .A2(MEM_stage_inst_dmem_n21239), .ZN(MEM_stage_inst_dmem_n8878) );
NAND2_X1 MEM_stage_inst_dmem_U21154 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n21246), .ZN(MEM_stage_inst_dmem_n21239) );
NAND2_X1 MEM_stage_inst_dmem_U21153 ( .A1(MEM_stage_inst_dmem_ram_3699), .A2(MEM_stage_inst_dmem_n21245), .ZN(MEM_stage_inst_dmem_n21240) );
NAND2_X1 MEM_stage_inst_dmem_U21152 ( .A1(MEM_stage_inst_dmem_n21238), .A2(MEM_stage_inst_dmem_n21237), .ZN(MEM_stage_inst_dmem_n8879) );
NAND2_X1 MEM_stage_inst_dmem_U21151 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n21246), .ZN(MEM_stage_inst_dmem_n21237) );
NAND2_X1 MEM_stage_inst_dmem_U21150 ( .A1(MEM_stage_inst_dmem_ram_3700), .A2(MEM_stage_inst_dmem_n21245), .ZN(MEM_stage_inst_dmem_n21238) );
NAND2_X1 MEM_stage_inst_dmem_U21149 ( .A1(MEM_stage_inst_dmem_n21236), .A2(MEM_stage_inst_dmem_n21235), .ZN(MEM_stage_inst_dmem_n8880) );
NAND2_X1 MEM_stage_inst_dmem_U21148 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n21246), .ZN(MEM_stage_inst_dmem_n21235) );
NAND2_X1 MEM_stage_inst_dmem_U21147 ( .A1(MEM_stage_inst_dmem_ram_3701), .A2(MEM_stage_inst_dmem_n21245), .ZN(MEM_stage_inst_dmem_n21236) );
NAND2_X1 MEM_stage_inst_dmem_U21146 ( .A1(MEM_stage_inst_dmem_n21234), .A2(MEM_stage_inst_dmem_n21233), .ZN(MEM_stage_inst_dmem_n8881) );
NAND2_X1 MEM_stage_inst_dmem_U21145 ( .A1(MEM_stage_inst_dmem_n21340), .A2(MEM_stage_inst_dmem_n21246), .ZN(MEM_stage_inst_dmem_n21233) );
NAND2_X1 MEM_stage_inst_dmem_U21144 ( .A1(MEM_stage_inst_dmem_ram_3702), .A2(MEM_stage_inst_dmem_n21245), .ZN(MEM_stage_inst_dmem_n21234) );
NAND2_X1 MEM_stage_inst_dmem_U21143 ( .A1(MEM_stage_inst_dmem_n21232), .A2(MEM_stage_inst_dmem_n21231), .ZN(MEM_stage_inst_dmem_n8882) );
NAND2_X1 MEM_stage_inst_dmem_U21142 ( .A1(MEM_stage_inst_dmem_n18), .A2(MEM_stage_inst_dmem_n21246), .ZN(MEM_stage_inst_dmem_n21231) );
NAND2_X1 MEM_stage_inst_dmem_U21141 ( .A1(MEM_stage_inst_dmem_ram_3703), .A2(MEM_stage_inst_dmem_n21245), .ZN(MEM_stage_inst_dmem_n21232) );
NAND2_X1 MEM_stage_inst_dmem_U21140 ( .A1(MEM_stage_inst_dmem_n21230), .A2(MEM_stage_inst_dmem_n21229), .ZN(MEM_stage_inst_dmem_n8883) );
NAND2_X1 MEM_stage_inst_dmem_U21139 ( .A1(MEM_stage_inst_dmem_n21335), .A2(MEM_stage_inst_dmem_n21246), .ZN(MEM_stage_inst_dmem_n21229) );
NAND2_X1 MEM_stage_inst_dmem_U21138 ( .A1(MEM_stage_inst_dmem_ram_3704), .A2(MEM_stage_inst_dmem_n21245), .ZN(MEM_stage_inst_dmem_n21230) );
NAND2_X1 MEM_stage_inst_dmem_U21137 ( .A1(MEM_stage_inst_dmem_n21228), .A2(MEM_stage_inst_dmem_n21227), .ZN(MEM_stage_inst_dmem_n8884) );
NAND2_X1 MEM_stage_inst_dmem_U21136 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n21246), .ZN(MEM_stage_inst_dmem_n21227) );
NAND2_X1 MEM_stage_inst_dmem_U21135 ( .A1(MEM_stage_inst_dmem_ram_3705), .A2(MEM_stage_inst_dmem_n21245), .ZN(MEM_stage_inst_dmem_n21228) );
NAND2_X1 MEM_stage_inst_dmem_U21134 ( .A1(MEM_stage_inst_dmem_n21226), .A2(MEM_stage_inst_dmem_n21225), .ZN(MEM_stage_inst_dmem_n8885) );
NAND2_X1 MEM_stage_inst_dmem_U21133 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n21246), .ZN(MEM_stage_inst_dmem_n21225) );
NAND2_X1 MEM_stage_inst_dmem_U21132 ( .A1(MEM_stage_inst_dmem_ram_3706), .A2(MEM_stage_inst_dmem_n21245), .ZN(MEM_stage_inst_dmem_n21226) );
NAND2_X1 MEM_stage_inst_dmem_U21131 ( .A1(MEM_stage_inst_dmem_n21224), .A2(MEM_stage_inst_dmem_n21223), .ZN(MEM_stage_inst_dmem_n8886) );
NAND2_X1 MEM_stage_inst_dmem_U21130 ( .A1(MEM_stage_inst_dmem_n13044), .A2(MEM_stage_inst_dmem_n21246), .ZN(MEM_stage_inst_dmem_n21223) );
NAND2_X1 MEM_stage_inst_dmem_U21129 ( .A1(MEM_stage_inst_dmem_ram_3707), .A2(MEM_stage_inst_dmem_n21245), .ZN(MEM_stage_inst_dmem_n21224) );
NAND2_X1 MEM_stage_inst_dmem_U21128 ( .A1(MEM_stage_inst_dmem_n21222), .A2(MEM_stage_inst_dmem_n21221), .ZN(MEM_stage_inst_dmem_n8887) );
NAND2_X1 MEM_stage_inst_dmem_U21127 ( .A1(MEM_stage_inst_dmem_n13041), .A2(MEM_stage_inst_dmem_n21246), .ZN(MEM_stage_inst_dmem_n21221) );
NAND2_X1 MEM_stage_inst_dmem_U21126 ( .A1(MEM_stage_inst_dmem_ram_3708), .A2(MEM_stage_inst_dmem_n21245), .ZN(MEM_stage_inst_dmem_n21222) );
NAND2_X1 MEM_stage_inst_dmem_U21125 ( .A1(MEM_stage_inst_dmem_n21220), .A2(MEM_stage_inst_dmem_n21219), .ZN(MEM_stage_inst_dmem_n8888) );
NAND2_X1 MEM_stage_inst_dmem_U21124 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n21246), .ZN(MEM_stage_inst_dmem_n21219) );
NAND2_X1 MEM_stage_inst_dmem_U21123 ( .A1(MEM_stage_inst_dmem_ram_3709), .A2(MEM_stage_inst_dmem_n21245), .ZN(MEM_stage_inst_dmem_n21220) );
NAND2_X1 MEM_stage_inst_dmem_U21122 ( .A1(MEM_stage_inst_dmem_n21218), .A2(MEM_stage_inst_dmem_n21217), .ZN(MEM_stage_inst_dmem_n8889) );
NAND2_X1 MEM_stage_inst_dmem_U21121 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n21246), .ZN(MEM_stage_inst_dmem_n21217) );
NAND2_X1 MEM_stage_inst_dmem_U21120 ( .A1(MEM_stage_inst_dmem_ram_3710), .A2(MEM_stage_inst_dmem_n21245), .ZN(MEM_stage_inst_dmem_n21218) );
NAND2_X1 MEM_stage_inst_dmem_U21119 ( .A1(MEM_stage_inst_dmem_n21216), .A2(MEM_stage_inst_dmem_n21215), .ZN(MEM_stage_inst_dmem_n8890) );
NAND2_X1 MEM_stage_inst_dmem_U21118 ( .A1(MEM_stage_inst_dmem_n21320), .A2(MEM_stage_inst_dmem_n21246), .ZN(MEM_stage_inst_dmem_n21215) );
INV_X1 MEM_stage_inst_dmem_U21117 ( .A(MEM_stage_inst_dmem_n21245), .ZN(MEM_stage_inst_dmem_n21246) );
NAND2_X1 MEM_stage_inst_dmem_U21116 ( .A1(MEM_stage_inst_dmem_ram_3711), .A2(MEM_stage_inst_dmem_n21245), .ZN(MEM_stage_inst_dmem_n21216) );
NAND2_X1 MEM_stage_inst_dmem_U21115 ( .A1(MEM_stage_inst_dmem_n21214), .A2(MEM_stage_inst_dmem_n21464), .ZN(MEM_stage_inst_dmem_n21245) );
NAND2_X1 MEM_stage_inst_dmem_U21114 ( .A1(MEM_stage_inst_dmem_n21213), .A2(MEM_stage_inst_dmem_n21212), .ZN(MEM_stage_inst_dmem_n8891) );
NAND2_X1 MEM_stage_inst_dmem_U21113 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n21211), .ZN(MEM_stage_inst_dmem_n21212) );
NAND2_X1 MEM_stage_inst_dmem_U21112 ( .A1(MEM_stage_inst_dmem_ram_3712), .A2(MEM_stage_inst_dmem_n21210), .ZN(MEM_stage_inst_dmem_n21213) );
NAND2_X1 MEM_stage_inst_dmem_U21111 ( .A1(MEM_stage_inst_dmem_n21209), .A2(MEM_stage_inst_dmem_n21208), .ZN(MEM_stage_inst_dmem_n8892) );
NAND2_X1 MEM_stage_inst_dmem_U21110 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n21211), .ZN(MEM_stage_inst_dmem_n21208) );
NAND2_X1 MEM_stage_inst_dmem_U21109 ( .A1(MEM_stage_inst_dmem_ram_3713), .A2(MEM_stage_inst_dmem_n21210), .ZN(MEM_stage_inst_dmem_n21209) );
NAND2_X1 MEM_stage_inst_dmem_U21108 ( .A1(MEM_stage_inst_dmem_n21207), .A2(MEM_stage_inst_dmem_n21206), .ZN(MEM_stage_inst_dmem_n8893) );
NAND2_X1 MEM_stage_inst_dmem_U21107 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n21211), .ZN(MEM_stage_inst_dmem_n21206) );
NAND2_X1 MEM_stage_inst_dmem_U21106 ( .A1(MEM_stage_inst_dmem_ram_3714), .A2(MEM_stage_inst_dmem_n21210), .ZN(MEM_stage_inst_dmem_n21207) );
NAND2_X1 MEM_stage_inst_dmem_U21105 ( .A1(MEM_stage_inst_dmem_n21205), .A2(MEM_stage_inst_dmem_n21204), .ZN(MEM_stage_inst_dmem_n8894) );
NAND2_X1 MEM_stage_inst_dmem_U21104 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n21211), .ZN(MEM_stage_inst_dmem_n21204) );
NAND2_X1 MEM_stage_inst_dmem_U21103 ( .A1(MEM_stage_inst_dmem_ram_3715), .A2(MEM_stage_inst_dmem_n21210), .ZN(MEM_stage_inst_dmem_n21205) );
NAND2_X1 MEM_stage_inst_dmem_U21102 ( .A1(MEM_stage_inst_dmem_n21203), .A2(MEM_stage_inst_dmem_n21202), .ZN(MEM_stage_inst_dmem_n8895) );
NAND2_X1 MEM_stage_inst_dmem_U21101 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n21211), .ZN(MEM_stage_inst_dmem_n21202) );
NAND2_X1 MEM_stage_inst_dmem_U21100 ( .A1(MEM_stage_inst_dmem_ram_3716), .A2(MEM_stage_inst_dmem_n21210), .ZN(MEM_stage_inst_dmem_n21203) );
NAND2_X1 MEM_stage_inst_dmem_U21099 ( .A1(MEM_stage_inst_dmem_n21201), .A2(MEM_stage_inst_dmem_n21200), .ZN(MEM_stage_inst_dmem_n8896) );
NAND2_X1 MEM_stage_inst_dmem_U21098 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n21211), .ZN(MEM_stage_inst_dmem_n21200) );
NAND2_X1 MEM_stage_inst_dmem_U21097 ( .A1(MEM_stage_inst_dmem_ram_3717), .A2(MEM_stage_inst_dmem_n21210), .ZN(MEM_stage_inst_dmem_n21201) );
NAND2_X1 MEM_stage_inst_dmem_U21096 ( .A1(MEM_stage_inst_dmem_n21199), .A2(MEM_stage_inst_dmem_n21198), .ZN(MEM_stage_inst_dmem_n8897) );
NAND2_X1 MEM_stage_inst_dmem_U21095 ( .A1(MEM_stage_inst_dmem_n21340), .A2(MEM_stage_inst_dmem_n21211), .ZN(MEM_stage_inst_dmem_n21198) );
NAND2_X1 MEM_stage_inst_dmem_U21094 ( .A1(MEM_stage_inst_dmem_ram_3718), .A2(MEM_stage_inst_dmem_n21210), .ZN(MEM_stage_inst_dmem_n21199) );
NAND2_X1 MEM_stage_inst_dmem_U21093 ( .A1(MEM_stage_inst_dmem_n21197), .A2(MEM_stage_inst_dmem_n21196), .ZN(MEM_stage_inst_dmem_n8898) );
NAND2_X1 MEM_stage_inst_dmem_U21092 ( .A1(MEM_stage_inst_dmem_n17), .A2(MEM_stage_inst_dmem_n21211), .ZN(MEM_stage_inst_dmem_n21196) );
NAND2_X1 MEM_stage_inst_dmem_U21091 ( .A1(MEM_stage_inst_dmem_ram_3719), .A2(MEM_stage_inst_dmem_n21210), .ZN(MEM_stage_inst_dmem_n21197) );
NAND2_X1 MEM_stage_inst_dmem_U21090 ( .A1(MEM_stage_inst_dmem_n21195), .A2(MEM_stage_inst_dmem_n21194), .ZN(MEM_stage_inst_dmem_n8899) );
NAND2_X1 MEM_stage_inst_dmem_U21089 ( .A1(MEM_stage_inst_dmem_n21335), .A2(MEM_stage_inst_dmem_n21211), .ZN(MEM_stage_inst_dmem_n21194) );
NAND2_X1 MEM_stage_inst_dmem_U21088 ( .A1(MEM_stage_inst_dmem_ram_3720), .A2(MEM_stage_inst_dmem_n21210), .ZN(MEM_stage_inst_dmem_n21195) );
NAND2_X1 MEM_stage_inst_dmem_U21087 ( .A1(MEM_stage_inst_dmem_n21193), .A2(MEM_stage_inst_dmem_n21192), .ZN(MEM_stage_inst_dmem_n8900) );
NAND2_X1 MEM_stage_inst_dmem_U21086 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n21211), .ZN(MEM_stage_inst_dmem_n21192) );
NAND2_X1 MEM_stage_inst_dmem_U21085 ( .A1(MEM_stage_inst_dmem_ram_3721), .A2(MEM_stage_inst_dmem_n21210), .ZN(MEM_stage_inst_dmem_n21193) );
NAND2_X1 MEM_stage_inst_dmem_U21084 ( .A1(MEM_stage_inst_dmem_n21191), .A2(MEM_stage_inst_dmem_n21190), .ZN(MEM_stage_inst_dmem_n8901) );
NAND2_X1 MEM_stage_inst_dmem_U21083 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n21211), .ZN(MEM_stage_inst_dmem_n21190) );
NAND2_X1 MEM_stage_inst_dmem_U21082 ( .A1(MEM_stage_inst_dmem_ram_3722), .A2(MEM_stage_inst_dmem_n21210), .ZN(MEM_stage_inst_dmem_n21191) );
NAND2_X1 MEM_stage_inst_dmem_U21081 ( .A1(MEM_stage_inst_dmem_n21189), .A2(MEM_stage_inst_dmem_n21188), .ZN(MEM_stage_inst_dmem_n8902) );
NAND2_X1 MEM_stage_inst_dmem_U21080 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n21211), .ZN(MEM_stage_inst_dmem_n21188) );
NAND2_X1 MEM_stage_inst_dmem_U21079 ( .A1(MEM_stage_inst_dmem_ram_3723), .A2(MEM_stage_inst_dmem_n21210), .ZN(MEM_stage_inst_dmem_n21189) );
NAND2_X1 MEM_stage_inst_dmem_U21078 ( .A1(MEM_stage_inst_dmem_n21187), .A2(MEM_stage_inst_dmem_n21186), .ZN(MEM_stage_inst_dmem_n8903) );
NAND2_X1 MEM_stage_inst_dmem_U21077 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n21211), .ZN(MEM_stage_inst_dmem_n21186) );
NAND2_X1 MEM_stage_inst_dmem_U21076 ( .A1(MEM_stage_inst_dmem_ram_3724), .A2(MEM_stage_inst_dmem_n21210), .ZN(MEM_stage_inst_dmem_n21187) );
NAND2_X1 MEM_stage_inst_dmem_U21075 ( .A1(MEM_stage_inst_dmem_n21185), .A2(MEM_stage_inst_dmem_n21184), .ZN(MEM_stage_inst_dmem_n8904) );
NAND2_X1 MEM_stage_inst_dmem_U21074 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n21211), .ZN(MEM_stage_inst_dmem_n21184) );
NAND2_X1 MEM_stage_inst_dmem_U21073 ( .A1(MEM_stage_inst_dmem_ram_3725), .A2(MEM_stage_inst_dmem_n21210), .ZN(MEM_stage_inst_dmem_n21185) );
NAND2_X1 MEM_stage_inst_dmem_U21072 ( .A1(MEM_stage_inst_dmem_n21183), .A2(MEM_stage_inst_dmem_n21182), .ZN(MEM_stage_inst_dmem_n8905) );
NAND2_X1 MEM_stage_inst_dmem_U21071 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n21211), .ZN(MEM_stage_inst_dmem_n21182) );
NAND2_X1 MEM_stage_inst_dmem_U21070 ( .A1(MEM_stage_inst_dmem_ram_3726), .A2(MEM_stage_inst_dmem_n21210), .ZN(MEM_stage_inst_dmem_n21183) );
NAND2_X1 MEM_stage_inst_dmem_U21069 ( .A1(MEM_stage_inst_dmem_n21181), .A2(MEM_stage_inst_dmem_n21180), .ZN(MEM_stage_inst_dmem_n8906) );
NAND2_X1 MEM_stage_inst_dmem_U21068 ( .A1(MEM_stage_inst_dmem_n21320), .A2(MEM_stage_inst_dmem_n21211), .ZN(MEM_stage_inst_dmem_n21180) );
INV_X1 MEM_stage_inst_dmem_U21067 ( .A(MEM_stage_inst_dmem_n21210), .ZN(MEM_stage_inst_dmem_n21211) );
NAND2_X1 MEM_stage_inst_dmem_U21066 ( .A1(MEM_stage_inst_dmem_ram_3727), .A2(MEM_stage_inst_dmem_n21210), .ZN(MEM_stage_inst_dmem_n21181) );
NAND2_X1 MEM_stage_inst_dmem_U21065 ( .A1(MEM_stage_inst_dmem_n21179), .A2(MEM_stage_inst_dmem_n21464), .ZN(MEM_stage_inst_dmem_n21210) );
NAND2_X1 MEM_stage_inst_dmem_U21064 ( .A1(MEM_stage_inst_dmem_n21178), .A2(MEM_stage_inst_dmem_n21177), .ZN(MEM_stage_inst_dmem_n8907) );
NAND2_X1 MEM_stage_inst_dmem_U21063 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n21176), .ZN(MEM_stage_inst_dmem_n21177) );
NAND2_X1 MEM_stage_inst_dmem_U21062 ( .A1(MEM_stage_inst_dmem_ram_3728), .A2(MEM_stage_inst_dmem_n21175), .ZN(MEM_stage_inst_dmem_n21178) );
NAND2_X1 MEM_stage_inst_dmem_U21061 ( .A1(MEM_stage_inst_dmem_n21174), .A2(MEM_stage_inst_dmem_n21173), .ZN(MEM_stage_inst_dmem_n8908) );
NAND2_X1 MEM_stage_inst_dmem_U21060 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n21176), .ZN(MEM_stage_inst_dmem_n21173) );
NAND2_X1 MEM_stage_inst_dmem_U21059 ( .A1(MEM_stage_inst_dmem_ram_3729), .A2(MEM_stage_inst_dmem_n21175), .ZN(MEM_stage_inst_dmem_n21174) );
NAND2_X1 MEM_stage_inst_dmem_U21058 ( .A1(MEM_stage_inst_dmem_n21172), .A2(MEM_stage_inst_dmem_n21171), .ZN(MEM_stage_inst_dmem_n8909) );
NAND2_X1 MEM_stage_inst_dmem_U21057 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n21176), .ZN(MEM_stage_inst_dmem_n21171) );
NAND2_X1 MEM_stage_inst_dmem_U21056 ( .A1(MEM_stage_inst_dmem_ram_3730), .A2(MEM_stage_inst_dmem_n21175), .ZN(MEM_stage_inst_dmem_n21172) );
NAND2_X1 MEM_stage_inst_dmem_U21055 ( .A1(MEM_stage_inst_dmem_n21170), .A2(MEM_stage_inst_dmem_n21169), .ZN(MEM_stage_inst_dmem_n8910) );
NAND2_X1 MEM_stage_inst_dmem_U21054 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n21176), .ZN(MEM_stage_inst_dmem_n21169) );
NAND2_X1 MEM_stage_inst_dmem_U21053 ( .A1(MEM_stage_inst_dmem_ram_3731), .A2(MEM_stage_inst_dmem_n21175), .ZN(MEM_stage_inst_dmem_n21170) );
NAND2_X1 MEM_stage_inst_dmem_U21052 ( .A1(MEM_stage_inst_dmem_n21168), .A2(MEM_stage_inst_dmem_n21167), .ZN(MEM_stage_inst_dmem_n8911) );
NAND2_X1 MEM_stage_inst_dmem_U21051 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n21176), .ZN(MEM_stage_inst_dmem_n21167) );
NAND2_X1 MEM_stage_inst_dmem_U21050 ( .A1(MEM_stage_inst_dmem_ram_3732), .A2(MEM_stage_inst_dmem_n21175), .ZN(MEM_stage_inst_dmem_n21168) );
NAND2_X1 MEM_stage_inst_dmem_U21049 ( .A1(MEM_stage_inst_dmem_n21166), .A2(MEM_stage_inst_dmem_n21165), .ZN(MEM_stage_inst_dmem_n8912) );
NAND2_X1 MEM_stage_inst_dmem_U21048 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n21176), .ZN(MEM_stage_inst_dmem_n21165) );
NAND2_X1 MEM_stage_inst_dmem_U21047 ( .A1(MEM_stage_inst_dmem_ram_3733), .A2(MEM_stage_inst_dmem_n21175), .ZN(MEM_stage_inst_dmem_n21166) );
NAND2_X1 MEM_stage_inst_dmem_U21046 ( .A1(MEM_stage_inst_dmem_n21164), .A2(MEM_stage_inst_dmem_n21163), .ZN(MEM_stage_inst_dmem_n8913) );
NAND2_X1 MEM_stage_inst_dmem_U21045 ( .A1(MEM_stage_inst_dmem_n21340), .A2(MEM_stage_inst_dmem_n21176), .ZN(MEM_stage_inst_dmem_n21163) );
NAND2_X1 MEM_stage_inst_dmem_U21044 ( .A1(MEM_stage_inst_dmem_ram_3734), .A2(MEM_stage_inst_dmem_n21175), .ZN(MEM_stage_inst_dmem_n21164) );
NAND2_X1 MEM_stage_inst_dmem_U21043 ( .A1(MEM_stage_inst_dmem_n21162), .A2(MEM_stage_inst_dmem_n21161), .ZN(MEM_stage_inst_dmem_n8914) );
NAND2_X1 MEM_stage_inst_dmem_U21042 ( .A1(MEM_stage_inst_dmem_n18), .A2(MEM_stage_inst_dmem_n21176), .ZN(MEM_stage_inst_dmem_n21161) );
NAND2_X1 MEM_stage_inst_dmem_U21041 ( .A1(MEM_stage_inst_dmem_ram_3735), .A2(MEM_stage_inst_dmem_n21175), .ZN(MEM_stage_inst_dmem_n21162) );
NAND2_X1 MEM_stage_inst_dmem_U21040 ( .A1(MEM_stage_inst_dmem_n21160), .A2(MEM_stage_inst_dmem_n21159), .ZN(MEM_stage_inst_dmem_n8915) );
NAND2_X1 MEM_stage_inst_dmem_U21039 ( .A1(MEM_stage_inst_dmem_n21335), .A2(MEM_stage_inst_dmem_n21176), .ZN(MEM_stage_inst_dmem_n21159) );
NAND2_X1 MEM_stage_inst_dmem_U21038 ( .A1(MEM_stage_inst_dmem_ram_3736), .A2(MEM_stage_inst_dmem_n21175), .ZN(MEM_stage_inst_dmem_n21160) );
NAND2_X1 MEM_stage_inst_dmem_U21037 ( .A1(MEM_stage_inst_dmem_n21158), .A2(MEM_stage_inst_dmem_n21157), .ZN(MEM_stage_inst_dmem_n8916) );
NAND2_X1 MEM_stage_inst_dmem_U21036 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n21176), .ZN(MEM_stage_inst_dmem_n21157) );
NAND2_X1 MEM_stage_inst_dmem_U21035 ( .A1(MEM_stage_inst_dmem_ram_3737), .A2(MEM_stage_inst_dmem_n21175), .ZN(MEM_stage_inst_dmem_n21158) );
NAND2_X1 MEM_stage_inst_dmem_U21034 ( .A1(MEM_stage_inst_dmem_n21156), .A2(MEM_stage_inst_dmem_n21155), .ZN(MEM_stage_inst_dmem_n8917) );
NAND2_X1 MEM_stage_inst_dmem_U21033 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n21176), .ZN(MEM_stage_inst_dmem_n21155) );
NAND2_X1 MEM_stage_inst_dmem_U21032 ( .A1(MEM_stage_inst_dmem_ram_3738), .A2(MEM_stage_inst_dmem_n21175), .ZN(MEM_stage_inst_dmem_n21156) );
NAND2_X1 MEM_stage_inst_dmem_U21031 ( .A1(MEM_stage_inst_dmem_n21154), .A2(MEM_stage_inst_dmem_n21153), .ZN(MEM_stage_inst_dmem_n8918) );
NAND2_X1 MEM_stage_inst_dmem_U21030 ( .A1(MEM_stage_inst_dmem_n20904), .A2(MEM_stage_inst_dmem_n21176), .ZN(MEM_stage_inst_dmem_n21153) );
NAND2_X1 MEM_stage_inst_dmem_U21029 ( .A1(MEM_stage_inst_dmem_ram_3739), .A2(MEM_stage_inst_dmem_n21175), .ZN(MEM_stage_inst_dmem_n21154) );
NAND2_X1 MEM_stage_inst_dmem_U21028 ( .A1(MEM_stage_inst_dmem_n21152), .A2(MEM_stage_inst_dmem_n21151), .ZN(MEM_stage_inst_dmem_n8919) );
NAND2_X1 MEM_stage_inst_dmem_U21027 ( .A1(MEM_stage_inst_dmem_n21474), .A2(MEM_stage_inst_dmem_n21176), .ZN(MEM_stage_inst_dmem_n21151) );
NAND2_X1 MEM_stage_inst_dmem_U21026 ( .A1(MEM_stage_inst_dmem_ram_3740), .A2(MEM_stage_inst_dmem_n21175), .ZN(MEM_stage_inst_dmem_n21152) );
NAND2_X1 MEM_stage_inst_dmem_U21025 ( .A1(MEM_stage_inst_dmem_n21150), .A2(MEM_stage_inst_dmem_n21149), .ZN(MEM_stage_inst_dmem_n8920) );
NAND2_X1 MEM_stage_inst_dmem_U21024 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n21176), .ZN(MEM_stage_inst_dmem_n21149) );
NAND2_X1 MEM_stage_inst_dmem_U21023 ( .A1(MEM_stage_inst_dmem_ram_3741), .A2(MEM_stage_inst_dmem_n21175), .ZN(MEM_stage_inst_dmem_n21150) );
NAND2_X1 MEM_stage_inst_dmem_U21022 ( .A1(MEM_stage_inst_dmem_n21148), .A2(MEM_stage_inst_dmem_n21147), .ZN(MEM_stage_inst_dmem_n8921) );
NAND2_X1 MEM_stage_inst_dmem_U21021 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n21176), .ZN(MEM_stage_inst_dmem_n21147) );
NAND2_X1 MEM_stage_inst_dmem_U21020 ( .A1(MEM_stage_inst_dmem_ram_3742), .A2(MEM_stage_inst_dmem_n21175), .ZN(MEM_stage_inst_dmem_n21148) );
NAND2_X1 MEM_stage_inst_dmem_U21019 ( .A1(MEM_stage_inst_dmem_n21146), .A2(MEM_stage_inst_dmem_n21145), .ZN(MEM_stage_inst_dmem_n8922) );
NAND2_X1 MEM_stage_inst_dmem_U21018 ( .A1(MEM_stage_inst_dmem_n21320), .A2(MEM_stage_inst_dmem_n21176), .ZN(MEM_stage_inst_dmem_n21145) );
INV_X1 MEM_stage_inst_dmem_U21017 ( .A(MEM_stage_inst_dmem_n21175), .ZN(MEM_stage_inst_dmem_n21176) );
NAND2_X1 MEM_stage_inst_dmem_U21016 ( .A1(MEM_stage_inst_dmem_ram_3743), .A2(MEM_stage_inst_dmem_n21175), .ZN(MEM_stage_inst_dmem_n21146) );
NAND2_X1 MEM_stage_inst_dmem_U21015 ( .A1(MEM_stage_inst_dmem_n21144), .A2(MEM_stage_inst_dmem_n21464), .ZN(MEM_stage_inst_dmem_n21175) );
NAND2_X1 MEM_stage_inst_dmem_U21014 ( .A1(MEM_stage_inst_dmem_n21143), .A2(MEM_stage_inst_dmem_n21142), .ZN(MEM_stage_inst_dmem_n8923) );
NAND2_X1 MEM_stage_inst_dmem_U21013 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n21141), .ZN(MEM_stage_inst_dmem_n21142) );
NAND2_X1 MEM_stage_inst_dmem_U21012 ( .A1(MEM_stage_inst_dmem_ram_3744), .A2(MEM_stage_inst_dmem_n21140), .ZN(MEM_stage_inst_dmem_n21143) );
NAND2_X1 MEM_stage_inst_dmem_U21011 ( .A1(MEM_stage_inst_dmem_n21139), .A2(MEM_stage_inst_dmem_n21138), .ZN(MEM_stage_inst_dmem_n8924) );
NAND2_X1 MEM_stage_inst_dmem_U21010 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n21141), .ZN(MEM_stage_inst_dmem_n21138) );
NAND2_X1 MEM_stage_inst_dmem_U21009 ( .A1(MEM_stage_inst_dmem_ram_3745), .A2(MEM_stage_inst_dmem_n21140), .ZN(MEM_stage_inst_dmem_n21139) );
NAND2_X1 MEM_stage_inst_dmem_U21008 ( .A1(MEM_stage_inst_dmem_n21137), .A2(MEM_stage_inst_dmem_n21136), .ZN(MEM_stage_inst_dmem_n8925) );
NAND2_X1 MEM_stage_inst_dmem_U21007 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n21141), .ZN(MEM_stage_inst_dmem_n21136) );
NAND2_X1 MEM_stage_inst_dmem_U21006 ( .A1(MEM_stage_inst_dmem_ram_3746), .A2(MEM_stage_inst_dmem_n21140), .ZN(MEM_stage_inst_dmem_n21137) );
NAND2_X1 MEM_stage_inst_dmem_U21005 ( .A1(MEM_stage_inst_dmem_n21135), .A2(MEM_stage_inst_dmem_n21134), .ZN(MEM_stage_inst_dmem_n8926) );
NAND2_X1 MEM_stage_inst_dmem_U21004 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n21141), .ZN(MEM_stage_inst_dmem_n21134) );
NAND2_X1 MEM_stage_inst_dmem_U21003 ( .A1(MEM_stage_inst_dmem_ram_3747), .A2(MEM_stage_inst_dmem_n21140), .ZN(MEM_stage_inst_dmem_n21135) );
NAND2_X1 MEM_stage_inst_dmem_U21002 ( .A1(MEM_stage_inst_dmem_n21133), .A2(MEM_stage_inst_dmem_n21132), .ZN(MEM_stage_inst_dmem_n8927) );
NAND2_X1 MEM_stage_inst_dmem_U21001 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n21141), .ZN(MEM_stage_inst_dmem_n21132) );
NAND2_X1 MEM_stage_inst_dmem_U21000 ( .A1(MEM_stage_inst_dmem_ram_3748), .A2(MEM_stage_inst_dmem_n21140), .ZN(MEM_stage_inst_dmem_n21133) );
NAND2_X1 MEM_stage_inst_dmem_U20999 ( .A1(MEM_stage_inst_dmem_n21131), .A2(MEM_stage_inst_dmem_n21130), .ZN(MEM_stage_inst_dmem_n8928) );
NAND2_X1 MEM_stage_inst_dmem_U20998 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n21141), .ZN(MEM_stage_inst_dmem_n21130) );
NAND2_X1 MEM_stage_inst_dmem_U20997 ( .A1(MEM_stage_inst_dmem_ram_3749), .A2(MEM_stage_inst_dmem_n21140), .ZN(MEM_stage_inst_dmem_n21131) );
NAND2_X1 MEM_stage_inst_dmem_U20996 ( .A1(MEM_stage_inst_dmem_n21129), .A2(MEM_stage_inst_dmem_n21128), .ZN(MEM_stage_inst_dmem_n8929) );
NAND2_X1 MEM_stage_inst_dmem_U20995 ( .A1(MEM_stage_inst_dmem_n21340), .A2(MEM_stage_inst_dmem_n21141), .ZN(MEM_stage_inst_dmem_n21128) );
NAND2_X1 MEM_stage_inst_dmem_U20994 ( .A1(MEM_stage_inst_dmem_ram_3750), .A2(MEM_stage_inst_dmem_n21140), .ZN(MEM_stage_inst_dmem_n21129) );
NAND2_X1 MEM_stage_inst_dmem_U20993 ( .A1(MEM_stage_inst_dmem_n21127), .A2(MEM_stage_inst_dmem_n21126), .ZN(MEM_stage_inst_dmem_n8930) );
NAND2_X1 MEM_stage_inst_dmem_U20992 ( .A1(MEM_stage_inst_dmem_n17), .A2(MEM_stage_inst_dmem_n21141), .ZN(MEM_stage_inst_dmem_n21126) );
NAND2_X1 MEM_stage_inst_dmem_U20991 ( .A1(MEM_stage_inst_dmem_ram_3751), .A2(MEM_stage_inst_dmem_n21140), .ZN(MEM_stage_inst_dmem_n21127) );
NAND2_X1 MEM_stage_inst_dmem_U20990 ( .A1(MEM_stage_inst_dmem_n21125), .A2(MEM_stage_inst_dmem_n21124), .ZN(MEM_stage_inst_dmem_n8931) );
NAND2_X1 MEM_stage_inst_dmem_U20989 ( .A1(MEM_stage_inst_dmem_n21335), .A2(MEM_stage_inst_dmem_n21141), .ZN(MEM_stage_inst_dmem_n21124) );
NAND2_X1 MEM_stage_inst_dmem_U20988 ( .A1(MEM_stage_inst_dmem_ram_3752), .A2(MEM_stage_inst_dmem_n21140), .ZN(MEM_stage_inst_dmem_n21125) );
NAND2_X1 MEM_stage_inst_dmem_U20987 ( .A1(MEM_stage_inst_dmem_n21123), .A2(MEM_stage_inst_dmem_n21122), .ZN(MEM_stage_inst_dmem_n8932) );
NAND2_X1 MEM_stage_inst_dmem_U20986 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n21141), .ZN(MEM_stage_inst_dmem_n21122) );
NAND2_X1 MEM_stage_inst_dmem_U20985 ( .A1(MEM_stage_inst_dmem_ram_3753), .A2(MEM_stage_inst_dmem_n21140), .ZN(MEM_stage_inst_dmem_n21123) );
NAND2_X1 MEM_stage_inst_dmem_U20984 ( .A1(MEM_stage_inst_dmem_n21121), .A2(MEM_stage_inst_dmem_n21120), .ZN(MEM_stage_inst_dmem_n8933) );
NAND2_X1 MEM_stage_inst_dmem_U20983 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n21141), .ZN(MEM_stage_inst_dmem_n21120) );
NAND2_X1 MEM_stage_inst_dmem_U20982 ( .A1(MEM_stage_inst_dmem_ram_3754), .A2(MEM_stage_inst_dmem_n21140), .ZN(MEM_stage_inst_dmem_n21121) );
NAND2_X1 MEM_stage_inst_dmem_U20981 ( .A1(MEM_stage_inst_dmem_n21119), .A2(MEM_stage_inst_dmem_n21118), .ZN(MEM_stage_inst_dmem_n8934) );
NAND2_X1 MEM_stage_inst_dmem_U20980 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n21141), .ZN(MEM_stage_inst_dmem_n21118) );
NAND2_X1 MEM_stage_inst_dmem_U20979 ( .A1(MEM_stage_inst_dmem_ram_3755), .A2(MEM_stage_inst_dmem_n21140), .ZN(MEM_stage_inst_dmem_n21119) );
NAND2_X1 MEM_stage_inst_dmem_U20978 ( .A1(MEM_stage_inst_dmem_n21117), .A2(MEM_stage_inst_dmem_n21116), .ZN(MEM_stage_inst_dmem_n8935) );
NAND2_X1 MEM_stage_inst_dmem_U20977 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n21141), .ZN(MEM_stage_inst_dmem_n21116) );
NAND2_X1 MEM_stage_inst_dmem_U20976 ( .A1(MEM_stage_inst_dmem_ram_3756), .A2(MEM_stage_inst_dmem_n21140), .ZN(MEM_stage_inst_dmem_n21117) );
NAND2_X1 MEM_stage_inst_dmem_U20975 ( .A1(MEM_stage_inst_dmem_n21115), .A2(MEM_stage_inst_dmem_n21114), .ZN(MEM_stage_inst_dmem_n8936) );
NAND2_X1 MEM_stage_inst_dmem_U20974 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n21141), .ZN(MEM_stage_inst_dmem_n21114) );
NAND2_X1 MEM_stage_inst_dmem_U20973 ( .A1(MEM_stage_inst_dmem_ram_3757), .A2(MEM_stage_inst_dmem_n21140), .ZN(MEM_stage_inst_dmem_n21115) );
NAND2_X1 MEM_stage_inst_dmem_U20972 ( .A1(MEM_stage_inst_dmem_n21113), .A2(MEM_stage_inst_dmem_n21112), .ZN(MEM_stage_inst_dmem_n8937) );
NAND2_X1 MEM_stage_inst_dmem_U20971 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n21141), .ZN(MEM_stage_inst_dmem_n21112) );
NAND2_X1 MEM_stage_inst_dmem_U20970 ( .A1(MEM_stage_inst_dmem_ram_3758), .A2(MEM_stage_inst_dmem_n21140), .ZN(MEM_stage_inst_dmem_n21113) );
NAND2_X1 MEM_stage_inst_dmem_U20969 ( .A1(MEM_stage_inst_dmem_n21111), .A2(MEM_stage_inst_dmem_n21110), .ZN(MEM_stage_inst_dmem_n8938) );
NAND2_X1 MEM_stage_inst_dmem_U20968 ( .A1(MEM_stage_inst_dmem_n21320), .A2(MEM_stage_inst_dmem_n21141), .ZN(MEM_stage_inst_dmem_n21110) );
NAND2_X1 MEM_stage_inst_dmem_U20967 ( .A1(MEM_stage_inst_dmem_ram_3759), .A2(MEM_stage_inst_dmem_n21140), .ZN(MEM_stage_inst_dmem_n21111) );
NAND2_X1 MEM_stage_inst_dmem_U20966 ( .A1(MEM_stage_inst_dmem_n21109), .A2(MEM_stage_inst_dmem_n21464), .ZN(MEM_stage_inst_dmem_n21140) );
NAND2_X1 MEM_stage_inst_dmem_U20965 ( .A1(MEM_stage_inst_dmem_n21108), .A2(MEM_stage_inst_dmem_n21107), .ZN(MEM_stage_inst_dmem_n8939) );
NAND2_X1 MEM_stage_inst_dmem_U20964 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n21106), .ZN(MEM_stage_inst_dmem_n21107) );
NAND2_X1 MEM_stage_inst_dmem_U20963 ( .A1(MEM_stage_inst_dmem_ram_3760), .A2(MEM_stage_inst_dmem_n21105), .ZN(MEM_stage_inst_dmem_n21108) );
NAND2_X1 MEM_stage_inst_dmem_U20962 ( .A1(MEM_stage_inst_dmem_n21104), .A2(MEM_stage_inst_dmem_n21103), .ZN(MEM_stage_inst_dmem_n8940) );
NAND2_X1 MEM_stage_inst_dmem_U20961 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n21106), .ZN(MEM_stage_inst_dmem_n21103) );
NAND2_X1 MEM_stage_inst_dmem_U20960 ( .A1(MEM_stage_inst_dmem_ram_3761), .A2(MEM_stage_inst_dmem_n21105), .ZN(MEM_stage_inst_dmem_n21104) );
NAND2_X1 MEM_stage_inst_dmem_U20959 ( .A1(MEM_stage_inst_dmem_n21102), .A2(MEM_stage_inst_dmem_n21101), .ZN(MEM_stage_inst_dmem_n8941) );
NAND2_X1 MEM_stage_inst_dmem_U20958 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n21106), .ZN(MEM_stage_inst_dmem_n21101) );
NAND2_X1 MEM_stage_inst_dmem_U20957 ( .A1(MEM_stage_inst_dmem_ram_3762), .A2(MEM_stage_inst_dmem_n21105), .ZN(MEM_stage_inst_dmem_n21102) );
NAND2_X1 MEM_stage_inst_dmem_U20956 ( .A1(MEM_stage_inst_dmem_n21100), .A2(MEM_stage_inst_dmem_n21099), .ZN(MEM_stage_inst_dmem_n8942) );
NAND2_X1 MEM_stage_inst_dmem_U20955 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n21106), .ZN(MEM_stage_inst_dmem_n21099) );
NAND2_X1 MEM_stage_inst_dmem_U20954 ( .A1(MEM_stage_inst_dmem_ram_3763), .A2(MEM_stage_inst_dmem_n21105), .ZN(MEM_stage_inst_dmem_n21100) );
NAND2_X1 MEM_stage_inst_dmem_U20953 ( .A1(MEM_stage_inst_dmem_n21098), .A2(MEM_stage_inst_dmem_n21097), .ZN(MEM_stage_inst_dmem_n8943) );
NAND2_X1 MEM_stage_inst_dmem_U20952 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n21106), .ZN(MEM_stage_inst_dmem_n21097) );
NAND2_X1 MEM_stage_inst_dmem_U20951 ( .A1(MEM_stage_inst_dmem_ram_3764), .A2(MEM_stage_inst_dmem_n21105), .ZN(MEM_stage_inst_dmem_n21098) );
NAND2_X1 MEM_stage_inst_dmem_U20950 ( .A1(MEM_stage_inst_dmem_n21096), .A2(MEM_stage_inst_dmem_n21095), .ZN(MEM_stage_inst_dmem_n8944) );
NAND2_X1 MEM_stage_inst_dmem_U20949 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n21106), .ZN(MEM_stage_inst_dmem_n21095) );
NAND2_X1 MEM_stage_inst_dmem_U20948 ( .A1(MEM_stage_inst_dmem_ram_3765), .A2(MEM_stage_inst_dmem_n21105), .ZN(MEM_stage_inst_dmem_n21096) );
NAND2_X1 MEM_stage_inst_dmem_U20947 ( .A1(MEM_stage_inst_dmem_n21094), .A2(MEM_stage_inst_dmem_n21093), .ZN(MEM_stage_inst_dmem_n8945) );
NAND2_X1 MEM_stage_inst_dmem_U20946 ( .A1(MEM_stage_inst_dmem_n21340), .A2(MEM_stage_inst_dmem_n21106), .ZN(MEM_stage_inst_dmem_n21093) );
NAND2_X1 MEM_stage_inst_dmem_U20945 ( .A1(MEM_stage_inst_dmem_ram_3766), .A2(MEM_stage_inst_dmem_n21105), .ZN(MEM_stage_inst_dmem_n21094) );
NAND2_X1 MEM_stage_inst_dmem_U20944 ( .A1(MEM_stage_inst_dmem_n21092), .A2(MEM_stage_inst_dmem_n21091), .ZN(MEM_stage_inst_dmem_n8946) );
NAND2_X1 MEM_stage_inst_dmem_U20943 ( .A1(MEM_stage_inst_dmem_n18), .A2(MEM_stage_inst_dmem_n21106), .ZN(MEM_stage_inst_dmem_n21091) );
NAND2_X1 MEM_stage_inst_dmem_U20942 ( .A1(MEM_stage_inst_dmem_ram_3767), .A2(MEM_stage_inst_dmem_n21105), .ZN(MEM_stage_inst_dmem_n21092) );
NAND2_X1 MEM_stage_inst_dmem_U20941 ( .A1(MEM_stage_inst_dmem_n21090), .A2(MEM_stage_inst_dmem_n21089), .ZN(MEM_stage_inst_dmem_n8947) );
NAND2_X1 MEM_stage_inst_dmem_U20940 ( .A1(MEM_stage_inst_dmem_n21335), .A2(MEM_stage_inst_dmem_n21106), .ZN(MEM_stage_inst_dmem_n21089) );
NAND2_X1 MEM_stage_inst_dmem_U20939 ( .A1(MEM_stage_inst_dmem_ram_3768), .A2(MEM_stage_inst_dmem_n21105), .ZN(MEM_stage_inst_dmem_n21090) );
NAND2_X1 MEM_stage_inst_dmem_U20938 ( .A1(MEM_stage_inst_dmem_n21088), .A2(MEM_stage_inst_dmem_n21087), .ZN(MEM_stage_inst_dmem_n8948) );
NAND2_X1 MEM_stage_inst_dmem_U20937 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n21106), .ZN(MEM_stage_inst_dmem_n21087) );
NAND2_X1 MEM_stage_inst_dmem_U20936 ( .A1(MEM_stage_inst_dmem_ram_3769), .A2(MEM_stage_inst_dmem_n21105), .ZN(MEM_stage_inst_dmem_n21088) );
NAND2_X1 MEM_stage_inst_dmem_U20935 ( .A1(MEM_stage_inst_dmem_n21086), .A2(MEM_stage_inst_dmem_n21085), .ZN(MEM_stage_inst_dmem_n8949) );
NAND2_X1 MEM_stage_inst_dmem_U20934 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n21106), .ZN(MEM_stage_inst_dmem_n21085) );
NAND2_X1 MEM_stage_inst_dmem_U20933 ( .A1(MEM_stage_inst_dmem_ram_3770), .A2(MEM_stage_inst_dmem_n21105), .ZN(MEM_stage_inst_dmem_n21086) );
NAND2_X1 MEM_stage_inst_dmem_U20932 ( .A1(MEM_stage_inst_dmem_n21084), .A2(MEM_stage_inst_dmem_n21083), .ZN(MEM_stage_inst_dmem_n8950) );
NAND2_X1 MEM_stage_inst_dmem_U20931 ( .A1(MEM_stage_inst_dmem_n14705), .A2(MEM_stage_inst_dmem_n21106), .ZN(MEM_stage_inst_dmem_n21083) );
NAND2_X1 MEM_stage_inst_dmem_U20930 ( .A1(MEM_stage_inst_dmem_ram_3771), .A2(MEM_stage_inst_dmem_n21105), .ZN(MEM_stage_inst_dmem_n21084) );
NAND2_X1 MEM_stage_inst_dmem_U20929 ( .A1(MEM_stage_inst_dmem_n21082), .A2(MEM_stage_inst_dmem_n21081), .ZN(MEM_stage_inst_dmem_n8951) );
NAND2_X1 MEM_stage_inst_dmem_U20928 ( .A1(MEM_stage_inst_dmem_n14702), .A2(MEM_stage_inst_dmem_n21106), .ZN(MEM_stage_inst_dmem_n21081) );
NAND2_X1 MEM_stage_inst_dmem_U20927 ( .A1(MEM_stage_inst_dmem_ram_3772), .A2(MEM_stage_inst_dmem_n21105), .ZN(MEM_stage_inst_dmem_n21082) );
NAND2_X1 MEM_stage_inst_dmem_U20926 ( .A1(MEM_stage_inst_dmem_n21080), .A2(MEM_stage_inst_dmem_n21079), .ZN(MEM_stage_inst_dmem_n8952) );
NAND2_X1 MEM_stage_inst_dmem_U20925 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n21106), .ZN(MEM_stage_inst_dmem_n21079) );
NAND2_X1 MEM_stage_inst_dmem_U20924 ( .A1(MEM_stage_inst_dmem_ram_3773), .A2(MEM_stage_inst_dmem_n21105), .ZN(MEM_stage_inst_dmem_n21080) );
NAND2_X1 MEM_stage_inst_dmem_U20923 ( .A1(MEM_stage_inst_dmem_n21078), .A2(MEM_stage_inst_dmem_n21077), .ZN(MEM_stage_inst_dmem_n8953) );
NAND2_X1 MEM_stage_inst_dmem_U20922 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n21106), .ZN(MEM_stage_inst_dmem_n21077) );
NAND2_X1 MEM_stage_inst_dmem_U20921 ( .A1(MEM_stage_inst_dmem_ram_3774), .A2(MEM_stage_inst_dmem_n21105), .ZN(MEM_stage_inst_dmem_n21078) );
NAND2_X1 MEM_stage_inst_dmem_U20920 ( .A1(MEM_stage_inst_dmem_n21076), .A2(MEM_stage_inst_dmem_n21075), .ZN(MEM_stage_inst_dmem_n8954) );
NAND2_X1 MEM_stage_inst_dmem_U20919 ( .A1(MEM_stage_inst_dmem_n21320), .A2(MEM_stage_inst_dmem_n21106), .ZN(MEM_stage_inst_dmem_n21075) );
INV_X1 MEM_stage_inst_dmem_U20918 ( .A(MEM_stage_inst_dmem_n21105), .ZN(MEM_stage_inst_dmem_n21106) );
NAND2_X1 MEM_stage_inst_dmem_U20917 ( .A1(MEM_stage_inst_dmem_ram_3775), .A2(MEM_stage_inst_dmem_n21105), .ZN(MEM_stage_inst_dmem_n21076) );
NAND2_X1 MEM_stage_inst_dmem_U20916 ( .A1(MEM_stage_inst_dmem_n21074), .A2(MEM_stage_inst_dmem_n21464), .ZN(MEM_stage_inst_dmem_n21105) );
NAND2_X1 MEM_stage_inst_dmem_U20915 ( .A1(MEM_stage_inst_dmem_n21073), .A2(MEM_stage_inst_dmem_n21072), .ZN(MEM_stage_inst_dmem_n8955) );
NAND2_X1 MEM_stage_inst_dmem_U20914 ( .A1(MEM_stage_inst_dmem_n15145), .A2(MEM_stage_inst_dmem_n21071), .ZN(MEM_stage_inst_dmem_n21072) );
NAND2_X1 MEM_stage_inst_dmem_U20913 ( .A1(MEM_stage_inst_dmem_ram_3776), .A2(MEM_stage_inst_dmem_n21070), .ZN(MEM_stage_inst_dmem_n21073) );
NAND2_X1 MEM_stage_inst_dmem_U20912 ( .A1(MEM_stage_inst_dmem_n21069), .A2(MEM_stage_inst_dmem_n21068), .ZN(MEM_stage_inst_dmem_n8956) );
NAND2_X1 MEM_stage_inst_dmem_U20911 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n21071), .ZN(MEM_stage_inst_dmem_n21068) );
NAND2_X1 MEM_stage_inst_dmem_U20910 ( .A1(MEM_stage_inst_dmem_ram_3777), .A2(MEM_stage_inst_dmem_n21070), .ZN(MEM_stage_inst_dmem_n21069) );
NAND2_X1 MEM_stage_inst_dmem_U20909 ( .A1(MEM_stage_inst_dmem_n21067), .A2(MEM_stage_inst_dmem_n21066), .ZN(MEM_stage_inst_dmem_n8957) );
NAND2_X1 MEM_stage_inst_dmem_U20908 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n21071), .ZN(MEM_stage_inst_dmem_n21066) );
NAND2_X1 MEM_stage_inst_dmem_U20907 ( .A1(MEM_stage_inst_dmem_ram_3778), .A2(MEM_stage_inst_dmem_n21070), .ZN(MEM_stage_inst_dmem_n21067) );
NAND2_X1 MEM_stage_inst_dmem_U20906 ( .A1(MEM_stage_inst_dmem_n21065), .A2(MEM_stage_inst_dmem_n21064), .ZN(MEM_stage_inst_dmem_n8958) );
NAND2_X1 MEM_stage_inst_dmem_U20905 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n21071), .ZN(MEM_stage_inst_dmem_n21064) );
NAND2_X1 MEM_stage_inst_dmem_U20904 ( .A1(MEM_stage_inst_dmem_ram_3779), .A2(MEM_stage_inst_dmem_n21070), .ZN(MEM_stage_inst_dmem_n21065) );
NAND2_X1 MEM_stage_inst_dmem_U20903 ( .A1(MEM_stage_inst_dmem_n21063), .A2(MEM_stage_inst_dmem_n21062), .ZN(MEM_stage_inst_dmem_n8959) );
NAND2_X1 MEM_stage_inst_dmem_U20902 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n21071), .ZN(MEM_stage_inst_dmem_n21062) );
NAND2_X1 MEM_stage_inst_dmem_U20901 ( .A1(MEM_stage_inst_dmem_ram_3780), .A2(MEM_stage_inst_dmem_n21070), .ZN(MEM_stage_inst_dmem_n21063) );
NAND2_X1 MEM_stage_inst_dmem_U20900 ( .A1(MEM_stage_inst_dmem_n21061), .A2(MEM_stage_inst_dmem_n21060), .ZN(MEM_stage_inst_dmem_n8960) );
NAND2_X1 MEM_stage_inst_dmem_U20899 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n21071), .ZN(MEM_stage_inst_dmem_n21060) );
NAND2_X1 MEM_stage_inst_dmem_U20898 ( .A1(MEM_stage_inst_dmem_ram_3781), .A2(MEM_stage_inst_dmem_n21070), .ZN(MEM_stage_inst_dmem_n21061) );
NAND2_X1 MEM_stage_inst_dmem_U20897 ( .A1(MEM_stage_inst_dmem_n21059), .A2(MEM_stage_inst_dmem_n21058), .ZN(MEM_stage_inst_dmem_n8961) );
NAND2_X1 MEM_stage_inst_dmem_U20896 ( .A1(MEM_stage_inst_dmem_n21340), .A2(MEM_stage_inst_dmem_n21071), .ZN(MEM_stage_inst_dmem_n21058) );
NAND2_X1 MEM_stage_inst_dmem_U20895 ( .A1(MEM_stage_inst_dmem_ram_3782), .A2(MEM_stage_inst_dmem_n21070), .ZN(MEM_stage_inst_dmem_n21059) );
NAND2_X1 MEM_stage_inst_dmem_U20894 ( .A1(MEM_stage_inst_dmem_n21057), .A2(MEM_stage_inst_dmem_n21056), .ZN(MEM_stage_inst_dmem_n8962) );
NAND2_X1 MEM_stage_inst_dmem_U20893 ( .A1(MEM_stage_inst_dmem_n17), .A2(MEM_stage_inst_dmem_n21071), .ZN(MEM_stage_inst_dmem_n21056) );
NAND2_X1 MEM_stage_inst_dmem_U20892 ( .A1(MEM_stage_inst_dmem_ram_3783), .A2(MEM_stage_inst_dmem_n21070), .ZN(MEM_stage_inst_dmem_n21057) );
NAND2_X1 MEM_stage_inst_dmem_U20891 ( .A1(MEM_stage_inst_dmem_n21055), .A2(MEM_stage_inst_dmem_n21054), .ZN(MEM_stage_inst_dmem_n8963) );
NAND2_X1 MEM_stage_inst_dmem_U20890 ( .A1(MEM_stage_inst_dmem_n21335), .A2(MEM_stage_inst_dmem_n21071), .ZN(MEM_stage_inst_dmem_n21054) );
NAND2_X1 MEM_stage_inst_dmem_U20889 ( .A1(MEM_stage_inst_dmem_ram_3784), .A2(MEM_stage_inst_dmem_n21070), .ZN(MEM_stage_inst_dmem_n21055) );
NAND2_X1 MEM_stage_inst_dmem_U20888 ( .A1(MEM_stage_inst_dmem_n21053), .A2(MEM_stage_inst_dmem_n21052), .ZN(MEM_stage_inst_dmem_n8964) );
NAND2_X1 MEM_stage_inst_dmem_U20887 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n21071), .ZN(MEM_stage_inst_dmem_n21052) );
NAND2_X1 MEM_stage_inst_dmem_U20886 ( .A1(MEM_stage_inst_dmem_ram_3785), .A2(MEM_stage_inst_dmem_n21070), .ZN(MEM_stage_inst_dmem_n21053) );
NAND2_X1 MEM_stage_inst_dmem_U20885 ( .A1(MEM_stage_inst_dmem_n21051), .A2(MEM_stage_inst_dmem_n21050), .ZN(MEM_stage_inst_dmem_n8965) );
NAND2_X1 MEM_stage_inst_dmem_U20884 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n21071), .ZN(MEM_stage_inst_dmem_n21050) );
NAND2_X1 MEM_stage_inst_dmem_U20883 ( .A1(MEM_stage_inst_dmem_ram_3786), .A2(MEM_stage_inst_dmem_n21070), .ZN(MEM_stage_inst_dmem_n21051) );
NAND2_X1 MEM_stage_inst_dmem_U20882 ( .A1(MEM_stage_inst_dmem_n21049), .A2(MEM_stage_inst_dmem_n21048), .ZN(MEM_stage_inst_dmem_n8966) );
NAND2_X1 MEM_stage_inst_dmem_U20881 ( .A1(MEM_stage_inst_dmem_n13044), .A2(MEM_stage_inst_dmem_n21071), .ZN(MEM_stage_inst_dmem_n21048) );
NAND2_X1 MEM_stage_inst_dmem_U20880 ( .A1(MEM_stage_inst_dmem_ram_3787), .A2(MEM_stage_inst_dmem_n21070), .ZN(MEM_stage_inst_dmem_n21049) );
NAND2_X1 MEM_stage_inst_dmem_U20879 ( .A1(MEM_stage_inst_dmem_n21047), .A2(MEM_stage_inst_dmem_n21046), .ZN(MEM_stage_inst_dmem_n8967) );
NAND2_X1 MEM_stage_inst_dmem_U20878 ( .A1(MEM_stage_inst_dmem_n13041), .A2(MEM_stage_inst_dmem_n21071), .ZN(MEM_stage_inst_dmem_n21046) );
NAND2_X1 MEM_stage_inst_dmem_U20877 ( .A1(MEM_stage_inst_dmem_ram_3788), .A2(MEM_stage_inst_dmem_n21070), .ZN(MEM_stage_inst_dmem_n21047) );
NAND2_X1 MEM_stage_inst_dmem_U20876 ( .A1(MEM_stage_inst_dmem_n21045), .A2(MEM_stage_inst_dmem_n21044), .ZN(MEM_stage_inst_dmem_n8968) );
NAND2_X1 MEM_stage_inst_dmem_U20875 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n21071), .ZN(MEM_stage_inst_dmem_n21044) );
NAND2_X1 MEM_stage_inst_dmem_U20874 ( .A1(MEM_stage_inst_dmem_ram_3789), .A2(MEM_stage_inst_dmem_n21070), .ZN(MEM_stage_inst_dmem_n21045) );
NAND2_X1 MEM_stage_inst_dmem_U20873 ( .A1(MEM_stage_inst_dmem_n21043), .A2(MEM_stage_inst_dmem_n21042), .ZN(MEM_stage_inst_dmem_n8969) );
NAND2_X1 MEM_stage_inst_dmem_U20872 ( .A1(MEM_stage_inst_dmem_n15113), .A2(MEM_stage_inst_dmem_n21071), .ZN(MEM_stage_inst_dmem_n21042) );
NAND2_X1 MEM_stage_inst_dmem_U20871 ( .A1(MEM_stage_inst_dmem_ram_3790), .A2(MEM_stage_inst_dmem_n21070), .ZN(MEM_stage_inst_dmem_n21043) );
NAND2_X1 MEM_stage_inst_dmem_U20870 ( .A1(MEM_stage_inst_dmem_n21041), .A2(MEM_stage_inst_dmem_n21040), .ZN(MEM_stage_inst_dmem_n8970) );
NAND2_X1 MEM_stage_inst_dmem_U20869 ( .A1(MEM_stage_inst_dmem_n21320), .A2(MEM_stage_inst_dmem_n21071), .ZN(MEM_stage_inst_dmem_n21040) );
INV_X1 MEM_stage_inst_dmem_U20868 ( .A(MEM_stage_inst_dmem_n21070), .ZN(MEM_stage_inst_dmem_n21071) );
NAND2_X1 MEM_stage_inst_dmem_U20867 ( .A1(MEM_stage_inst_dmem_ram_3791), .A2(MEM_stage_inst_dmem_n21070), .ZN(MEM_stage_inst_dmem_n21041) );
NAND2_X1 MEM_stage_inst_dmem_U20866 ( .A1(MEM_stage_inst_dmem_n21039), .A2(MEM_stage_inst_dmem_n21464), .ZN(MEM_stage_inst_dmem_n21070) );
NAND2_X1 MEM_stage_inst_dmem_U20865 ( .A1(MEM_stage_inst_dmem_n21038), .A2(MEM_stage_inst_dmem_n21037), .ZN(MEM_stage_inst_dmem_n8971) );
NAND2_X1 MEM_stage_inst_dmem_U20864 ( .A1(MEM_stage_inst_dmem_n19275), .A2(MEM_stage_inst_dmem_n21036), .ZN(MEM_stage_inst_dmem_n21037) );
NAND2_X1 MEM_stage_inst_dmem_U20863 ( .A1(MEM_stage_inst_dmem_ram_3792), .A2(MEM_stage_inst_dmem_n21035), .ZN(MEM_stage_inst_dmem_n21038) );
NAND2_X1 MEM_stage_inst_dmem_U20862 ( .A1(MEM_stage_inst_dmem_n21034), .A2(MEM_stage_inst_dmem_n21033), .ZN(MEM_stage_inst_dmem_n8972) );
NAND2_X1 MEM_stage_inst_dmem_U20861 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n21036), .ZN(MEM_stage_inst_dmem_n21033) );
NAND2_X1 MEM_stage_inst_dmem_U20860 ( .A1(MEM_stage_inst_dmem_ram_3793), .A2(MEM_stage_inst_dmem_n21035), .ZN(MEM_stage_inst_dmem_n21034) );
NAND2_X1 MEM_stage_inst_dmem_U20859 ( .A1(MEM_stage_inst_dmem_n21032), .A2(MEM_stage_inst_dmem_n21031), .ZN(MEM_stage_inst_dmem_n8973) );
NAND2_X1 MEM_stage_inst_dmem_U20858 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n21036), .ZN(MEM_stage_inst_dmem_n21031) );
NAND2_X1 MEM_stage_inst_dmem_U20857 ( .A1(MEM_stage_inst_dmem_ram_3794), .A2(MEM_stage_inst_dmem_n21035), .ZN(MEM_stage_inst_dmem_n21032) );
NAND2_X1 MEM_stage_inst_dmem_U20856 ( .A1(MEM_stage_inst_dmem_n21030), .A2(MEM_stage_inst_dmem_n21029), .ZN(MEM_stage_inst_dmem_n8974) );
NAND2_X1 MEM_stage_inst_dmem_U20855 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n21036), .ZN(MEM_stage_inst_dmem_n21029) );
NAND2_X1 MEM_stage_inst_dmem_U20854 ( .A1(MEM_stage_inst_dmem_ram_3795), .A2(MEM_stage_inst_dmem_n21035), .ZN(MEM_stage_inst_dmem_n21030) );
NAND2_X1 MEM_stage_inst_dmem_U20853 ( .A1(MEM_stage_inst_dmem_n21028), .A2(MEM_stage_inst_dmem_n21027), .ZN(MEM_stage_inst_dmem_n8975) );
NAND2_X1 MEM_stage_inst_dmem_U20852 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n21036), .ZN(MEM_stage_inst_dmem_n21027) );
NAND2_X1 MEM_stage_inst_dmem_U20851 ( .A1(MEM_stage_inst_dmem_ram_3796), .A2(MEM_stage_inst_dmem_n21035), .ZN(MEM_stage_inst_dmem_n21028) );
NAND2_X1 MEM_stage_inst_dmem_U20850 ( .A1(MEM_stage_inst_dmem_n21026), .A2(MEM_stage_inst_dmem_n21025), .ZN(MEM_stage_inst_dmem_n8976) );
NAND2_X1 MEM_stage_inst_dmem_U20849 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n21036), .ZN(MEM_stage_inst_dmem_n21025) );
NAND2_X1 MEM_stage_inst_dmem_U20848 ( .A1(MEM_stage_inst_dmem_ram_3797), .A2(MEM_stage_inst_dmem_n21035), .ZN(MEM_stage_inst_dmem_n21026) );
NAND2_X1 MEM_stage_inst_dmem_U20847 ( .A1(MEM_stage_inst_dmem_n21024), .A2(MEM_stage_inst_dmem_n21023), .ZN(MEM_stage_inst_dmem_n8977) );
NAND2_X1 MEM_stage_inst_dmem_U20846 ( .A1(MEM_stage_inst_dmem_n21340), .A2(MEM_stage_inst_dmem_n21036), .ZN(MEM_stage_inst_dmem_n21023) );
NAND2_X1 MEM_stage_inst_dmem_U20845 ( .A1(MEM_stage_inst_dmem_ram_3798), .A2(MEM_stage_inst_dmem_n21035), .ZN(MEM_stage_inst_dmem_n21024) );
NAND2_X1 MEM_stage_inst_dmem_U20844 ( .A1(MEM_stage_inst_dmem_n21022), .A2(MEM_stage_inst_dmem_n21021), .ZN(MEM_stage_inst_dmem_n8978) );
NAND2_X1 MEM_stage_inst_dmem_U20843 ( .A1(MEM_stage_inst_dmem_n18), .A2(MEM_stage_inst_dmem_n21036), .ZN(MEM_stage_inst_dmem_n21021) );
NAND2_X1 MEM_stage_inst_dmem_U20842 ( .A1(MEM_stage_inst_dmem_ram_3799), .A2(MEM_stage_inst_dmem_n21035), .ZN(MEM_stage_inst_dmem_n21022) );
NAND2_X1 MEM_stage_inst_dmem_U20841 ( .A1(MEM_stage_inst_dmem_n21020), .A2(MEM_stage_inst_dmem_n21019), .ZN(MEM_stage_inst_dmem_n8979) );
NAND2_X1 MEM_stage_inst_dmem_U20840 ( .A1(MEM_stage_inst_dmem_n21335), .A2(MEM_stage_inst_dmem_n21036), .ZN(MEM_stage_inst_dmem_n21019) );
NAND2_X1 MEM_stage_inst_dmem_U20839 ( .A1(MEM_stage_inst_dmem_ram_3800), .A2(MEM_stage_inst_dmem_n21035), .ZN(MEM_stage_inst_dmem_n21020) );
NAND2_X1 MEM_stage_inst_dmem_U20838 ( .A1(MEM_stage_inst_dmem_n21018), .A2(MEM_stage_inst_dmem_n21017), .ZN(MEM_stage_inst_dmem_n8980) );
NAND2_X1 MEM_stage_inst_dmem_U20837 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n21036), .ZN(MEM_stage_inst_dmem_n21017) );
NAND2_X1 MEM_stage_inst_dmem_U20836 ( .A1(MEM_stage_inst_dmem_ram_3801), .A2(MEM_stage_inst_dmem_n21035), .ZN(MEM_stage_inst_dmem_n21018) );
NAND2_X1 MEM_stage_inst_dmem_U20835 ( .A1(MEM_stage_inst_dmem_n21016), .A2(MEM_stage_inst_dmem_n21015), .ZN(MEM_stage_inst_dmem_n8981) );
NAND2_X1 MEM_stage_inst_dmem_U20834 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n21036), .ZN(MEM_stage_inst_dmem_n21015) );
NAND2_X1 MEM_stage_inst_dmem_U20833 ( .A1(MEM_stage_inst_dmem_ram_3802), .A2(MEM_stage_inst_dmem_n21035), .ZN(MEM_stage_inst_dmem_n21016) );
NAND2_X1 MEM_stage_inst_dmem_U20832 ( .A1(MEM_stage_inst_dmem_n21014), .A2(MEM_stage_inst_dmem_n21013), .ZN(MEM_stage_inst_dmem_n8982) );
NAND2_X1 MEM_stage_inst_dmem_U20831 ( .A1(MEM_stage_inst_dmem_n13044), .A2(MEM_stage_inst_dmem_n21036), .ZN(MEM_stage_inst_dmem_n21013) );
NAND2_X1 MEM_stage_inst_dmem_U20830 ( .A1(MEM_stage_inst_dmem_ram_3803), .A2(MEM_stage_inst_dmem_n21035), .ZN(MEM_stage_inst_dmem_n21014) );
NAND2_X1 MEM_stage_inst_dmem_U20829 ( .A1(MEM_stage_inst_dmem_n21012), .A2(MEM_stage_inst_dmem_n21011), .ZN(MEM_stage_inst_dmem_n8983) );
NAND2_X1 MEM_stage_inst_dmem_U20828 ( .A1(MEM_stage_inst_dmem_n13041), .A2(MEM_stage_inst_dmem_n21036), .ZN(MEM_stage_inst_dmem_n21011) );
NAND2_X1 MEM_stage_inst_dmem_U20827 ( .A1(MEM_stage_inst_dmem_ram_3804), .A2(MEM_stage_inst_dmem_n21035), .ZN(MEM_stage_inst_dmem_n21012) );
NAND2_X1 MEM_stage_inst_dmem_U20826 ( .A1(MEM_stage_inst_dmem_n21010), .A2(MEM_stage_inst_dmem_n21009), .ZN(MEM_stage_inst_dmem_n8984) );
NAND2_X1 MEM_stage_inst_dmem_U20825 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n21036), .ZN(MEM_stage_inst_dmem_n21009) );
NAND2_X1 MEM_stage_inst_dmem_U20824 ( .A1(MEM_stage_inst_dmem_ram_3805), .A2(MEM_stage_inst_dmem_n21035), .ZN(MEM_stage_inst_dmem_n21010) );
NAND2_X1 MEM_stage_inst_dmem_U20823 ( .A1(MEM_stage_inst_dmem_n21008), .A2(MEM_stage_inst_dmem_n21007), .ZN(MEM_stage_inst_dmem_n8985) );
NAND2_X1 MEM_stage_inst_dmem_U20822 ( .A1(MEM_stage_inst_dmem_n115), .A2(MEM_stage_inst_dmem_n21036), .ZN(MEM_stage_inst_dmem_n21007) );
NAND2_X1 MEM_stage_inst_dmem_U20821 ( .A1(MEM_stage_inst_dmem_ram_3806), .A2(MEM_stage_inst_dmem_n21035), .ZN(MEM_stage_inst_dmem_n21008) );
NAND2_X1 MEM_stage_inst_dmem_U20820 ( .A1(MEM_stage_inst_dmem_n21006), .A2(MEM_stage_inst_dmem_n21005), .ZN(MEM_stage_inst_dmem_n8986) );
NAND2_X1 MEM_stage_inst_dmem_U20819 ( .A1(MEM_stage_inst_dmem_n21320), .A2(MEM_stage_inst_dmem_n21036), .ZN(MEM_stage_inst_dmem_n21005) );
INV_X1 MEM_stage_inst_dmem_U20818 ( .A(MEM_stage_inst_dmem_n21035), .ZN(MEM_stage_inst_dmem_n21036) );
NAND2_X1 MEM_stage_inst_dmem_U20817 ( .A1(MEM_stage_inst_dmem_ram_3807), .A2(MEM_stage_inst_dmem_n21035), .ZN(MEM_stage_inst_dmem_n21006) );
NAND2_X1 MEM_stage_inst_dmem_U20816 ( .A1(MEM_stage_inst_dmem_n21004), .A2(MEM_stage_inst_dmem_n21464), .ZN(MEM_stage_inst_dmem_n21035) );
NAND2_X1 MEM_stage_inst_dmem_U20815 ( .A1(MEM_stage_inst_dmem_n21003), .A2(MEM_stage_inst_dmem_n21002), .ZN(MEM_stage_inst_dmem_n8987) );
NAND2_X1 MEM_stage_inst_dmem_U20814 ( .A1(MEM_stage_inst_dmem_n20551), .A2(MEM_stage_inst_dmem_n21001), .ZN(MEM_stage_inst_dmem_n21002) );
NAND2_X1 MEM_stage_inst_dmem_U20813 ( .A1(MEM_stage_inst_dmem_ram_3808), .A2(MEM_stage_inst_dmem_n21000), .ZN(MEM_stage_inst_dmem_n21003) );
NAND2_X1 MEM_stage_inst_dmem_U20812 ( .A1(MEM_stage_inst_dmem_n20999), .A2(MEM_stage_inst_dmem_n20998), .ZN(MEM_stage_inst_dmem_n8988) );
NAND2_X1 MEM_stage_inst_dmem_U20811 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n21001), .ZN(MEM_stage_inst_dmem_n20998) );
NAND2_X1 MEM_stage_inst_dmem_U20810 ( .A1(MEM_stage_inst_dmem_ram_3809), .A2(MEM_stage_inst_dmem_n21000), .ZN(MEM_stage_inst_dmem_n20999) );
NAND2_X1 MEM_stage_inst_dmem_U20809 ( .A1(MEM_stage_inst_dmem_n20997), .A2(MEM_stage_inst_dmem_n20996), .ZN(MEM_stage_inst_dmem_n8989) );
NAND2_X1 MEM_stage_inst_dmem_U20808 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n21001), .ZN(MEM_stage_inst_dmem_n20996) );
NAND2_X1 MEM_stage_inst_dmem_U20807 ( .A1(MEM_stage_inst_dmem_ram_3810), .A2(MEM_stage_inst_dmem_n21000), .ZN(MEM_stage_inst_dmem_n20997) );
NAND2_X1 MEM_stage_inst_dmem_U20806 ( .A1(MEM_stage_inst_dmem_n20995), .A2(MEM_stage_inst_dmem_n20994), .ZN(MEM_stage_inst_dmem_n8990) );
NAND2_X1 MEM_stage_inst_dmem_U20805 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n21001), .ZN(MEM_stage_inst_dmem_n20994) );
NAND2_X1 MEM_stage_inst_dmem_U20804 ( .A1(MEM_stage_inst_dmem_ram_3811), .A2(MEM_stage_inst_dmem_n21000), .ZN(MEM_stage_inst_dmem_n20995) );
NAND2_X1 MEM_stage_inst_dmem_U20803 ( .A1(MEM_stage_inst_dmem_n20993), .A2(MEM_stage_inst_dmem_n20992), .ZN(MEM_stage_inst_dmem_n8991) );
NAND2_X1 MEM_stage_inst_dmem_U20802 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n21001), .ZN(MEM_stage_inst_dmem_n20992) );
NAND2_X1 MEM_stage_inst_dmem_U20801 ( .A1(MEM_stage_inst_dmem_ram_3812), .A2(MEM_stage_inst_dmem_n21000), .ZN(MEM_stage_inst_dmem_n20993) );
NAND2_X1 MEM_stage_inst_dmem_U20800 ( .A1(MEM_stage_inst_dmem_n20991), .A2(MEM_stage_inst_dmem_n20990), .ZN(MEM_stage_inst_dmem_n8992) );
NAND2_X1 MEM_stage_inst_dmem_U20799 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n21001), .ZN(MEM_stage_inst_dmem_n20990) );
NAND2_X1 MEM_stage_inst_dmem_U20798 ( .A1(MEM_stage_inst_dmem_ram_3813), .A2(MEM_stage_inst_dmem_n21000), .ZN(MEM_stage_inst_dmem_n20991) );
NAND2_X1 MEM_stage_inst_dmem_U20797 ( .A1(MEM_stage_inst_dmem_n20989), .A2(MEM_stage_inst_dmem_n20988), .ZN(MEM_stage_inst_dmem_n8993) );
NAND2_X1 MEM_stage_inst_dmem_U20796 ( .A1(MEM_stage_inst_dmem_n21340), .A2(MEM_stage_inst_dmem_n21001), .ZN(MEM_stage_inst_dmem_n20988) );
NAND2_X1 MEM_stage_inst_dmem_U20795 ( .A1(MEM_stage_inst_dmem_ram_3814), .A2(MEM_stage_inst_dmem_n21000), .ZN(MEM_stage_inst_dmem_n20989) );
NAND2_X1 MEM_stage_inst_dmem_U20794 ( .A1(MEM_stage_inst_dmem_n20987), .A2(MEM_stage_inst_dmem_n20986), .ZN(MEM_stage_inst_dmem_n8994) );
NAND2_X1 MEM_stage_inst_dmem_U20793 ( .A1(MEM_stage_inst_dmem_n17), .A2(MEM_stage_inst_dmem_n21001), .ZN(MEM_stage_inst_dmem_n20986) );
NAND2_X1 MEM_stage_inst_dmem_U20792 ( .A1(MEM_stage_inst_dmem_ram_3815), .A2(MEM_stage_inst_dmem_n21000), .ZN(MEM_stage_inst_dmem_n20987) );
NAND2_X1 MEM_stage_inst_dmem_U20791 ( .A1(MEM_stage_inst_dmem_n20985), .A2(MEM_stage_inst_dmem_n20984), .ZN(MEM_stage_inst_dmem_n8995) );
NAND2_X1 MEM_stage_inst_dmem_U20790 ( .A1(MEM_stage_inst_dmem_n21335), .A2(MEM_stage_inst_dmem_n21001), .ZN(MEM_stage_inst_dmem_n20984) );
NAND2_X1 MEM_stage_inst_dmem_U20789 ( .A1(MEM_stage_inst_dmem_ram_3816), .A2(MEM_stage_inst_dmem_n21000), .ZN(MEM_stage_inst_dmem_n20985) );
NAND2_X1 MEM_stage_inst_dmem_U20788 ( .A1(MEM_stage_inst_dmem_n20983), .A2(MEM_stage_inst_dmem_n20982), .ZN(MEM_stage_inst_dmem_n8996) );
NAND2_X1 MEM_stage_inst_dmem_U20787 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n21001), .ZN(MEM_stage_inst_dmem_n20982) );
NAND2_X1 MEM_stage_inst_dmem_U20786 ( .A1(MEM_stage_inst_dmem_ram_3817), .A2(MEM_stage_inst_dmem_n21000), .ZN(MEM_stage_inst_dmem_n20983) );
NAND2_X1 MEM_stage_inst_dmem_U20785 ( .A1(MEM_stage_inst_dmem_n20981), .A2(MEM_stage_inst_dmem_n20980), .ZN(MEM_stage_inst_dmem_n8997) );
NAND2_X1 MEM_stage_inst_dmem_U20784 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n21001), .ZN(MEM_stage_inst_dmem_n20980) );
NAND2_X1 MEM_stage_inst_dmem_U20783 ( .A1(MEM_stage_inst_dmem_ram_3818), .A2(MEM_stage_inst_dmem_n21000), .ZN(MEM_stage_inst_dmem_n20981) );
NAND2_X1 MEM_stage_inst_dmem_U20782 ( .A1(MEM_stage_inst_dmem_n20979), .A2(MEM_stage_inst_dmem_n20978), .ZN(MEM_stage_inst_dmem_n8998) );
NAND2_X1 MEM_stage_inst_dmem_U20781 ( .A1(MEM_stage_inst_dmem_n14705), .A2(MEM_stage_inst_dmem_n21001), .ZN(MEM_stage_inst_dmem_n20978) );
NAND2_X1 MEM_stage_inst_dmem_U20780 ( .A1(MEM_stage_inst_dmem_ram_3819), .A2(MEM_stage_inst_dmem_n21000), .ZN(MEM_stage_inst_dmem_n20979) );
NAND2_X1 MEM_stage_inst_dmem_U20779 ( .A1(MEM_stage_inst_dmem_n20977), .A2(MEM_stage_inst_dmem_n20976), .ZN(MEM_stage_inst_dmem_n8999) );
NAND2_X1 MEM_stage_inst_dmem_U20778 ( .A1(MEM_stage_inst_dmem_n14702), .A2(MEM_stage_inst_dmem_n21001), .ZN(MEM_stage_inst_dmem_n20976) );
NAND2_X1 MEM_stage_inst_dmem_U20777 ( .A1(MEM_stage_inst_dmem_ram_3820), .A2(MEM_stage_inst_dmem_n21000), .ZN(MEM_stage_inst_dmem_n20977) );
NAND2_X1 MEM_stage_inst_dmem_U20776 ( .A1(MEM_stage_inst_dmem_n20975), .A2(MEM_stage_inst_dmem_n20974), .ZN(MEM_stage_inst_dmem_n9000) );
NAND2_X1 MEM_stage_inst_dmem_U20775 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n21001), .ZN(MEM_stage_inst_dmem_n20974) );
NAND2_X1 MEM_stage_inst_dmem_U20774 ( .A1(MEM_stage_inst_dmem_ram_3821), .A2(MEM_stage_inst_dmem_n21000), .ZN(MEM_stage_inst_dmem_n20975) );
NAND2_X1 MEM_stage_inst_dmem_U20773 ( .A1(MEM_stage_inst_dmem_n20973), .A2(MEM_stage_inst_dmem_n20972), .ZN(MEM_stage_inst_dmem_n9001) );
NAND2_X1 MEM_stage_inst_dmem_U20772 ( .A1(MEM_stage_inst_dmem_n20509), .A2(MEM_stage_inst_dmem_n21001), .ZN(MEM_stage_inst_dmem_n20972) );
NAND2_X1 MEM_stage_inst_dmem_U20771 ( .A1(MEM_stage_inst_dmem_ram_3822), .A2(MEM_stage_inst_dmem_n21000), .ZN(MEM_stage_inst_dmem_n20973) );
NAND2_X1 MEM_stage_inst_dmem_U20770 ( .A1(MEM_stage_inst_dmem_n20971), .A2(MEM_stage_inst_dmem_n20970), .ZN(MEM_stage_inst_dmem_n9002) );
NAND2_X1 MEM_stage_inst_dmem_U20769 ( .A1(MEM_stage_inst_dmem_n21320), .A2(MEM_stage_inst_dmem_n21001), .ZN(MEM_stage_inst_dmem_n20970) );
INV_X1 MEM_stage_inst_dmem_U20768 ( .A(MEM_stage_inst_dmem_n21000), .ZN(MEM_stage_inst_dmem_n21001) );
NAND2_X1 MEM_stage_inst_dmem_U20767 ( .A1(MEM_stage_inst_dmem_ram_3823), .A2(MEM_stage_inst_dmem_n21000), .ZN(MEM_stage_inst_dmem_n20971) );
NAND2_X1 MEM_stage_inst_dmem_U20766 ( .A1(MEM_stage_inst_dmem_n20969), .A2(MEM_stage_inst_dmem_n21464), .ZN(MEM_stage_inst_dmem_n21000) );
NAND2_X1 MEM_stage_inst_dmem_U20765 ( .A1(MEM_stage_inst_dmem_n20968), .A2(MEM_stage_inst_dmem_n20967), .ZN(MEM_stage_inst_dmem_n9003) );
NAND2_X1 MEM_stage_inst_dmem_U20764 ( .A1(EX_pipeline_reg_out_5), .A2(MEM_stage_inst_dmem_n20966), .ZN(MEM_stage_inst_dmem_n20967) );
NAND2_X1 MEM_stage_inst_dmem_U20763 ( .A1(MEM_stage_inst_dmem_ram_3824), .A2(MEM_stage_inst_dmem_n20965), .ZN(MEM_stage_inst_dmem_n20968) );
NAND2_X1 MEM_stage_inst_dmem_U20762 ( .A1(MEM_stage_inst_dmem_n20964), .A2(MEM_stage_inst_dmem_n20963), .ZN(MEM_stage_inst_dmem_n9004) );
NAND2_X1 MEM_stage_inst_dmem_U20761 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n20966), .ZN(MEM_stage_inst_dmem_n20963) );
NAND2_X1 MEM_stage_inst_dmem_U20760 ( .A1(MEM_stage_inst_dmem_ram_3825), .A2(MEM_stage_inst_dmem_n20965), .ZN(MEM_stage_inst_dmem_n20964) );
NAND2_X1 MEM_stage_inst_dmem_U20759 ( .A1(MEM_stage_inst_dmem_n20962), .A2(MEM_stage_inst_dmem_n20961), .ZN(MEM_stage_inst_dmem_n9005) );
NAND2_X1 MEM_stage_inst_dmem_U20758 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n20966), .ZN(MEM_stage_inst_dmem_n20961) );
NAND2_X1 MEM_stage_inst_dmem_U20757 ( .A1(MEM_stage_inst_dmem_ram_3826), .A2(MEM_stage_inst_dmem_n20965), .ZN(MEM_stage_inst_dmem_n20962) );
NAND2_X1 MEM_stage_inst_dmem_U20756 ( .A1(MEM_stage_inst_dmem_n20960), .A2(MEM_stage_inst_dmem_n20959), .ZN(MEM_stage_inst_dmem_n9006) );
NAND2_X1 MEM_stage_inst_dmem_U20755 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n20966), .ZN(MEM_stage_inst_dmem_n20959) );
NAND2_X1 MEM_stage_inst_dmem_U20754 ( .A1(MEM_stage_inst_dmem_ram_3827), .A2(MEM_stage_inst_dmem_n20965), .ZN(MEM_stage_inst_dmem_n20960) );
NAND2_X1 MEM_stage_inst_dmem_U20753 ( .A1(MEM_stage_inst_dmem_n20958), .A2(MEM_stage_inst_dmem_n20957), .ZN(MEM_stage_inst_dmem_n9007) );
NAND2_X1 MEM_stage_inst_dmem_U20752 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n20966), .ZN(MEM_stage_inst_dmem_n20957) );
NAND2_X1 MEM_stage_inst_dmem_U20751 ( .A1(MEM_stage_inst_dmem_ram_3828), .A2(MEM_stage_inst_dmem_n20965), .ZN(MEM_stage_inst_dmem_n20958) );
NAND2_X1 MEM_stage_inst_dmem_U20750 ( .A1(MEM_stage_inst_dmem_n20956), .A2(MEM_stage_inst_dmem_n20955), .ZN(MEM_stage_inst_dmem_n9008) );
NAND2_X1 MEM_stage_inst_dmem_U20749 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n20966), .ZN(MEM_stage_inst_dmem_n20955) );
NAND2_X1 MEM_stage_inst_dmem_U20748 ( .A1(MEM_stage_inst_dmem_ram_3829), .A2(MEM_stage_inst_dmem_n20965), .ZN(MEM_stage_inst_dmem_n20956) );
NAND2_X1 MEM_stage_inst_dmem_U20747 ( .A1(MEM_stage_inst_dmem_n20954), .A2(MEM_stage_inst_dmem_n20953), .ZN(MEM_stage_inst_dmem_n9009) );
NAND2_X1 MEM_stage_inst_dmem_U20746 ( .A1(MEM_stage_inst_dmem_n21340), .A2(MEM_stage_inst_dmem_n20966), .ZN(MEM_stage_inst_dmem_n20953) );
NAND2_X1 MEM_stage_inst_dmem_U20745 ( .A1(MEM_stage_inst_dmem_ram_3830), .A2(MEM_stage_inst_dmem_n20965), .ZN(MEM_stage_inst_dmem_n20954) );
NAND2_X1 MEM_stage_inst_dmem_U20744 ( .A1(MEM_stage_inst_dmem_n20952), .A2(MEM_stage_inst_dmem_n20951), .ZN(MEM_stage_inst_dmem_n9010) );
NAND2_X1 MEM_stage_inst_dmem_U20743 ( .A1(MEM_stage_inst_dmem_n18), .A2(MEM_stage_inst_dmem_n20966), .ZN(MEM_stage_inst_dmem_n20951) );
NAND2_X1 MEM_stage_inst_dmem_U20742 ( .A1(MEM_stage_inst_dmem_ram_3831), .A2(MEM_stage_inst_dmem_n20965), .ZN(MEM_stage_inst_dmem_n20952) );
NAND2_X1 MEM_stage_inst_dmem_U20741 ( .A1(MEM_stage_inst_dmem_n20950), .A2(MEM_stage_inst_dmem_n20949), .ZN(MEM_stage_inst_dmem_n9011) );
NAND2_X1 MEM_stage_inst_dmem_U20740 ( .A1(MEM_stage_inst_dmem_n21335), .A2(MEM_stage_inst_dmem_n20966), .ZN(MEM_stage_inst_dmem_n20949) );
NAND2_X1 MEM_stage_inst_dmem_U20739 ( .A1(MEM_stage_inst_dmem_ram_3832), .A2(MEM_stage_inst_dmem_n20965), .ZN(MEM_stage_inst_dmem_n20950) );
NAND2_X1 MEM_stage_inst_dmem_U20738 ( .A1(MEM_stage_inst_dmem_n20948), .A2(MEM_stage_inst_dmem_n20947), .ZN(MEM_stage_inst_dmem_n9012) );
NAND2_X1 MEM_stage_inst_dmem_U20737 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n20966), .ZN(MEM_stage_inst_dmem_n20947) );
NAND2_X1 MEM_stage_inst_dmem_U20736 ( .A1(MEM_stage_inst_dmem_ram_3833), .A2(MEM_stage_inst_dmem_n20965), .ZN(MEM_stage_inst_dmem_n20948) );
NAND2_X1 MEM_stage_inst_dmem_U20735 ( .A1(MEM_stage_inst_dmem_n20946), .A2(MEM_stage_inst_dmem_n20945), .ZN(MEM_stage_inst_dmem_n9013) );
NAND2_X1 MEM_stage_inst_dmem_U20734 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n20966), .ZN(MEM_stage_inst_dmem_n20945) );
NAND2_X1 MEM_stage_inst_dmem_U20733 ( .A1(MEM_stage_inst_dmem_ram_3834), .A2(MEM_stage_inst_dmem_n20965), .ZN(MEM_stage_inst_dmem_n20946) );
NAND2_X1 MEM_stage_inst_dmem_U20732 ( .A1(MEM_stage_inst_dmem_n20944), .A2(MEM_stage_inst_dmem_n20943), .ZN(MEM_stage_inst_dmem_n9014) );
NAND2_X1 MEM_stage_inst_dmem_U20731 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n20966), .ZN(MEM_stage_inst_dmem_n20943) );
NAND2_X1 MEM_stage_inst_dmem_U20730 ( .A1(MEM_stage_inst_dmem_ram_3835), .A2(MEM_stage_inst_dmem_n20965), .ZN(MEM_stage_inst_dmem_n20944) );
NAND2_X1 MEM_stage_inst_dmem_U20729 ( .A1(MEM_stage_inst_dmem_n20942), .A2(MEM_stage_inst_dmem_n20941), .ZN(MEM_stage_inst_dmem_n9015) );
NAND2_X1 MEM_stage_inst_dmem_U20728 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n20966), .ZN(MEM_stage_inst_dmem_n20941) );
NAND2_X1 MEM_stage_inst_dmem_U20727 ( .A1(MEM_stage_inst_dmem_ram_3836), .A2(MEM_stage_inst_dmem_n20965), .ZN(MEM_stage_inst_dmem_n20942) );
NAND2_X1 MEM_stage_inst_dmem_U20726 ( .A1(MEM_stage_inst_dmem_n20940), .A2(MEM_stage_inst_dmem_n20939), .ZN(MEM_stage_inst_dmem_n9016) );
NAND2_X1 MEM_stage_inst_dmem_U20725 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n20966), .ZN(MEM_stage_inst_dmem_n20939) );
NAND2_X1 MEM_stage_inst_dmem_U20724 ( .A1(MEM_stage_inst_dmem_ram_3837), .A2(MEM_stage_inst_dmem_n20965), .ZN(MEM_stage_inst_dmem_n20940) );
NAND2_X1 MEM_stage_inst_dmem_U20723 ( .A1(MEM_stage_inst_dmem_n20938), .A2(MEM_stage_inst_dmem_n20937), .ZN(MEM_stage_inst_dmem_n9017) );
NAND2_X1 MEM_stage_inst_dmem_U20722 ( .A1(EX_pipeline_reg_out_19), .A2(MEM_stage_inst_dmem_n20966), .ZN(MEM_stage_inst_dmem_n20937) );
NAND2_X1 MEM_stage_inst_dmem_U20721 ( .A1(MEM_stage_inst_dmem_ram_3838), .A2(MEM_stage_inst_dmem_n20965), .ZN(MEM_stage_inst_dmem_n20938) );
NAND2_X1 MEM_stage_inst_dmem_U20720 ( .A1(MEM_stage_inst_dmem_n20936), .A2(MEM_stage_inst_dmem_n20935), .ZN(MEM_stage_inst_dmem_n9018) );
NAND2_X1 MEM_stage_inst_dmem_U20719 ( .A1(MEM_stage_inst_dmem_n21320), .A2(MEM_stage_inst_dmem_n20966), .ZN(MEM_stage_inst_dmem_n20935) );
INV_X1 MEM_stage_inst_dmem_U20718 ( .A(MEM_stage_inst_dmem_n20965), .ZN(MEM_stage_inst_dmem_n20966) );
NAND2_X1 MEM_stage_inst_dmem_U20717 ( .A1(MEM_stage_inst_dmem_ram_3839), .A2(MEM_stage_inst_dmem_n20965), .ZN(MEM_stage_inst_dmem_n20936) );
NAND2_X1 MEM_stage_inst_dmem_U20716 ( .A1(MEM_stage_inst_dmem_n20934), .A2(MEM_stage_inst_dmem_n21464), .ZN(MEM_stage_inst_dmem_n20965) );
NOR2_X2 MEM_stage_inst_dmem_U20715 ( .A1(MEM_stage_inst_dmem_n20933), .A2(MEM_stage_inst_dmem_n20932), .ZN(MEM_stage_inst_dmem_n21464) );
NAND2_X1 MEM_stage_inst_dmem_U20714 ( .A1(MEM_stage_inst_dmem_n20931), .A2(MEM_stage_inst_dmem_n20930), .ZN(MEM_stage_inst_dmem_n9019) );
NAND2_X1 MEM_stage_inst_dmem_U20713 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n20929), .ZN(MEM_stage_inst_dmem_n20930) );
NAND2_X1 MEM_stage_inst_dmem_U20712 ( .A1(MEM_stage_inst_dmem_ram_3840), .A2(MEM_stage_inst_dmem_n20928), .ZN(MEM_stage_inst_dmem_n20931) );
NAND2_X1 MEM_stage_inst_dmem_U20711 ( .A1(MEM_stage_inst_dmem_n20927), .A2(MEM_stage_inst_dmem_n20926), .ZN(MEM_stage_inst_dmem_n9020) );
NAND2_X1 MEM_stage_inst_dmem_U20710 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n20929), .ZN(MEM_stage_inst_dmem_n20926) );
NAND2_X1 MEM_stage_inst_dmem_U20709 ( .A1(MEM_stage_inst_dmem_ram_3841), .A2(MEM_stage_inst_dmem_n20928), .ZN(MEM_stage_inst_dmem_n20927) );
NAND2_X1 MEM_stage_inst_dmem_U20708 ( .A1(MEM_stage_inst_dmem_n20925), .A2(MEM_stage_inst_dmem_n20924), .ZN(MEM_stage_inst_dmem_n9021) );
NAND2_X1 MEM_stage_inst_dmem_U20707 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n20929), .ZN(MEM_stage_inst_dmem_n20924) );
NAND2_X1 MEM_stage_inst_dmem_U20706 ( .A1(MEM_stage_inst_dmem_ram_3842), .A2(MEM_stage_inst_dmem_n20928), .ZN(MEM_stage_inst_dmem_n20925) );
NAND2_X1 MEM_stage_inst_dmem_U20705 ( .A1(MEM_stage_inst_dmem_n20923), .A2(MEM_stage_inst_dmem_n20922), .ZN(MEM_stage_inst_dmem_n9022) );
NAND2_X1 MEM_stage_inst_dmem_U20704 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n20929), .ZN(MEM_stage_inst_dmem_n20922) );
NAND2_X1 MEM_stage_inst_dmem_U20703 ( .A1(MEM_stage_inst_dmem_ram_3843), .A2(MEM_stage_inst_dmem_n20928), .ZN(MEM_stage_inst_dmem_n20923) );
NAND2_X1 MEM_stage_inst_dmem_U20702 ( .A1(MEM_stage_inst_dmem_n20921), .A2(MEM_stage_inst_dmem_n20920), .ZN(MEM_stage_inst_dmem_n9023) );
NAND2_X1 MEM_stage_inst_dmem_U20701 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n20929), .ZN(MEM_stage_inst_dmem_n20920) );
NAND2_X1 MEM_stage_inst_dmem_U20700 ( .A1(MEM_stage_inst_dmem_ram_3844), .A2(MEM_stage_inst_dmem_n20928), .ZN(MEM_stage_inst_dmem_n20921) );
NAND2_X1 MEM_stage_inst_dmem_U20699 ( .A1(MEM_stage_inst_dmem_n20918), .A2(MEM_stage_inst_dmem_n20917), .ZN(MEM_stage_inst_dmem_n9024) );
NAND2_X1 MEM_stage_inst_dmem_U20698 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n20929), .ZN(MEM_stage_inst_dmem_n20917) );
NAND2_X1 MEM_stage_inst_dmem_U20697 ( .A1(MEM_stage_inst_dmem_ram_3845), .A2(MEM_stage_inst_dmem_n20928), .ZN(MEM_stage_inst_dmem_n20918) );
NAND2_X1 MEM_stage_inst_dmem_U20696 ( .A1(MEM_stage_inst_dmem_n20916), .A2(MEM_stage_inst_dmem_n20915), .ZN(MEM_stage_inst_dmem_n9025) );
NAND2_X1 MEM_stage_inst_dmem_U20695 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n20929), .ZN(MEM_stage_inst_dmem_n20915) );
NAND2_X1 MEM_stage_inst_dmem_U20694 ( .A1(MEM_stage_inst_dmem_ram_3846), .A2(MEM_stage_inst_dmem_n20928), .ZN(MEM_stage_inst_dmem_n20916) );
NAND2_X1 MEM_stage_inst_dmem_U20693 ( .A1(MEM_stage_inst_dmem_n20914), .A2(MEM_stage_inst_dmem_n20913), .ZN(MEM_stage_inst_dmem_n9026) );
NAND2_X1 MEM_stage_inst_dmem_U20692 ( .A1(MEM_stage_inst_dmem_n17), .A2(MEM_stage_inst_dmem_n20929), .ZN(MEM_stage_inst_dmem_n20913) );
NAND2_X1 MEM_stage_inst_dmem_U20691 ( .A1(MEM_stage_inst_dmem_ram_3847), .A2(MEM_stage_inst_dmem_n20928), .ZN(MEM_stage_inst_dmem_n20914) );
NAND2_X1 MEM_stage_inst_dmem_U20690 ( .A1(MEM_stage_inst_dmem_n20912), .A2(MEM_stage_inst_dmem_n20911), .ZN(MEM_stage_inst_dmem_n9027) );
NAND2_X1 MEM_stage_inst_dmem_U20689 ( .A1(MEM_stage_inst_dmem_n13051), .A2(MEM_stage_inst_dmem_n20929), .ZN(MEM_stage_inst_dmem_n20911) );
NAND2_X1 MEM_stage_inst_dmem_U20688 ( .A1(MEM_stage_inst_dmem_ram_3848), .A2(MEM_stage_inst_dmem_n20928), .ZN(MEM_stage_inst_dmem_n20912) );
NAND2_X1 MEM_stage_inst_dmem_U20687 ( .A1(MEM_stage_inst_dmem_n20910), .A2(MEM_stage_inst_dmem_n20909), .ZN(MEM_stage_inst_dmem_n9028) );
NAND2_X1 MEM_stage_inst_dmem_U20686 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n20929), .ZN(MEM_stage_inst_dmem_n20909) );
NAND2_X1 MEM_stage_inst_dmem_U20685 ( .A1(MEM_stage_inst_dmem_ram_3849), .A2(MEM_stage_inst_dmem_n20928), .ZN(MEM_stage_inst_dmem_n20910) );
NAND2_X1 MEM_stage_inst_dmem_U20684 ( .A1(MEM_stage_inst_dmem_n20908), .A2(MEM_stage_inst_dmem_n20907), .ZN(MEM_stage_inst_dmem_n9029) );
NAND2_X1 MEM_stage_inst_dmem_U20683 ( .A1(MEM_stage_inst_dmem_n18867), .A2(MEM_stage_inst_dmem_n20929), .ZN(MEM_stage_inst_dmem_n20907) );
NAND2_X1 MEM_stage_inst_dmem_U20682 ( .A1(MEM_stage_inst_dmem_ram_3850), .A2(MEM_stage_inst_dmem_n20928), .ZN(MEM_stage_inst_dmem_n20908) );
NAND2_X1 MEM_stage_inst_dmem_U20681 ( .A1(MEM_stage_inst_dmem_n20906), .A2(MEM_stage_inst_dmem_n20905), .ZN(MEM_stage_inst_dmem_n9030) );
NAND2_X1 MEM_stage_inst_dmem_U20680 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n20929), .ZN(MEM_stage_inst_dmem_n20905) );
NAND2_X1 MEM_stage_inst_dmem_U20679 ( .A1(MEM_stage_inst_dmem_ram_3851), .A2(MEM_stage_inst_dmem_n20928), .ZN(MEM_stage_inst_dmem_n20906) );
NAND2_X1 MEM_stage_inst_dmem_U20678 ( .A1(MEM_stage_inst_dmem_n20903), .A2(MEM_stage_inst_dmem_n20902), .ZN(MEM_stage_inst_dmem_n9031) );
NAND2_X1 MEM_stage_inst_dmem_U20677 ( .A1(MEM_stage_inst_dmem_n14702), .A2(MEM_stage_inst_dmem_n20929), .ZN(MEM_stage_inst_dmem_n20902) );
NAND2_X1 MEM_stage_inst_dmem_U20676 ( .A1(MEM_stage_inst_dmem_ram_3852), .A2(MEM_stage_inst_dmem_n20928), .ZN(MEM_stage_inst_dmem_n20903) );
NAND2_X1 MEM_stage_inst_dmem_U20675 ( .A1(MEM_stage_inst_dmem_n20901), .A2(MEM_stage_inst_dmem_n20900), .ZN(MEM_stage_inst_dmem_n9032) );
NAND2_X1 MEM_stage_inst_dmem_U20674 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n20929), .ZN(MEM_stage_inst_dmem_n20900) );
NAND2_X1 MEM_stage_inst_dmem_U20673 ( .A1(MEM_stage_inst_dmem_ram_3853), .A2(MEM_stage_inst_dmem_n20928), .ZN(MEM_stage_inst_dmem_n20901) );
NAND2_X1 MEM_stage_inst_dmem_U20672 ( .A1(MEM_stage_inst_dmem_n20899), .A2(MEM_stage_inst_dmem_n20898), .ZN(MEM_stage_inst_dmem_n9033) );
NAND2_X1 MEM_stage_inst_dmem_U20671 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n20929), .ZN(MEM_stage_inst_dmem_n20898) );
NAND2_X1 MEM_stage_inst_dmem_U20670 ( .A1(MEM_stage_inst_dmem_ram_3854), .A2(MEM_stage_inst_dmem_n20928), .ZN(MEM_stage_inst_dmem_n20899) );
NAND2_X1 MEM_stage_inst_dmem_U20669 ( .A1(MEM_stage_inst_dmem_n20897), .A2(MEM_stage_inst_dmem_n20896), .ZN(MEM_stage_inst_dmem_n9034) );
NAND2_X1 MEM_stage_inst_dmem_U20668 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n20929), .ZN(MEM_stage_inst_dmem_n20896) );
INV_X1 MEM_stage_inst_dmem_U20667 ( .A(MEM_stage_inst_dmem_n20928), .ZN(MEM_stage_inst_dmem_n20929) );
NAND2_X1 MEM_stage_inst_dmem_U20666 ( .A1(MEM_stage_inst_dmem_ram_3855), .A2(MEM_stage_inst_dmem_n20928), .ZN(MEM_stage_inst_dmem_n20897) );
NAND2_X1 MEM_stage_inst_dmem_U20665 ( .A1(MEM_stage_inst_dmem_n21465), .A2(MEM_stage_inst_dmem_n20895), .ZN(MEM_stage_inst_dmem_n20928) );
NAND2_X1 MEM_stage_inst_dmem_U20664 ( .A1(MEM_stage_inst_dmem_n20894), .A2(MEM_stage_inst_dmem_n20893), .ZN(MEM_stage_inst_dmem_n9035) );
NAND2_X1 MEM_stage_inst_dmem_U20663 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n20892), .ZN(MEM_stage_inst_dmem_n20893) );
NAND2_X1 MEM_stage_inst_dmem_U20662 ( .A1(MEM_stage_inst_dmem_ram_3856), .A2(MEM_stage_inst_dmem_n20891), .ZN(MEM_stage_inst_dmem_n20894) );
NAND2_X1 MEM_stage_inst_dmem_U20661 ( .A1(MEM_stage_inst_dmem_n20890), .A2(MEM_stage_inst_dmem_n20889), .ZN(MEM_stage_inst_dmem_n9036) );
NAND2_X1 MEM_stage_inst_dmem_U20660 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n20892), .ZN(MEM_stage_inst_dmem_n20889) );
NAND2_X1 MEM_stage_inst_dmem_U20659 ( .A1(MEM_stage_inst_dmem_ram_3857), .A2(MEM_stage_inst_dmem_n20891), .ZN(MEM_stage_inst_dmem_n20890) );
NAND2_X1 MEM_stage_inst_dmem_U20658 ( .A1(MEM_stage_inst_dmem_n20888), .A2(MEM_stage_inst_dmem_n20887), .ZN(MEM_stage_inst_dmem_n9037) );
NAND2_X1 MEM_stage_inst_dmem_U20657 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n20892), .ZN(MEM_stage_inst_dmem_n20887) );
NAND2_X1 MEM_stage_inst_dmem_U20656 ( .A1(MEM_stage_inst_dmem_ram_3858), .A2(MEM_stage_inst_dmem_n20891), .ZN(MEM_stage_inst_dmem_n20888) );
NAND2_X1 MEM_stage_inst_dmem_U20655 ( .A1(MEM_stage_inst_dmem_n20886), .A2(MEM_stage_inst_dmem_n20885), .ZN(MEM_stage_inst_dmem_n9038) );
NAND2_X1 MEM_stage_inst_dmem_U20654 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n20892), .ZN(MEM_stage_inst_dmem_n20885) );
NAND2_X1 MEM_stage_inst_dmem_U20653 ( .A1(MEM_stage_inst_dmem_ram_3859), .A2(MEM_stage_inst_dmem_n20891), .ZN(MEM_stage_inst_dmem_n20886) );
NAND2_X1 MEM_stage_inst_dmem_U20652 ( .A1(MEM_stage_inst_dmem_n20884), .A2(MEM_stage_inst_dmem_n20883), .ZN(MEM_stage_inst_dmem_n9039) );
NAND2_X1 MEM_stage_inst_dmem_U20651 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n20892), .ZN(MEM_stage_inst_dmem_n20883) );
NAND2_X1 MEM_stage_inst_dmem_U20650 ( .A1(MEM_stage_inst_dmem_ram_3860), .A2(MEM_stage_inst_dmem_n20891), .ZN(MEM_stage_inst_dmem_n20884) );
NAND2_X1 MEM_stage_inst_dmem_U20649 ( .A1(MEM_stage_inst_dmem_n20882), .A2(MEM_stage_inst_dmem_n20881), .ZN(MEM_stage_inst_dmem_n9040) );
NAND2_X1 MEM_stage_inst_dmem_U20648 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n20892), .ZN(MEM_stage_inst_dmem_n20881) );
NAND2_X1 MEM_stage_inst_dmem_U20647 ( .A1(MEM_stage_inst_dmem_ram_3861), .A2(MEM_stage_inst_dmem_n20891), .ZN(MEM_stage_inst_dmem_n20882) );
NAND2_X1 MEM_stage_inst_dmem_U20646 ( .A1(MEM_stage_inst_dmem_n20880), .A2(MEM_stage_inst_dmem_n20879), .ZN(MEM_stage_inst_dmem_n9041) );
NAND2_X1 MEM_stage_inst_dmem_U20645 ( .A1(MEM_stage_inst_dmem_n14717), .A2(MEM_stage_inst_dmem_n20892), .ZN(MEM_stage_inst_dmem_n20879) );
NAND2_X1 MEM_stage_inst_dmem_U20644 ( .A1(MEM_stage_inst_dmem_ram_3862), .A2(MEM_stage_inst_dmem_n20891), .ZN(MEM_stage_inst_dmem_n20880) );
NAND2_X1 MEM_stage_inst_dmem_U20643 ( .A1(MEM_stage_inst_dmem_n20878), .A2(MEM_stage_inst_dmem_n20877), .ZN(MEM_stage_inst_dmem_n9042) );
NAND2_X1 MEM_stage_inst_dmem_U20642 ( .A1(EX_pipeline_reg_out_12), .A2(MEM_stage_inst_dmem_n20892), .ZN(MEM_stage_inst_dmem_n20877) );
NAND2_X1 MEM_stage_inst_dmem_U20641 ( .A1(MEM_stage_inst_dmem_ram_3863), .A2(MEM_stage_inst_dmem_n20891), .ZN(MEM_stage_inst_dmem_n20878) );
NAND2_X1 MEM_stage_inst_dmem_U20640 ( .A1(MEM_stage_inst_dmem_n20876), .A2(MEM_stage_inst_dmem_n20875), .ZN(MEM_stage_inst_dmem_n9043) );
NAND2_X1 MEM_stage_inst_dmem_U20639 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n20892), .ZN(MEM_stage_inst_dmem_n20875) );
NAND2_X1 MEM_stage_inst_dmem_U20638 ( .A1(MEM_stage_inst_dmem_ram_3864), .A2(MEM_stage_inst_dmem_n20891), .ZN(MEM_stage_inst_dmem_n20876) );
NAND2_X1 MEM_stage_inst_dmem_U20637 ( .A1(MEM_stage_inst_dmem_n20874), .A2(MEM_stage_inst_dmem_n20873), .ZN(MEM_stage_inst_dmem_n9044) );
NAND2_X1 MEM_stage_inst_dmem_U20636 ( .A1(MEM_stage_inst_dmem_n96), .A2(MEM_stage_inst_dmem_n20892), .ZN(MEM_stage_inst_dmem_n20873) );
NAND2_X1 MEM_stage_inst_dmem_U20635 ( .A1(MEM_stage_inst_dmem_ram_3865), .A2(MEM_stage_inst_dmem_n20891), .ZN(MEM_stage_inst_dmem_n20874) );
NAND2_X1 MEM_stage_inst_dmem_U20634 ( .A1(MEM_stage_inst_dmem_n20872), .A2(MEM_stage_inst_dmem_n20871), .ZN(MEM_stage_inst_dmem_n9045) );
NAND2_X1 MEM_stage_inst_dmem_U20633 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n20892), .ZN(MEM_stage_inst_dmem_n20871) );
NAND2_X1 MEM_stage_inst_dmem_U20632 ( .A1(MEM_stage_inst_dmem_ram_3866), .A2(MEM_stage_inst_dmem_n20891), .ZN(MEM_stage_inst_dmem_n20872) );
NAND2_X1 MEM_stage_inst_dmem_U20631 ( .A1(MEM_stage_inst_dmem_n20870), .A2(MEM_stage_inst_dmem_n20869), .ZN(MEM_stage_inst_dmem_n9046) );
NAND2_X1 MEM_stage_inst_dmem_U20630 ( .A1(MEM_stage_inst_dmem_n14705), .A2(MEM_stage_inst_dmem_n20892), .ZN(MEM_stage_inst_dmem_n20869) );
NAND2_X1 MEM_stage_inst_dmem_U20629 ( .A1(MEM_stage_inst_dmem_ram_3867), .A2(MEM_stage_inst_dmem_n20891), .ZN(MEM_stage_inst_dmem_n20870) );
NAND2_X1 MEM_stage_inst_dmem_U20628 ( .A1(MEM_stage_inst_dmem_n20868), .A2(MEM_stage_inst_dmem_n20867), .ZN(MEM_stage_inst_dmem_n9047) );
NAND2_X1 MEM_stage_inst_dmem_U20627 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n20892), .ZN(MEM_stage_inst_dmem_n20867) );
NAND2_X1 MEM_stage_inst_dmem_U20626 ( .A1(MEM_stage_inst_dmem_ram_3868), .A2(MEM_stage_inst_dmem_n20891), .ZN(MEM_stage_inst_dmem_n20868) );
NAND2_X1 MEM_stage_inst_dmem_U20625 ( .A1(MEM_stage_inst_dmem_n20866), .A2(MEM_stage_inst_dmem_n20865), .ZN(MEM_stage_inst_dmem_n9048) );
NAND2_X1 MEM_stage_inst_dmem_U20624 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n20892), .ZN(MEM_stage_inst_dmem_n20865) );
NAND2_X1 MEM_stage_inst_dmem_U20623 ( .A1(MEM_stage_inst_dmem_ram_3869), .A2(MEM_stage_inst_dmem_n20891), .ZN(MEM_stage_inst_dmem_n20866) );
NAND2_X1 MEM_stage_inst_dmem_U20622 ( .A1(MEM_stage_inst_dmem_n20864), .A2(MEM_stage_inst_dmem_n20863), .ZN(MEM_stage_inst_dmem_n9049) );
NAND2_X1 MEM_stage_inst_dmem_U20621 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n20892), .ZN(MEM_stage_inst_dmem_n20863) );
NAND2_X1 MEM_stage_inst_dmem_U20620 ( .A1(MEM_stage_inst_dmem_ram_3870), .A2(MEM_stage_inst_dmem_n20891), .ZN(MEM_stage_inst_dmem_n20864) );
NAND2_X1 MEM_stage_inst_dmem_U20619 ( .A1(MEM_stage_inst_dmem_n20862), .A2(MEM_stage_inst_dmem_n20861), .ZN(MEM_stage_inst_dmem_n9050) );
NAND2_X1 MEM_stage_inst_dmem_U20618 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n20892), .ZN(MEM_stage_inst_dmem_n20861) );
INV_X1 MEM_stage_inst_dmem_U20617 ( .A(MEM_stage_inst_dmem_n20891), .ZN(MEM_stage_inst_dmem_n20892) );
NAND2_X1 MEM_stage_inst_dmem_U20616 ( .A1(MEM_stage_inst_dmem_ram_3871), .A2(MEM_stage_inst_dmem_n20891), .ZN(MEM_stage_inst_dmem_n20862) );
NAND2_X1 MEM_stage_inst_dmem_U20615 ( .A1(MEM_stage_inst_dmem_n21429), .A2(MEM_stage_inst_dmem_n20895), .ZN(MEM_stage_inst_dmem_n20891) );
NAND2_X1 MEM_stage_inst_dmem_U20614 ( .A1(MEM_stage_inst_dmem_n20860), .A2(MEM_stage_inst_dmem_n20859), .ZN(MEM_stage_inst_dmem_n9051) );
NAND2_X1 MEM_stage_inst_dmem_U20613 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n20858), .ZN(MEM_stage_inst_dmem_n20859) );
NAND2_X1 MEM_stage_inst_dmem_U20612 ( .A1(MEM_stage_inst_dmem_ram_3872), .A2(MEM_stage_inst_dmem_n20857), .ZN(MEM_stage_inst_dmem_n20860) );
NAND2_X1 MEM_stage_inst_dmem_U20611 ( .A1(MEM_stage_inst_dmem_n20856), .A2(MEM_stage_inst_dmem_n20855), .ZN(MEM_stage_inst_dmem_n9052) );
NAND2_X1 MEM_stage_inst_dmem_U20610 ( .A1(MEM_stage_inst_dmem_n109), .A2(MEM_stage_inst_dmem_n20858), .ZN(MEM_stage_inst_dmem_n20855) );
NAND2_X1 MEM_stage_inst_dmem_U20609 ( .A1(MEM_stage_inst_dmem_ram_3873), .A2(MEM_stage_inst_dmem_n20857), .ZN(MEM_stage_inst_dmem_n20856) );
NAND2_X1 MEM_stage_inst_dmem_U20608 ( .A1(MEM_stage_inst_dmem_n20854), .A2(MEM_stage_inst_dmem_n20853), .ZN(MEM_stage_inst_dmem_n9053) );
NAND2_X1 MEM_stage_inst_dmem_U20607 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n20858), .ZN(MEM_stage_inst_dmem_n20853) );
NAND2_X1 MEM_stage_inst_dmem_U20606 ( .A1(MEM_stage_inst_dmem_ram_3874), .A2(MEM_stage_inst_dmem_n20857), .ZN(MEM_stage_inst_dmem_n20854) );
NAND2_X1 MEM_stage_inst_dmem_U20605 ( .A1(MEM_stage_inst_dmem_n20852), .A2(MEM_stage_inst_dmem_n20851), .ZN(MEM_stage_inst_dmem_n9054) );
NAND2_X1 MEM_stage_inst_dmem_U20604 ( .A1(MEM_stage_inst_dmem_n13064), .A2(MEM_stage_inst_dmem_n20858), .ZN(MEM_stage_inst_dmem_n20851) );
NAND2_X1 MEM_stage_inst_dmem_U20603 ( .A1(MEM_stage_inst_dmem_ram_3875), .A2(MEM_stage_inst_dmem_n20857), .ZN(MEM_stage_inst_dmem_n20852) );
NAND2_X1 MEM_stage_inst_dmem_U20602 ( .A1(MEM_stage_inst_dmem_n20850), .A2(MEM_stage_inst_dmem_n20849), .ZN(MEM_stage_inst_dmem_n9055) );
NAND2_X1 MEM_stage_inst_dmem_U20601 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n20858), .ZN(MEM_stage_inst_dmem_n20849) );
NAND2_X1 MEM_stage_inst_dmem_U20600 ( .A1(MEM_stage_inst_dmem_ram_3876), .A2(MEM_stage_inst_dmem_n20857), .ZN(MEM_stage_inst_dmem_n20850) );
NAND2_X1 MEM_stage_inst_dmem_U20599 ( .A1(MEM_stage_inst_dmem_n20848), .A2(MEM_stage_inst_dmem_n20847), .ZN(MEM_stage_inst_dmem_n9056) );
NAND2_X1 MEM_stage_inst_dmem_U20598 ( .A1(MEM_stage_inst_dmem_n13059), .A2(MEM_stage_inst_dmem_n20858), .ZN(MEM_stage_inst_dmem_n20847) );
NAND2_X1 MEM_stage_inst_dmem_U20597 ( .A1(MEM_stage_inst_dmem_ram_3877), .A2(MEM_stage_inst_dmem_n20857), .ZN(MEM_stage_inst_dmem_n20848) );
NAND2_X1 MEM_stage_inst_dmem_U20596 ( .A1(MEM_stage_inst_dmem_n20846), .A2(MEM_stage_inst_dmem_n20845), .ZN(MEM_stage_inst_dmem_n9057) );
NAND2_X1 MEM_stage_inst_dmem_U20595 ( .A1(MEM_stage_inst_dmem_n13056), .A2(MEM_stage_inst_dmem_n20858), .ZN(MEM_stage_inst_dmem_n20845) );
NAND2_X1 MEM_stage_inst_dmem_U20594 ( .A1(MEM_stage_inst_dmem_ram_3878), .A2(MEM_stage_inst_dmem_n20857), .ZN(MEM_stage_inst_dmem_n20846) );
NAND2_X1 MEM_stage_inst_dmem_U20593 ( .A1(MEM_stage_inst_dmem_n20844), .A2(MEM_stage_inst_dmem_n20843), .ZN(MEM_stage_inst_dmem_n9058) );
NAND2_X1 MEM_stage_inst_dmem_U20592 ( .A1(MEM_stage_inst_dmem_n13886), .A2(MEM_stage_inst_dmem_n20858), .ZN(MEM_stage_inst_dmem_n20843) );
NAND2_X1 MEM_stage_inst_dmem_U20591 ( .A1(MEM_stage_inst_dmem_ram_3879), .A2(MEM_stage_inst_dmem_n20857), .ZN(MEM_stage_inst_dmem_n20844) );
NAND2_X1 MEM_stage_inst_dmem_U20590 ( .A1(MEM_stage_inst_dmem_n20842), .A2(MEM_stage_inst_dmem_n20841), .ZN(MEM_stage_inst_dmem_n9059) );
NAND2_X1 MEM_stage_inst_dmem_U20589 ( .A1(MEM_stage_inst_dmem_n21335), .A2(MEM_stage_inst_dmem_n20858), .ZN(MEM_stage_inst_dmem_n20841) );
NAND2_X1 MEM_stage_inst_dmem_U20588 ( .A1(MEM_stage_inst_dmem_ram_3880), .A2(MEM_stage_inst_dmem_n20857), .ZN(MEM_stage_inst_dmem_n20842) );
NAND2_X1 MEM_stage_inst_dmem_U20587 ( .A1(MEM_stage_inst_dmem_n20840), .A2(MEM_stage_inst_dmem_n20839), .ZN(MEM_stage_inst_dmem_n9060) );
NAND2_X1 MEM_stage_inst_dmem_U20586 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n20858), .ZN(MEM_stage_inst_dmem_n20839) );
NAND2_X1 MEM_stage_inst_dmem_U20585 ( .A1(MEM_stage_inst_dmem_ram_3881), .A2(MEM_stage_inst_dmem_n20857), .ZN(MEM_stage_inst_dmem_n20840) );
NAND2_X1 MEM_stage_inst_dmem_U20584 ( .A1(MEM_stage_inst_dmem_n20838), .A2(MEM_stage_inst_dmem_n20837), .ZN(MEM_stage_inst_dmem_n9061) );
NAND2_X1 MEM_stage_inst_dmem_U20583 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n20858), .ZN(MEM_stage_inst_dmem_n20837) );
NAND2_X1 MEM_stage_inst_dmem_U20582 ( .A1(MEM_stage_inst_dmem_ram_3882), .A2(MEM_stage_inst_dmem_n20857), .ZN(MEM_stage_inst_dmem_n20838) );
NAND2_X1 MEM_stage_inst_dmem_U20581 ( .A1(MEM_stage_inst_dmem_n20836), .A2(MEM_stage_inst_dmem_n20835), .ZN(MEM_stage_inst_dmem_n9062) );
NAND2_X1 MEM_stage_inst_dmem_U20580 ( .A1(MEM_stage_inst_dmem_n20904), .A2(MEM_stage_inst_dmem_n20858), .ZN(MEM_stage_inst_dmem_n20835) );
NAND2_X1 MEM_stage_inst_dmem_U20579 ( .A1(MEM_stage_inst_dmem_ram_3883), .A2(MEM_stage_inst_dmem_n20857), .ZN(MEM_stage_inst_dmem_n20836) );
NAND2_X1 MEM_stage_inst_dmem_U20578 ( .A1(MEM_stage_inst_dmem_n20834), .A2(MEM_stage_inst_dmem_n20833), .ZN(MEM_stage_inst_dmem_n9063) );
NAND2_X1 MEM_stage_inst_dmem_U20577 ( .A1(MEM_stage_inst_dmem_n13041), .A2(MEM_stage_inst_dmem_n20858), .ZN(MEM_stage_inst_dmem_n20833) );
NAND2_X1 MEM_stage_inst_dmem_U20576 ( .A1(MEM_stage_inst_dmem_ram_3884), .A2(MEM_stage_inst_dmem_n20857), .ZN(MEM_stage_inst_dmem_n20834) );
NAND2_X1 MEM_stage_inst_dmem_U20575 ( .A1(MEM_stage_inst_dmem_n20832), .A2(MEM_stage_inst_dmem_n20831), .ZN(MEM_stage_inst_dmem_n9064) );
NAND2_X1 MEM_stage_inst_dmem_U20574 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n20858), .ZN(MEM_stage_inst_dmem_n20831) );
NAND2_X1 MEM_stage_inst_dmem_U20573 ( .A1(MEM_stage_inst_dmem_ram_3885), .A2(MEM_stage_inst_dmem_n20857), .ZN(MEM_stage_inst_dmem_n20832) );
NAND2_X1 MEM_stage_inst_dmem_U20572 ( .A1(MEM_stage_inst_dmem_n20830), .A2(MEM_stage_inst_dmem_n20829), .ZN(MEM_stage_inst_dmem_n9065) );
NAND2_X1 MEM_stage_inst_dmem_U20571 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n20858), .ZN(MEM_stage_inst_dmem_n20829) );
NAND2_X1 MEM_stage_inst_dmem_U20570 ( .A1(MEM_stage_inst_dmem_ram_3886), .A2(MEM_stage_inst_dmem_n20857), .ZN(MEM_stage_inst_dmem_n20830) );
NAND2_X1 MEM_stage_inst_dmem_U20569 ( .A1(MEM_stage_inst_dmem_n20828), .A2(MEM_stage_inst_dmem_n20827), .ZN(MEM_stage_inst_dmem_n9066) );
NAND2_X1 MEM_stage_inst_dmem_U20568 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n20858), .ZN(MEM_stage_inst_dmem_n20827) );
NAND2_X1 MEM_stage_inst_dmem_U20567 ( .A1(MEM_stage_inst_dmem_ram_3887), .A2(MEM_stage_inst_dmem_n20857), .ZN(MEM_stage_inst_dmem_n20828) );
NAND2_X1 MEM_stage_inst_dmem_U20566 ( .A1(MEM_stage_inst_dmem_n21394), .A2(MEM_stage_inst_dmem_n20895), .ZN(MEM_stage_inst_dmem_n20857) );
NAND2_X1 MEM_stage_inst_dmem_U20565 ( .A1(MEM_stage_inst_dmem_n20826), .A2(MEM_stage_inst_dmem_n20825), .ZN(MEM_stage_inst_dmem_n9067) );
NAND2_X1 MEM_stage_inst_dmem_U20564 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n20824), .ZN(MEM_stage_inst_dmem_n20825) );
NAND2_X1 MEM_stage_inst_dmem_U20563 ( .A1(MEM_stage_inst_dmem_ram_3888), .A2(MEM_stage_inst_dmem_n20823), .ZN(MEM_stage_inst_dmem_n20826) );
NAND2_X1 MEM_stage_inst_dmem_U20562 ( .A1(MEM_stage_inst_dmem_n20822), .A2(MEM_stage_inst_dmem_n20821), .ZN(MEM_stage_inst_dmem_n9068) );
NAND2_X1 MEM_stage_inst_dmem_U20561 ( .A1(MEM_stage_inst_dmem_n109), .A2(MEM_stage_inst_dmem_n20824), .ZN(MEM_stage_inst_dmem_n20821) );
NAND2_X1 MEM_stage_inst_dmem_U20560 ( .A1(MEM_stage_inst_dmem_ram_3889), .A2(MEM_stage_inst_dmem_n20823), .ZN(MEM_stage_inst_dmem_n20822) );
NAND2_X1 MEM_stage_inst_dmem_U20559 ( .A1(MEM_stage_inst_dmem_n20820), .A2(MEM_stage_inst_dmem_n20819), .ZN(MEM_stage_inst_dmem_n9069) );
NAND2_X1 MEM_stage_inst_dmem_U20558 ( .A1(MEM_stage_inst_dmem_n16789), .A2(MEM_stage_inst_dmem_n20824), .ZN(MEM_stage_inst_dmem_n20819) );
NAND2_X1 MEM_stage_inst_dmem_U20557 ( .A1(MEM_stage_inst_dmem_ram_3890), .A2(MEM_stage_inst_dmem_n20823), .ZN(MEM_stage_inst_dmem_n20820) );
NAND2_X1 MEM_stage_inst_dmem_U20556 ( .A1(MEM_stage_inst_dmem_n20818), .A2(MEM_stage_inst_dmem_n20817), .ZN(MEM_stage_inst_dmem_n9070) );
NAND2_X1 MEM_stage_inst_dmem_U20555 ( .A1(MEM_stage_inst_dmem_n13064), .A2(MEM_stage_inst_dmem_n20824), .ZN(MEM_stage_inst_dmem_n20817) );
NAND2_X1 MEM_stage_inst_dmem_U20554 ( .A1(MEM_stage_inst_dmem_ram_3891), .A2(MEM_stage_inst_dmem_n20823), .ZN(MEM_stage_inst_dmem_n20818) );
NAND2_X1 MEM_stage_inst_dmem_U20553 ( .A1(MEM_stage_inst_dmem_n20816), .A2(MEM_stage_inst_dmem_n20815), .ZN(MEM_stage_inst_dmem_n9071) );
NAND2_X1 MEM_stage_inst_dmem_U20552 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n20824), .ZN(MEM_stage_inst_dmem_n20815) );
NAND2_X1 MEM_stage_inst_dmem_U20551 ( .A1(MEM_stage_inst_dmem_ram_3892), .A2(MEM_stage_inst_dmem_n20823), .ZN(MEM_stage_inst_dmem_n20816) );
NAND2_X1 MEM_stage_inst_dmem_U20550 ( .A1(MEM_stage_inst_dmem_n20814), .A2(MEM_stage_inst_dmem_n20813), .ZN(MEM_stage_inst_dmem_n9072) );
NAND2_X1 MEM_stage_inst_dmem_U20549 ( .A1(MEM_stage_inst_dmem_n13059), .A2(MEM_stage_inst_dmem_n20824), .ZN(MEM_stage_inst_dmem_n20813) );
NAND2_X1 MEM_stage_inst_dmem_U20548 ( .A1(MEM_stage_inst_dmem_ram_3893), .A2(MEM_stage_inst_dmem_n20823), .ZN(MEM_stage_inst_dmem_n20814) );
NAND2_X1 MEM_stage_inst_dmem_U20547 ( .A1(MEM_stage_inst_dmem_n20812), .A2(MEM_stage_inst_dmem_n20811), .ZN(MEM_stage_inst_dmem_n9073) );
NAND2_X1 MEM_stage_inst_dmem_U20546 ( .A1(MEM_stage_inst_dmem_n13056), .A2(MEM_stage_inst_dmem_n20824), .ZN(MEM_stage_inst_dmem_n20811) );
NAND2_X1 MEM_stage_inst_dmem_U20545 ( .A1(MEM_stage_inst_dmem_ram_3894), .A2(MEM_stage_inst_dmem_n20823), .ZN(MEM_stage_inst_dmem_n20812) );
NAND2_X1 MEM_stage_inst_dmem_U20544 ( .A1(MEM_stage_inst_dmem_n20810), .A2(MEM_stage_inst_dmem_n20809), .ZN(MEM_stage_inst_dmem_n9074) );
NAND2_X1 MEM_stage_inst_dmem_U20543 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n20824), .ZN(MEM_stage_inst_dmem_n20809) );
NAND2_X1 MEM_stage_inst_dmem_U20542 ( .A1(MEM_stage_inst_dmem_ram_3895), .A2(MEM_stage_inst_dmem_n20823), .ZN(MEM_stage_inst_dmem_n20810) );
NAND2_X1 MEM_stage_inst_dmem_U20541 ( .A1(MEM_stage_inst_dmem_n20808), .A2(MEM_stage_inst_dmem_n20807), .ZN(MEM_stage_inst_dmem_n9075) );
NAND2_X1 MEM_stage_inst_dmem_U20540 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n20824), .ZN(MEM_stage_inst_dmem_n20807) );
NAND2_X1 MEM_stage_inst_dmem_U20539 ( .A1(MEM_stage_inst_dmem_ram_3896), .A2(MEM_stage_inst_dmem_n20823), .ZN(MEM_stage_inst_dmem_n20808) );
NAND2_X1 MEM_stage_inst_dmem_U20538 ( .A1(MEM_stage_inst_dmem_n20806), .A2(MEM_stage_inst_dmem_n20805), .ZN(MEM_stage_inst_dmem_n9076) );
NAND2_X1 MEM_stage_inst_dmem_U20537 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n20824), .ZN(MEM_stage_inst_dmem_n20805) );
NAND2_X1 MEM_stage_inst_dmem_U20536 ( .A1(MEM_stage_inst_dmem_ram_3897), .A2(MEM_stage_inst_dmem_n20823), .ZN(MEM_stage_inst_dmem_n20806) );
NAND2_X1 MEM_stage_inst_dmem_U20535 ( .A1(MEM_stage_inst_dmem_n20804), .A2(MEM_stage_inst_dmem_n20803), .ZN(MEM_stage_inst_dmem_n9077) );
NAND2_X1 MEM_stage_inst_dmem_U20534 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n20824), .ZN(MEM_stage_inst_dmem_n20803) );
NAND2_X1 MEM_stage_inst_dmem_U20533 ( .A1(MEM_stage_inst_dmem_ram_3898), .A2(MEM_stage_inst_dmem_n20823), .ZN(MEM_stage_inst_dmem_n20804) );
NAND2_X1 MEM_stage_inst_dmem_U20532 ( .A1(MEM_stage_inst_dmem_n20802), .A2(MEM_stage_inst_dmem_n20801), .ZN(MEM_stage_inst_dmem_n9078) );
NAND2_X1 MEM_stage_inst_dmem_U20531 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n20824), .ZN(MEM_stage_inst_dmem_n20801) );
NAND2_X1 MEM_stage_inst_dmem_U20530 ( .A1(MEM_stage_inst_dmem_ram_3899), .A2(MEM_stage_inst_dmem_n20823), .ZN(MEM_stage_inst_dmem_n20802) );
NAND2_X1 MEM_stage_inst_dmem_U20529 ( .A1(MEM_stage_inst_dmem_n20800), .A2(MEM_stage_inst_dmem_n20799), .ZN(MEM_stage_inst_dmem_n9079) );
NAND2_X1 MEM_stage_inst_dmem_U20528 ( .A1(MEM_stage_inst_dmem_n18001), .A2(MEM_stage_inst_dmem_n20824), .ZN(MEM_stage_inst_dmem_n20799) );
NAND2_X1 MEM_stage_inst_dmem_U20527 ( .A1(MEM_stage_inst_dmem_ram_3900), .A2(MEM_stage_inst_dmem_n20823), .ZN(MEM_stage_inst_dmem_n20800) );
NAND2_X1 MEM_stage_inst_dmem_U20526 ( .A1(MEM_stage_inst_dmem_n20798), .A2(MEM_stage_inst_dmem_n20797), .ZN(MEM_stage_inst_dmem_n9080) );
NAND2_X1 MEM_stage_inst_dmem_U20525 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n20824), .ZN(MEM_stage_inst_dmem_n20797) );
NAND2_X1 MEM_stage_inst_dmem_U20524 ( .A1(MEM_stage_inst_dmem_ram_3901), .A2(MEM_stage_inst_dmem_n20823), .ZN(MEM_stage_inst_dmem_n20798) );
NAND2_X1 MEM_stage_inst_dmem_U20523 ( .A1(MEM_stage_inst_dmem_n20796), .A2(MEM_stage_inst_dmem_n20795), .ZN(MEM_stage_inst_dmem_n9081) );
NAND2_X1 MEM_stage_inst_dmem_U20522 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n20824), .ZN(MEM_stage_inst_dmem_n20795) );
NAND2_X1 MEM_stage_inst_dmem_U20521 ( .A1(MEM_stage_inst_dmem_ram_3902), .A2(MEM_stage_inst_dmem_n20823), .ZN(MEM_stage_inst_dmem_n20796) );
NAND2_X1 MEM_stage_inst_dmem_U20520 ( .A1(MEM_stage_inst_dmem_n20794), .A2(MEM_stage_inst_dmem_n20793), .ZN(MEM_stage_inst_dmem_n9082) );
NAND2_X1 MEM_stage_inst_dmem_U20519 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n20824), .ZN(MEM_stage_inst_dmem_n20793) );
INV_X1 MEM_stage_inst_dmem_U20518 ( .A(MEM_stage_inst_dmem_n20823), .ZN(MEM_stage_inst_dmem_n20824) );
NAND2_X1 MEM_stage_inst_dmem_U20517 ( .A1(MEM_stage_inst_dmem_ram_3903), .A2(MEM_stage_inst_dmem_n20823), .ZN(MEM_stage_inst_dmem_n20794) );
NAND2_X1 MEM_stage_inst_dmem_U20516 ( .A1(MEM_stage_inst_dmem_n21359), .A2(MEM_stage_inst_dmem_n20895), .ZN(MEM_stage_inst_dmem_n20823) );
NAND2_X1 MEM_stage_inst_dmem_U20515 ( .A1(MEM_stage_inst_dmem_n20792), .A2(MEM_stage_inst_dmem_n20791), .ZN(MEM_stage_inst_dmem_n9083) );
NAND2_X1 MEM_stage_inst_dmem_U20514 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n20790), .ZN(MEM_stage_inst_dmem_n20791) );
NAND2_X1 MEM_stage_inst_dmem_U20513 ( .A1(MEM_stage_inst_dmem_ram_3904), .A2(MEM_stage_inst_dmem_n20789), .ZN(MEM_stage_inst_dmem_n20792) );
NAND2_X1 MEM_stage_inst_dmem_U20512 ( .A1(MEM_stage_inst_dmem_n20788), .A2(MEM_stage_inst_dmem_n20787), .ZN(MEM_stage_inst_dmem_n9084) );
NAND2_X1 MEM_stage_inst_dmem_U20511 ( .A1(MEM_stage_inst_dmem_n20547), .A2(MEM_stage_inst_dmem_n20790), .ZN(MEM_stage_inst_dmem_n20787) );
NAND2_X1 MEM_stage_inst_dmem_U20510 ( .A1(MEM_stage_inst_dmem_ram_3905), .A2(MEM_stage_inst_dmem_n20789), .ZN(MEM_stage_inst_dmem_n20788) );
NAND2_X1 MEM_stage_inst_dmem_U20509 ( .A1(MEM_stage_inst_dmem_n20786), .A2(MEM_stage_inst_dmem_n20785), .ZN(MEM_stage_inst_dmem_n9085) );
NAND2_X1 MEM_stage_inst_dmem_U20508 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n20790), .ZN(MEM_stage_inst_dmem_n20785) );
NAND2_X1 MEM_stage_inst_dmem_U20507 ( .A1(MEM_stage_inst_dmem_ram_3906), .A2(MEM_stage_inst_dmem_n20789), .ZN(MEM_stage_inst_dmem_n20786) );
NAND2_X1 MEM_stage_inst_dmem_U20506 ( .A1(MEM_stage_inst_dmem_n20784), .A2(MEM_stage_inst_dmem_n20783), .ZN(MEM_stage_inst_dmem_n9086) );
NAND2_X1 MEM_stage_inst_dmem_U20505 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n20790), .ZN(MEM_stage_inst_dmem_n20783) );
NAND2_X1 MEM_stage_inst_dmem_U20504 ( .A1(MEM_stage_inst_dmem_ram_3907), .A2(MEM_stage_inst_dmem_n20789), .ZN(MEM_stage_inst_dmem_n20784) );
NAND2_X1 MEM_stage_inst_dmem_U20503 ( .A1(MEM_stage_inst_dmem_n20782), .A2(MEM_stage_inst_dmem_n20781), .ZN(MEM_stage_inst_dmem_n9087) );
NAND2_X1 MEM_stage_inst_dmem_U20502 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n20790), .ZN(MEM_stage_inst_dmem_n20781) );
NAND2_X1 MEM_stage_inst_dmem_U20501 ( .A1(MEM_stage_inst_dmem_ram_3908), .A2(MEM_stage_inst_dmem_n20789), .ZN(MEM_stage_inst_dmem_n20782) );
NAND2_X1 MEM_stage_inst_dmem_U20500 ( .A1(MEM_stage_inst_dmem_n20780), .A2(MEM_stage_inst_dmem_n20779), .ZN(MEM_stage_inst_dmem_n9088) );
NAND2_X1 MEM_stage_inst_dmem_U20499 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n20790), .ZN(MEM_stage_inst_dmem_n20779) );
NAND2_X1 MEM_stage_inst_dmem_U20498 ( .A1(MEM_stage_inst_dmem_ram_3909), .A2(MEM_stage_inst_dmem_n20789), .ZN(MEM_stage_inst_dmem_n20780) );
NAND2_X1 MEM_stage_inst_dmem_U20497 ( .A1(MEM_stage_inst_dmem_n20778), .A2(MEM_stage_inst_dmem_n20777), .ZN(MEM_stage_inst_dmem_n9089) );
NAND2_X1 MEM_stage_inst_dmem_U20496 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n20790), .ZN(MEM_stage_inst_dmem_n20777) );
NAND2_X1 MEM_stage_inst_dmem_U20495 ( .A1(MEM_stage_inst_dmem_ram_3910), .A2(MEM_stage_inst_dmem_n20789), .ZN(MEM_stage_inst_dmem_n20778) );
NAND2_X1 MEM_stage_inst_dmem_U20494 ( .A1(MEM_stage_inst_dmem_n20776), .A2(MEM_stage_inst_dmem_n20775), .ZN(MEM_stage_inst_dmem_n9090) );
NAND2_X1 MEM_stage_inst_dmem_U20493 ( .A1(MEM_stage_inst_dmem_n16361), .A2(MEM_stage_inst_dmem_n20790), .ZN(MEM_stage_inst_dmem_n20775) );
NAND2_X1 MEM_stage_inst_dmem_U20492 ( .A1(MEM_stage_inst_dmem_ram_3911), .A2(MEM_stage_inst_dmem_n20789), .ZN(MEM_stage_inst_dmem_n20776) );
NAND2_X1 MEM_stage_inst_dmem_U20491 ( .A1(MEM_stage_inst_dmem_n20774), .A2(MEM_stage_inst_dmem_n20773), .ZN(MEM_stage_inst_dmem_n9091) );
NAND2_X1 MEM_stage_inst_dmem_U20490 ( .A1(MEM_stage_inst_dmem_n13051), .A2(MEM_stage_inst_dmem_n20790), .ZN(MEM_stage_inst_dmem_n20773) );
NAND2_X1 MEM_stage_inst_dmem_U20489 ( .A1(MEM_stage_inst_dmem_ram_3912), .A2(MEM_stage_inst_dmem_n20789), .ZN(MEM_stage_inst_dmem_n20774) );
NAND2_X1 MEM_stage_inst_dmem_U20488 ( .A1(MEM_stage_inst_dmem_n20772), .A2(MEM_stage_inst_dmem_n20771), .ZN(MEM_stage_inst_dmem_n9092) );
NAND2_X1 MEM_stage_inst_dmem_U20487 ( .A1(MEM_stage_inst_dmem_n20524), .A2(MEM_stage_inst_dmem_n20790), .ZN(MEM_stage_inst_dmem_n20771) );
NAND2_X1 MEM_stage_inst_dmem_U20486 ( .A1(MEM_stage_inst_dmem_ram_3913), .A2(MEM_stage_inst_dmem_n20789), .ZN(MEM_stage_inst_dmem_n20772) );
NAND2_X1 MEM_stage_inst_dmem_U20485 ( .A1(MEM_stage_inst_dmem_n20770), .A2(MEM_stage_inst_dmem_n20769), .ZN(MEM_stage_inst_dmem_n9093) );
NAND2_X1 MEM_stage_inst_dmem_U20484 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n20790), .ZN(MEM_stage_inst_dmem_n20769) );
NAND2_X1 MEM_stage_inst_dmem_U20483 ( .A1(MEM_stage_inst_dmem_ram_3914), .A2(MEM_stage_inst_dmem_n20789), .ZN(MEM_stage_inst_dmem_n20770) );
NAND2_X1 MEM_stage_inst_dmem_U20482 ( .A1(MEM_stage_inst_dmem_n20768), .A2(MEM_stage_inst_dmem_n20767), .ZN(MEM_stage_inst_dmem_n9094) );
NAND2_X1 MEM_stage_inst_dmem_U20481 ( .A1(MEM_stage_inst_dmem_n14705), .A2(MEM_stage_inst_dmem_n20790), .ZN(MEM_stage_inst_dmem_n20767) );
NAND2_X1 MEM_stage_inst_dmem_U20480 ( .A1(MEM_stage_inst_dmem_ram_3915), .A2(MEM_stage_inst_dmem_n20789), .ZN(MEM_stage_inst_dmem_n20768) );
NAND2_X1 MEM_stage_inst_dmem_U20479 ( .A1(MEM_stage_inst_dmem_n20766), .A2(MEM_stage_inst_dmem_n20765), .ZN(MEM_stage_inst_dmem_n9095) );
NAND2_X1 MEM_stage_inst_dmem_U20478 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n20790), .ZN(MEM_stage_inst_dmem_n20765) );
NAND2_X1 MEM_stage_inst_dmem_U20477 ( .A1(MEM_stage_inst_dmem_ram_3916), .A2(MEM_stage_inst_dmem_n20789), .ZN(MEM_stage_inst_dmem_n20766) );
NAND2_X1 MEM_stage_inst_dmem_U20476 ( .A1(MEM_stage_inst_dmem_n20764), .A2(MEM_stage_inst_dmem_n20763), .ZN(MEM_stage_inst_dmem_n9096) );
NAND2_X1 MEM_stage_inst_dmem_U20475 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n20790), .ZN(MEM_stage_inst_dmem_n20763) );
NAND2_X1 MEM_stage_inst_dmem_U20474 ( .A1(MEM_stage_inst_dmem_ram_3917), .A2(MEM_stage_inst_dmem_n20789), .ZN(MEM_stage_inst_dmem_n20764) );
NAND2_X1 MEM_stage_inst_dmem_U20473 ( .A1(MEM_stage_inst_dmem_n20762), .A2(MEM_stage_inst_dmem_n20761), .ZN(MEM_stage_inst_dmem_n9097) );
NAND2_X1 MEM_stage_inst_dmem_U20472 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n20790), .ZN(MEM_stage_inst_dmem_n20761) );
NAND2_X1 MEM_stage_inst_dmem_U20471 ( .A1(MEM_stage_inst_dmem_ram_3918), .A2(MEM_stage_inst_dmem_n20789), .ZN(MEM_stage_inst_dmem_n20762) );
NAND2_X1 MEM_stage_inst_dmem_U20470 ( .A1(MEM_stage_inst_dmem_n20760), .A2(MEM_stage_inst_dmem_n20759), .ZN(MEM_stage_inst_dmem_n9098) );
NAND2_X1 MEM_stage_inst_dmem_U20469 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n20790), .ZN(MEM_stage_inst_dmem_n20759) );
INV_X1 MEM_stage_inst_dmem_U20468 ( .A(MEM_stage_inst_dmem_n20789), .ZN(MEM_stage_inst_dmem_n20790) );
NAND2_X1 MEM_stage_inst_dmem_U20467 ( .A1(MEM_stage_inst_dmem_ram_3919), .A2(MEM_stage_inst_dmem_n20789), .ZN(MEM_stage_inst_dmem_n20760) );
NAND2_X1 MEM_stage_inst_dmem_U20466 ( .A1(MEM_stage_inst_dmem_n21319), .A2(MEM_stage_inst_dmem_n20895), .ZN(MEM_stage_inst_dmem_n20789) );
NAND2_X1 MEM_stage_inst_dmem_U20465 ( .A1(MEM_stage_inst_dmem_n20758), .A2(MEM_stage_inst_dmem_n20757), .ZN(MEM_stage_inst_dmem_n9099) );
NAND2_X1 MEM_stage_inst_dmem_U20464 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n20756), .ZN(MEM_stage_inst_dmem_n20757) );
NAND2_X1 MEM_stage_inst_dmem_U20463 ( .A1(MEM_stage_inst_dmem_ram_3920), .A2(MEM_stage_inst_dmem_n20755), .ZN(MEM_stage_inst_dmem_n20758) );
NAND2_X1 MEM_stage_inst_dmem_U20462 ( .A1(MEM_stage_inst_dmem_n20754), .A2(MEM_stage_inst_dmem_n20753), .ZN(MEM_stage_inst_dmem_n9100) );
NAND2_X1 MEM_stage_inst_dmem_U20461 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n20756), .ZN(MEM_stage_inst_dmem_n20753) );
NAND2_X1 MEM_stage_inst_dmem_U20460 ( .A1(MEM_stage_inst_dmem_ram_3921), .A2(MEM_stage_inst_dmem_n20755), .ZN(MEM_stage_inst_dmem_n20754) );
NAND2_X1 MEM_stage_inst_dmem_U20459 ( .A1(MEM_stage_inst_dmem_n20752), .A2(MEM_stage_inst_dmem_n20751), .ZN(MEM_stage_inst_dmem_n9101) );
NAND2_X1 MEM_stage_inst_dmem_U20458 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n20756), .ZN(MEM_stage_inst_dmem_n20751) );
NAND2_X1 MEM_stage_inst_dmem_U20457 ( .A1(MEM_stage_inst_dmem_ram_3922), .A2(MEM_stage_inst_dmem_n20755), .ZN(MEM_stage_inst_dmem_n20752) );
NAND2_X1 MEM_stage_inst_dmem_U20456 ( .A1(MEM_stage_inst_dmem_n20750), .A2(MEM_stage_inst_dmem_n20749), .ZN(MEM_stage_inst_dmem_n9102) );
NAND2_X1 MEM_stage_inst_dmem_U20455 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n20756), .ZN(MEM_stage_inst_dmem_n20749) );
NAND2_X1 MEM_stage_inst_dmem_U20454 ( .A1(MEM_stage_inst_dmem_ram_3923), .A2(MEM_stage_inst_dmem_n20755), .ZN(MEM_stage_inst_dmem_n20750) );
NAND2_X1 MEM_stage_inst_dmem_U20453 ( .A1(MEM_stage_inst_dmem_n20748), .A2(MEM_stage_inst_dmem_n20747), .ZN(MEM_stage_inst_dmem_n9103) );
NAND2_X1 MEM_stage_inst_dmem_U20452 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n20756), .ZN(MEM_stage_inst_dmem_n20747) );
NAND2_X1 MEM_stage_inst_dmem_U20451 ( .A1(MEM_stage_inst_dmem_ram_3924), .A2(MEM_stage_inst_dmem_n20755), .ZN(MEM_stage_inst_dmem_n20748) );
NAND2_X1 MEM_stage_inst_dmem_U20450 ( .A1(MEM_stage_inst_dmem_n20746), .A2(MEM_stage_inst_dmem_n20745), .ZN(MEM_stage_inst_dmem_n9104) );
NAND2_X1 MEM_stage_inst_dmem_U20449 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n20756), .ZN(MEM_stage_inst_dmem_n20745) );
NAND2_X1 MEM_stage_inst_dmem_U20448 ( .A1(MEM_stage_inst_dmem_ram_3925), .A2(MEM_stage_inst_dmem_n20755), .ZN(MEM_stage_inst_dmem_n20746) );
NAND2_X1 MEM_stage_inst_dmem_U20447 ( .A1(MEM_stage_inst_dmem_n20744), .A2(MEM_stage_inst_dmem_n20743), .ZN(MEM_stage_inst_dmem_n9105) );
NAND2_X1 MEM_stage_inst_dmem_U20446 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n20756), .ZN(MEM_stage_inst_dmem_n20743) );
NAND2_X1 MEM_stage_inst_dmem_U20445 ( .A1(MEM_stage_inst_dmem_ram_3926), .A2(MEM_stage_inst_dmem_n20755), .ZN(MEM_stage_inst_dmem_n20744) );
NAND2_X1 MEM_stage_inst_dmem_U20444 ( .A1(MEM_stage_inst_dmem_n20742), .A2(MEM_stage_inst_dmem_n20741), .ZN(MEM_stage_inst_dmem_n9106) );
NAND2_X1 MEM_stage_inst_dmem_U20443 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n20756), .ZN(MEM_stage_inst_dmem_n20741) );
NAND2_X1 MEM_stage_inst_dmem_U20442 ( .A1(MEM_stage_inst_dmem_ram_3927), .A2(MEM_stage_inst_dmem_n20755), .ZN(MEM_stage_inst_dmem_n20742) );
NAND2_X1 MEM_stage_inst_dmem_U20441 ( .A1(MEM_stage_inst_dmem_n20740), .A2(MEM_stage_inst_dmem_n20739), .ZN(MEM_stage_inst_dmem_n9107) );
NAND2_X1 MEM_stage_inst_dmem_U20440 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n20756), .ZN(MEM_stage_inst_dmem_n20739) );
NAND2_X1 MEM_stage_inst_dmem_U20439 ( .A1(MEM_stage_inst_dmem_ram_3928), .A2(MEM_stage_inst_dmem_n20755), .ZN(MEM_stage_inst_dmem_n20740) );
NAND2_X1 MEM_stage_inst_dmem_U20438 ( .A1(MEM_stage_inst_dmem_n20738), .A2(MEM_stage_inst_dmem_n20737), .ZN(MEM_stage_inst_dmem_n9108) );
NAND2_X1 MEM_stage_inst_dmem_U20437 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n20756), .ZN(MEM_stage_inst_dmem_n20737) );
NAND2_X1 MEM_stage_inst_dmem_U20436 ( .A1(MEM_stage_inst_dmem_ram_3929), .A2(MEM_stage_inst_dmem_n20755), .ZN(MEM_stage_inst_dmem_n20738) );
NAND2_X1 MEM_stage_inst_dmem_U20435 ( .A1(MEM_stage_inst_dmem_n20736), .A2(MEM_stage_inst_dmem_n20735), .ZN(MEM_stage_inst_dmem_n9109) );
NAND2_X1 MEM_stage_inst_dmem_U20434 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n20756), .ZN(MEM_stage_inst_dmem_n20735) );
NAND2_X1 MEM_stage_inst_dmem_U20433 ( .A1(MEM_stage_inst_dmem_ram_3930), .A2(MEM_stage_inst_dmem_n20755), .ZN(MEM_stage_inst_dmem_n20736) );
NAND2_X1 MEM_stage_inst_dmem_U20432 ( .A1(MEM_stage_inst_dmem_n20734), .A2(MEM_stage_inst_dmem_n20733), .ZN(MEM_stage_inst_dmem_n9110) );
NAND2_X1 MEM_stage_inst_dmem_U20431 ( .A1(MEM_stage_inst_dmem_n20904), .A2(MEM_stage_inst_dmem_n20756), .ZN(MEM_stage_inst_dmem_n20733) );
NAND2_X1 MEM_stage_inst_dmem_U20430 ( .A1(MEM_stage_inst_dmem_ram_3931), .A2(MEM_stage_inst_dmem_n20755), .ZN(MEM_stage_inst_dmem_n20734) );
NAND2_X1 MEM_stage_inst_dmem_U20429 ( .A1(MEM_stage_inst_dmem_n20732), .A2(MEM_stage_inst_dmem_n20731), .ZN(MEM_stage_inst_dmem_n9111) );
NAND2_X1 MEM_stage_inst_dmem_U20428 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n20756), .ZN(MEM_stage_inst_dmem_n20731) );
NAND2_X1 MEM_stage_inst_dmem_U20427 ( .A1(MEM_stage_inst_dmem_ram_3932), .A2(MEM_stage_inst_dmem_n20755), .ZN(MEM_stage_inst_dmem_n20732) );
NAND2_X1 MEM_stage_inst_dmem_U20426 ( .A1(MEM_stage_inst_dmem_n20730), .A2(MEM_stage_inst_dmem_n20729), .ZN(MEM_stage_inst_dmem_n9112) );
NAND2_X1 MEM_stage_inst_dmem_U20425 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n20756), .ZN(MEM_stage_inst_dmem_n20729) );
NAND2_X1 MEM_stage_inst_dmem_U20424 ( .A1(MEM_stage_inst_dmem_ram_3933), .A2(MEM_stage_inst_dmem_n20755), .ZN(MEM_stage_inst_dmem_n20730) );
NAND2_X1 MEM_stage_inst_dmem_U20423 ( .A1(MEM_stage_inst_dmem_n20728), .A2(MEM_stage_inst_dmem_n20727), .ZN(MEM_stage_inst_dmem_n9113) );
NAND2_X1 MEM_stage_inst_dmem_U20422 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n20756), .ZN(MEM_stage_inst_dmem_n20727) );
NAND2_X1 MEM_stage_inst_dmem_U20421 ( .A1(MEM_stage_inst_dmem_ram_3934), .A2(MEM_stage_inst_dmem_n20755), .ZN(MEM_stage_inst_dmem_n20728) );
NAND2_X1 MEM_stage_inst_dmem_U20420 ( .A1(MEM_stage_inst_dmem_n20726), .A2(MEM_stage_inst_dmem_n20725), .ZN(MEM_stage_inst_dmem_n9114) );
NAND2_X1 MEM_stage_inst_dmem_U20419 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n20756), .ZN(MEM_stage_inst_dmem_n20725) );
INV_X1 MEM_stage_inst_dmem_U20418 ( .A(MEM_stage_inst_dmem_n20755), .ZN(MEM_stage_inst_dmem_n20756) );
NAND2_X1 MEM_stage_inst_dmem_U20417 ( .A1(MEM_stage_inst_dmem_ram_3935), .A2(MEM_stage_inst_dmem_n20755), .ZN(MEM_stage_inst_dmem_n20726) );
NAND2_X1 MEM_stage_inst_dmem_U20416 ( .A1(MEM_stage_inst_dmem_n21284), .A2(MEM_stage_inst_dmem_n20895), .ZN(MEM_stage_inst_dmem_n20755) );
NAND2_X1 MEM_stage_inst_dmem_U20415 ( .A1(MEM_stage_inst_dmem_n20724), .A2(MEM_stage_inst_dmem_n20723), .ZN(MEM_stage_inst_dmem_n9115) );
NAND2_X1 MEM_stage_inst_dmem_U20414 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n20722), .ZN(MEM_stage_inst_dmem_n20723) );
NAND2_X1 MEM_stage_inst_dmem_U20413 ( .A1(MEM_stage_inst_dmem_ram_3936), .A2(MEM_stage_inst_dmem_n20721), .ZN(MEM_stage_inst_dmem_n20724) );
NAND2_X1 MEM_stage_inst_dmem_U20412 ( .A1(MEM_stage_inst_dmem_n20720), .A2(MEM_stage_inst_dmem_n20719), .ZN(MEM_stage_inst_dmem_n9116) );
NAND2_X1 MEM_stage_inst_dmem_U20411 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n20722), .ZN(MEM_stage_inst_dmem_n20719) );
NAND2_X1 MEM_stage_inst_dmem_U20410 ( .A1(MEM_stage_inst_dmem_ram_3937), .A2(MEM_stage_inst_dmem_n20721), .ZN(MEM_stage_inst_dmem_n20720) );
NAND2_X1 MEM_stage_inst_dmem_U20409 ( .A1(MEM_stage_inst_dmem_n20718), .A2(MEM_stage_inst_dmem_n20717), .ZN(MEM_stage_inst_dmem_n9117) );
NAND2_X1 MEM_stage_inst_dmem_U20408 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n20722), .ZN(MEM_stage_inst_dmem_n20717) );
NAND2_X1 MEM_stage_inst_dmem_U20407 ( .A1(MEM_stage_inst_dmem_ram_3938), .A2(MEM_stage_inst_dmem_n20721), .ZN(MEM_stage_inst_dmem_n20718) );
NAND2_X1 MEM_stage_inst_dmem_U20406 ( .A1(MEM_stage_inst_dmem_n20716), .A2(MEM_stage_inst_dmem_n20715), .ZN(MEM_stage_inst_dmem_n9118) );
NAND2_X1 MEM_stage_inst_dmem_U20405 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n20722), .ZN(MEM_stage_inst_dmem_n20715) );
NAND2_X1 MEM_stage_inst_dmem_U20404 ( .A1(MEM_stage_inst_dmem_ram_3939), .A2(MEM_stage_inst_dmem_n20721), .ZN(MEM_stage_inst_dmem_n20716) );
NAND2_X1 MEM_stage_inst_dmem_U20403 ( .A1(MEM_stage_inst_dmem_n20714), .A2(MEM_stage_inst_dmem_n20713), .ZN(MEM_stage_inst_dmem_n9119) );
NAND2_X1 MEM_stage_inst_dmem_U20402 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n20722), .ZN(MEM_stage_inst_dmem_n20713) );
NAND2_X1 MEM_stage_inst_dmem_U20401 ( .A1(MEM_stage_inst_dmem_ram_3940), .A2(MEM_stage_inst_dmem_n20721), .ZN(MEM_stage_inst_dmem_n20714) );
NAND2_X1 MEM_stage_inst_dmem_U20400 ( .A1(MEM_stage_inst_dmem_n20712), .A2(MEM_stage_inst_dmem_n20711), .ZN(MEM_stage_inst_dmem_n9120) );
NAND2_X1 MEM_stage_inst_dmem_U20399 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n20722), .ZN(MEM_stage_inst_dmem_n20711) );
NAND2_X1 MEM_stage_inst_dmem_U20398 ( .A1(MEM_stage_inst_dmem_ram_3941), .A2(MEM_stage_inst_dmem_n20721), .ZN(MEM_stage_inst_dmem_n20712) );
NAND2_X1 MEM_stage_inst_dmem_U20397 ( .A1(MEM_stage_inst_dmem_n20710), .A2(MEM_stage_inst_dmem_n20709), .ZN(MEM_stage_inst_dmem_n9121) );
NAND2_X1 MEM_stage_inst_dmem_U20396 ( .A1(MEM_stage_inst_dmem_n14717), .A2(MEM_stage_inst_dmem_n20722), .ZN(MEM_stage_inst_dmem_n20709) );
NAND2_X1 MEM_stage_inst_dmem_U20395 ( .A1(MEM_stage_inst_dmem_ram_3942), .A2(MEM_stage_inst_dmem_n20721), .ZN(MEM_stage_inst_dmem_n20710) );
NAND2_X1 MEM_stage_inst_dmem_U20394 ( .A1(MEM_stage_inst_dmem_n20708), .A2(MEM_stage_inst_dmem_n20707), .ZN(MEM_stage_inst_dmem_n9122) );
NAND2_X1 MEM_stage_inst_dmem_U20393 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n20722), .ZN(MEM_stage_inst_dmem_n20707) );
NAND2_X1 MEM_stage_inst_dmem_U20392 ( .A1(MEM_stage_inst_dmem_ram_3943), .A2(MEM_stage_inst_dmem_n20721), .ZN(MEM_stage_inst_dmem_n20708) );
NAND2_X1 MEM_stage_inst_dmem_U20391 ( .A1(MEM_stage_inst_dmem_n20706), .A2(MEM_stage_inst_dmem_n20705), .ZN(MEM_stage_inst_dmem_n9123) );
NAND2_X1 MEM_stage_inst_dmem_U20390 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n20722), .ZN(MEM_stage_inst_dmem_n20705) );
NAND2_X1 MEM_stage_inst_dmem_U20389 ( .A1(MEM_stage_inst_dmem_ram_3944), .A2(MEM_stage_inst_dmem_n20721), .ZN(MEM_stage_inst_dmem_n20706) );
NAND2_X1 MEM_stage_inst_dmem_U20388 ( .A1(MEM_stage_inst_dmem_n20704), .A2(MEM_stage_inst_dmem_n20703), .ZN(MEM_stage_inst_dmem_n9124) );
NAND2_X1 MEM_stage_inst_dmem_U20387 ( .A1(EX_pipeline_reg_out_14), .A2(MEM_stage_inst_dmem_n20722), .ZN(MEM_stage_inst_dmem_n20703) );
NAND2_X1 MEM_stage_inst_dmem_U20386 ( .A1(MEM_stage_inst_dmem_ram_3945), .A2(MEM_stage_inst_dmem_n20721), .ZN(MEM_stage_inst_dmem_n20704) );
NAND2_X1 MEM_stage_inst_dmem_U20385 ( .A1(MEM_stage_inst_dmem_n20702), .A2(MEM_stage_inst_dmem_n20701), .ZN(MEM_stage_inst_dmem_n9125) );
NAND2_X1 MEM_stage_inst_dmem_U20384 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n20722), .ZN(MEM_stage_inst_dmem_n20701) );
NAND2_X1 MEM_stage_inst_dmem_U20383 ( .A1(MEM_stage_inst_dmem_ram_3946), .A2(MEM_stage_inst_dmem_n20721), .ZN(MEM_stage_inst_dmem_n20702) );
NAND2_X1 MEM_stage_inst_dmem_U20382 ( .A1(MEM_stage_inst_dmem_n20700), .A2(MEM_stage_inst_dmem_n20699), .ZN(MEM_stage_inst_dmem_n9126) );
NAND2_X1 MEM_stage_inst_dmem_U20381 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n20722), .ZN(MEM_stage_inst_dmem_n20699) );
NAND2_X1 MEM_stage_inst_dmem_U20380 ( .A1(MEM_stage_inst_dmem_ram_3947), .A2(MEM_stage_inst_dmem_n20721), .ZN(MEM_stage_inst_dmem_n20700) );
NAND2_X1 MEM_stage_inst_dmem_U20379 ( .A1(MEM_stage_inst_dmem_n20698), .A2(MEM_stage_inst_dmem_n20697), .ZN(MEM_stage_inst_dmem_n9127) );
NAND2_X1 MEM_stage_inst_dmem_U20378 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n20722), .ZN(MEM_stage_inst_dmem_n20697) );
NAND2_X1 MEM_stage_inst_dmem_U20377 ( .A1(MEM_stage_inst_dmem_ram_3948), .A2(MEM_stage_inst_dmem_n20721), .ZN(MEM_stage_inst_dmem_n20698) );
NAND2_X1 MEM_stage_inst_dmem_U20376 ( .A1(MEM_stage_inst_dmem_n20696), .A2(MEM_stage_inst_dmem_n20695), .ZN(MEM_stage_inst_dmem_n9128) );
NAND2_X1 MEM_stage_inst_dmem_U20375 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n20722), .ZN(MEM_stage_inst_dmem_n20695) );
NAND2_X1 MEM_stage_inst_dmem_U20374 ( .A1(MEM_stage_inst_dmem_ram_3949), .A2(MEM_stage_inst_dmem_n20721), .ZN(MEM_stage_inst_dmem_n20696) );
NAND2_X1 MEM_stage_inst_dmem_U20373 ( .A1(MEM_stage_inst_dmem_n20694), .A2(MEM_stage_inst_dmem_n20693), .ZN(MEM_stage_inst_dmem_n9129) );
NAND2_X1 MEM_stage_inst_dmem_U20372 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n20722), .ZN(MEM_stage_inst_dmem_n20693) );
NAND2_X1 MEM_stage_inst_dmem_U20371 ( .A1(MEM_stage_inst_dmem_ram_3950), .A2(MEM_stage_inst_dmem_n20721), .ZN(MEM_stage_inst_dmem_n20694) );
NAND2_X1 MEM_stage_inst_dmem_U20370 ( .A1(MEM_stage_inst_dmem_n20692), .A2(MEM_stage_inst_dmem_n20691), .ZN(MEM_stage_inst_dmem_n9130) );
NAND2_X1 MEM_stage_inst_dmem_U20369 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n20722), .ZN(MEM_stage_inst_dmem_n20691) );
INV_X1 MEM_stage_inst_dmem_U20368 ( .A(MEM_stage_inst_dmem_n20721), .ZN(MEM_stage_inst_dmem_n20722) );
NAND2_X1 MEM_stage_inst_dmem_U20367 ( .A1(MEM_stage_inst_dmem_ram_3951), .A2(MEM_stage_inst_dmem_n20721), .ZN(MEM_stage_inst_dmem_n20692) );
NAND2_X1 MEM_stage_inst_dmem_U20366 ( .A1(MEM_stage_inst_dmem_n21249), .A2(MEM_stage_inst_dmem_n20895), .ZN(MEM_stage_inst_dmem_n20721) );
NAND2_X1 MEM_stage_inst_dmem_U20365 ( .A1(MEM_stage_inst_dmem_n20690), .A2(MEM_stage_inst_dmem_n20689), .ZN(MEM_stage_inst_dmem_n9131) );
NAND2_X1 MEM_stage_inst_dmem_U20364 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n20688), .ZN(MEM_stage_inst_dmem_n20689) );
NAND2_X1 MEM_stage_inst_dmem_U20363 ( .A1(MEM_stage_inst_dmem_ram_3952), .A2(MEM_stage_inst_dmem_n20687), .ZN(MEM_stage_inst_dmem_n20690) );
NAND2_X1 MEM_stage_inst_dmem_U20362 ( .A1(MEM_stage_inst_dmem_n20686), .A2(MEM_stage_inst_dmem_n20685), .ZN(MEM_stage_inst_dmem_n9132) );
NAND2_X1 MEM_stage_inst_dmem_U20361 ( .A1(MEM_stage_inst_dmem_n109), .A2(MEM_stage_inst_dmem_n20688), .ZN(MEM_stage_inst_dmem_n20685) );
NAND2_X1 MEM_stage_inst_dmem_U20360 ( .A1(MEM_stage_inst_dmem_ram_3953), .A2(MEM_stage_inst_dmem_n20687), .ZN(MEM_stage_inst_dmem_n20686) );
NAND2_X1 MEM_stage_inst_dmem_U20359 ( .A1(MEM_stage_inst_dmem_n20684), .A2(MEM_stage_inst_dmem_n20683), .ZN(MEM_stage_inst_dmem_n9133) );
NAND2_X1 MEM_stage_inst_dmem_U20358 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n20688), .ZN(MEM_stage_inst_dmem_n20683) );
NAND2_X1 MEM_stage_inst_dmem_U20357 ( .A1(MEM_stage_inst_dmem_ram_3954), .A2(MEM_stage_inst_dmem_n20687), .ZN(MEM_stage_inst_dmem_n20684) );
NAND2_X1 MEM_stage_inst_dmem_U20356 ( .A1(MEM_stage_inst_dmem_n20682), .A2(MEM_stage_inst_dmem_n20681), .ZN(MEM_stage_inst_dmem_n9134) );
NAND2_X1 MEM_stage_inst_dmem_U20355 ( .A1(MEM_stage_inst_dmem_n13064), .A2(MEM_stage_inst_dmem_n20688), .ZN(MEM_stage_inst_dmem_n20681) );
NAND2_X1 MEM_stage_inst_dmem_U20354 ( .A1(MEM_stage_inst_dmem_ram_3955), .A2(MEM_stage_inst_dmem_n20687), .ZN(MEM_stage_inst_dmem_n20682) );
NAND2_X1 MEM_stage_inst_dmem_U20353 ( .A1(MEM_stage_inst_dmem_n20680), .A2(MEM_stage_inst_dmem_n20679), .ZN(MEM_stage_inst_dmem_n9135) );
NAND2_X1 MEM_stage_inst_dmem_U20352 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n20688), .ZN(MEM_stage_inst_dmem_n20679) );
NAND2_X1 MEM_stage_inst_dmem_U20351 ( .A1(MEM_stage_inst_dmem_ram_3956), .A2(MEM_stage_inst_dmem_n20687), .ZN(MEM_stage_inst_dmem_n20680) );
NAND2_X1 MEM_stage_inst_dmem_U20350 ( .A1(MEM_stage_inst_dmem_n20678), .A2(MEM_stage_inst_dmem_n20677), .ZN(MEM_stage_inst_dmem_n9136) );
NAND2_X1 MEM_stage_inst_dmem_U20349 ( .A1(MEM_stage_inst_dmem_n13059), .A2(MEM_stage_inst_dmem_n20688), .ZN(MEM_stage_inst_dmem_n20677) );
NAND2_X1 MEM_stage_inst_dmem_U20348 ( .A1(MEM_stage_inst_dmem_ram_3957), .A2(MEM_stage_inst_dmem_n20687), .ZN(MEM_stage_inst_dmem_n20678) );
NAND2_X1 MEM_stage_inst_dmem_U20347 ( .A1(MEM_stage_inst_dmem_n20676), .A2(MEM_stage_inst_dmem_n20675), .ZN(MEM_stage_inst_dmem_n9137) );
NAND2_X1 MEM_stage_inst_dmem_U20346 ( .A1(MEM_stage_inst_dmem_n13056), .A2(MEM_stage_inst_dmem_n20688), .ZN(MEM_stage_inst_dmem_n20675) );
NAND2_X1 MEM_stage_inst_dmem_U20345 ( .A1(MEM_stage_inst_dmem_ram_3958), .A2(MEM_stage_inst_dmem_n20687), .ZN(MEM_stage_inst_dmem_n20676) );
NAND2_X1 MEM_stage_inst_dmem_U20344 ( .A1(MEM_stage_inst_dmem_n20674), .A2(MEM_stage_inst_dmem_n20673), .ZN(MEM_stage_inst_dmem_n9138) );
NAND2_X1 MEM_stage_inst_dmem_U20343 ( .A1(MEM_stage_inst_dmem_n18), .A2(MEM_stage_inst_dmem_n20688), .ZN(MEM_stage_inst_dmem_n20673) );
NAND2_X1 MEM_stage_inst_dmem_U20342 ( .A1(MEM_stage_inst_dmem_ram_3959), .A2(MEM_stage_inst_dmem_n20687), .ZN(MEM_stage_inst_dmem_n20674) );
NAND2_X1 MEM_stage_inst_dmem_U20341 ( .A1(MEM_stage_inst_dmem_n20672), .A2(MEM_stage_inst_dmem_n20671), .ZN(MEM_stage_inst_dmem_n9139) );
NAND2_X1 MEM_stage_inst_dmem_U20340 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n20688), .ZN(MEM_stage_inst_dmem_n20671) );
NAND2_X1 MEM_stage_inst_dmem_U20339 ( .A1(MEM_stage_inst_dmem_ram_3960), .A2(MEM_stage_inst_dmem_n20687), .ZN(MEM_stage_inst_dmem_n20672) );
NAND2_X1 MEM_stage_inst_dmem_U20338 ( .A1(MEM_stage_inst_dmem_n20670), .A2(MEM_stage_inst_dmem_n20669), .ZN(MEM_stage_inst_dmem_n9140) );
NAND2_X1 MEM_stage_inst_dmem_U20337 ( .A1(MEM_stage_inst_dmem_n20524), .A2(MEM_stage_inst_dmem_n20688), .ZN(MEM_stage_inst_dmem_n20669) );
NAND2_X1 MEM_stage_inst_dmem_U20336 ( .A1(MEM_stage_inst_dmem_ram_3961), .A2(MEM_stage_inst_dmem_n20687), .ZN(MEM_stage_inst_dmem_n20670) );
NAND2_X1 MEM_stage_inst_dmem_U20335 ( .A1(MEM_stage_inst_dmem_n20668), .A2(MEM_stage_inst_dmem_n20667), .ZN(MEM_stage_inst_dmem_n9141) );
NAND2_X1 MEM_stage_inst_dmem_U20334 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n20688), .ZN(MEM_stage_inst_dmem_n20667) );
NAND2_X1 MEM_stage_inst_dmem_U20333 ( .A1(MEM_stage_inst_dmem_ram_3962), .A2(MEM_stage_inst_dmem_n20687), .ZN(MEM_stage_inst_dmem_n20668) );
NAND2_X1 MEM_stage_inst_dmem_U20332 ( .A1(MEM_stage_inst_dmem_n20666), .A2(MEM_stage_inst_dmem_n20665), .ZN(MEM_stage_inst_dmem_n9142) );
NAND2_X1 MEM_stage_inst_dmem_U20331 ( .A1(MEM_stage_inst_dmem_n14705), .A2(MEM_stage_inst_dmem_n20688), .ZN(MEM_stage_inst_dmem_n20665) );
NAND2_X1 MEM_stage_inst_dmem_U20330 ( .A1(MEM_stage_inst_dmem_ram_3963), .A2(MEM_stage_inst_dmem_n20687), .ZN(MEM_stage_inst_dmem_n20666) );
NAND2_X1 MEM_stage_inst_dmem_U20329 ( .A1(MEM_stage_inst_dmem_n20664), .A2(MEM_stage_inst_dmem_n20663), .ZN(MEM_stage_inst_dmem_n9143) );
NAND2_X1 MEM_stage_inst_dmem_U20328 ( .A1(MEM_stage_inst_dmem_n13041), .A2(MEM_stage_inst_dmem_n20688), .ZN(MEM_stage_inst_dmem_n20663) );
NAND2_X1 MEM_stage_inst_dmem_U20327 ( .A1(MEM_stage_inst_dmem_ram_3964), .A2(MEM_stage_inst_dmem_n20687), .ZN(MEM_stage_inst_dmem_n20664) );
NAND2_X1 MEM_stage_inst_dmem_U20326 ( .A1(MEM_stage_inst_dmem_n20662), .A2(MEM_stage_inst_dmem_n20661), .ZN(MEM_stage_inst_dmem_n9144) );
NAND2_X1 MEM_stage_inst_dmem_U20325 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n20688), .ZN(MEM_stage_inst_dmem_n20661) );
NAND2_X1 MEM_stage_inst_dmem_U20324 ( .A1(MEM_stage_inst_dmem_ram_3965), .A2(MEM_stage_inst_dmem_n20687), .ZN(MEM_stage_inst_dmem_n20662) );
NAND2_X1 MEM_stage_inst_dmem_U20323 ( .A1(MEM_stage_inst_dmem_n20660), .A2(MEM_stage_inst_dmem_n20659), .ZN(MEM_stage_inst_dmem_n9145) );
NAND2_X1 MEM_stage_inst_dmem_U20322 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n20688), .ZN(MEM_stage_inst_dmem_n20659) );
NAND2_X1 MEM_stage_inst_dmem_U20321 ( .A1(MEM_stage_inst_dmem_ram_3966), .A2(MEM_stage_inst_dmem_n20687), .ZN(MEM_stage_inst_dmem_n20660) );
NAND2_X1 MEM_stage_inst_dmem_U20320 ( .A1(MEM_stage_inst_dmem_n20658), .A2(MEM_stage_inst_dmem_n20657), .ZN(MEM_stage_inst_dmem_n9146) );
NAND2_X1 MEM_stage_inst_dmem_U20319 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n20688), .ZN(MEM_stage_inst_dmem_n20657) );
INV_X1 MEM_stage_inst_dmem_U20318 ( .A(MEM_stage_inst_dmem_n20687), .ZN(MEM_stage_inst_dmem_n20688) );
NAND2_X1 MEM_stage_inst_dmem_U20317 ( .A1(MEM_stage_inst_dmem_ram_3967), .A2(MEM_stage_inst_dmem_n20687), .ZN(MEM_stage_inst_dmem_n20658) );
NAND2_X1 MEM_stage_inst_dmem_U20316 ( .A1(MEM_stage_inst_dmem_n21214), .A2(MEM_stage_inst_dmem_n20895), .ZN(MEM_stage_inst_dmem_n20687) );
NAND2_X1 MEM_stage_inst_dmem_U20315 ( .A1(MEM_stage_inst_dmem_n20656), .A2(MEM_stage_inst_dmem_n20655), .ZN(MEM_stage_inst_dmem_n9147) );
NAND2_X1 MEM_stage_inst_dmem_U20314 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n20654), .ZN(MEM_stage_inst_dmem_n20655) );
NAND2_X1 MEM_stage_inst_dmem_U20313 ( .A1(MEM_stage_inst_dmem_ram_3968), .A2(MEM_stage_inst_dmem_n20653), .ZN(MEM_stage_inst_dmem_n20656) );
NAND2_X1 MEM_stage_inst_dmem_U20312 ( .A1(MEM_stage_inst_dmem_n20652), .A2(MEM_stage_inst_dmem_n20651), .ZN(MEM_stage_inst_dmem_n9148) );
NAND2_X1 MEM_stage_inst_dmem_U20311 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n20654), .ZN(MEM_stage_inst_dmem_n20651) );
NAND2_X1 MEM_stage_inst_dmem_U20310 ( .A1(MEM_stage_inst_dmem_ram_3969), .A2(MEM_stage_inst_dmem_n20653), .ZN(MEM_stage_inst_dmem_n20652) );
NAND2_X1 MEM_stage_inst_dmem_U20309 ( .A1(MEM_stage_inst_dmem_n20650), .A2(MEM_stage_inst_dmem_n20649), .ZN(MEM_stage_inst_dmem_n9149) );
NAND2_X1 MEM_stage_inst_dmem_U20308 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n20654), .ZN(MEM_stage_inst_dmem_n20649) );
NAND2_X1 MEM_stage_inst_dmem_U20307 ( .A1(MEM_stage_inst_dmem_ram_3970), .A2(MEM_stage_inst_dmem_n20653), .ZN(MEM_stage_inst_dmem_n20650) );
NAND2_X1 MEM_stage_inst_dmem_U20306 ( .A1(MEM_stage_inst_dmem_n20648), .A2(MEM_stage_inst_dmem_n20647), .ZN(MEM_stage_inst_dmem_n9150) );
NAND2_X1 MEM_stage_inst_dmem_U20305 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n20654), .ZN(MEM_stage_inst_dmem_n20647) );
NAND2_X1 MEM_stage_inst_dmem_U20304 ( .A1(MEM_stage_inst_dmem_ram_3971), .A2(MEM_stage_inst_dmem_n20653), .ZN(MEM_stage_inst_dmem_n20648) );
NAND2_X1 MEM_stage_inst_dmem_U20303 ( .A1(MEM_stage_inst_dmem_n20646), .A2(MEM_stage_inst_dmem_n20645), .ZN(MEM_stage_inst_dmem_n9151) );
NAND2_X1 MEM_stage_inst_dmem_U20302 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n20654), .ZN(MEM_stage_inst_dmem_n20645) );
NAND2_X1 MEM_stage_inst_dmem_U20301 ( .A1(MEM_stage_inst_dmem_ram_3972), .A2(MEM_stage_inst_dmem_n20653), .ZN(MEM_stage_inst_dmem_n20646) );
NAND2_X1 MEM_stage_inst_dmem_U20300 ( .A1(MEM_stage_inst_dmem_n20644), .A2(MEM_stage_inst_dmem_n20643), .ZN(MEM_stage_inst_dmem_n9152) );
NAND2_X1 MEM_stage_inst_dmem_U20299 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n20654), .ZN(MEM_stage_inst_dmem_n20643) );
NAND2_X1 MEM_stage_inst_dmem_U20298 ( .A1(MEM_stage_inst_dmem_ram_3973), .A2(MEM_stage_inst_dmem_n20653), .ZN(MEM_stage_inst_dmem_n20644) );
NAND2_X1 MEM_stage_inst_dmem_U20297 ( .A1(MEM_stage_inst_dmem_n20642), .A2(MEM_stage_inst_dmem_n20641), .ZN(MEM_stage_inst_dmem_n9153) );
NAND2_X1 MEM_stage_inst_dmem_U20296 ( .A1(MEM_stage_inst_dmem_n14717), .A2(MEM_stage_inst_dmem_n20654), .ZN(MEM_stage_inst_dmem_n20641) );
NAND2_X1 MEM_stage_inst_dmem_U20295 ( .A1(MEM_stage_inst_dmem_ram_3974), .A2(MEM_stage_inst_dmem_n20653), .ZN(MEM_stage_inst_dmem_n20642) );
NAND2_X1 MEM_stage_inst_dmem_U20294 ( .A1(MEM_stage_inst_dmem_n20640), .A2(MEM_stage_inst_dmem_n20639), .ZN(MEM_stage_inst_dmem_n9154) );
NAND2_X1 MEM_stage_inst_dmem_U20293 ( .A1(EX_pipeline_reg_out_12), .A2(MEM_stage_inst_dmem_n20654), .ZN(MEM_stage_inst_dmem_n20639) );
NAND2_X1 MEM_stage_inst_dmem_U20292 ( .A1(MEM_stage_inst_dmem_ram_3975), .A2(MEM_stage_inst_dmem_n20653), .ZN(MEM_stage_inst_dmem_n20640) );
NAND2_X1 MEM_stage_inst_dmem_U20291 ( .A1(MEM_stage_inst_dmem_n20638), .A2(MEM_stage_inst_dmem_n20637), .ZN(MEM_stage_inst_dmem_n9155) );
NAND2_X1 MEM_stage_inst_dmem_U20290 ( .A1(MEM_stage_inst_dmem_n13051), .A2(MEM_stage_inst_dmem_n20654), .ZN(MEM_stage_inst_dmem_n20637) );
NAND2_X1 MEM_stage_inst_dmem_U20289 ( .A1(MEM_stage_inst_dmem_ram_3976), .A2(MEM_stage_inst_dmem_n20653), .ZN(MEM_stage_inst_dmem_n20638) );
NAND2_X1 MEM_stage_inst_dmem_U20288 ( .A1(MEM_stage_inst_dmem_n20636), .A2(MEM_stage_inst_dmem_n20635), .ZN(MEM_stage_inst_dmem_n9156) );
NAND2_X1 MEM_stage_inst_dmem_U20287 ( .A1(MEM_stage_inst_dmem_n19251), .A2(MEM_stage_inst_dmem_n20654), .ZN(MEM_stage_inst_dmem_n20635) );
NAND2_X1 MEM_stage_inst_dmem_U20286 ( .A1(MEM_stage_inst_dmem_ram_3977), .A2(MEM_stage_inst_dmem_n20653), .ZN(MEM_stage_inst_dmem_n20636) );
NAND2_X1 MEM_stage_inst_dmem_U20285 ( .A1(MEM_stage_inst_dmem_n20634), .A2(MEM_stage_inst_dmem_n20633), .ZN(MEM_stage_inst_dmem_n9157) );
NAND2_X1 MEM_stage_inst_dmem_U20284 ( .A1(MEM_stage_inst_dmem_n16769), .A2(MEM_stage_inst_dmem_n20654), .ZN(MEM_stage_inst_dmem_n20633) );
NAND2_X1 MEM_stage_inst_dmem_U20283 ( .A1(MEM_stage_inst_dmem_ram_3978), .A2(MEM_stage_inst_dmem_n20653), .ZN(MEM_stage_inst_dmem_n20634) );
NAND2_X1 MEM_stage_inst_dmem_U20282 ( .A1(MEM_stage_inst_dmem_n20632), .A2(MEM_stage_inst_dmem_n20631), .ZN(MEM_stage_inst_dmem_n9158) );
NAND2_X1 MEM_stage_inst_dmem_U20281 ( .A1(MEM_stage_inst_dmem_n20904), .A2(MEM_stage_inst_dmem_n20654), .ZN(MEM_stage_inst_dmem_n20631) );
NAND2_X1 MEM_stage_inst_dmem_U20280 ( .A1(MEM_stage_inst_dmem_ram_3979), .A2(MEM_stage_inst_dmem_n20653), .ZN(MEM_stage_inst_dmem_n20632) );
NAND2_X1 MEM_stage_inst_dmem_U20279 ( .A1(MEM_stage_inst_dmem_n20630), .A2(MEM_stage_inst_dmem_n20629), .ZN(MEM_stage_inst_dmem_n9159) );
NAND2_X1 MEM_stage_inst_dmem_U20278 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n20654), .ZN(MEM_stage_inst_dmem_n20629) );
NAND2_X1 MEM_stage_inst_dmem_U20277 ( .A1(MEM_stage_inst_dmem_ram_3980), .A2(MEM_stage_inst_dmem_n20653), .ZN(MEM_stage_inst_dmem_n20630) );
NAND2_X1 MEM_stage_inst_dmem_U20276 ( .A1(MEM_stage_inst_dmem_n20628), .A2(MEM_stage_inst_dmem_n20627), .ZN(MEM_stage_inst_dmem_n9160) );
NAND2_X1 MEM_stage_inst_dmem_U20275 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n20654), .ZN(MEM_stage_inst_dmem_n20627) );
NAND2_X1 MEM_stage_inst_dmem_U20274 ( .A1(MEM_stage_inst_dmem_ram_3981), .A2(MEM_stage_inst_dmem_n20653), .ZN(MEM_stage_inst_dmem_n20628) );
NAND2_X1 MEM_stage_inst_dmem_U20273 ( .A1(MEM_stage_inst_dmem_n20626), .A2(MEM_stage_inst_dmem_n20625), .ZN(MEM_stage_inst_dmem_n9161) );
NAND2_X1 MEM_stage_inst_dmem_U20272 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n20654), .ZN(MEM_stage_inst_dmem_n20625) );
NAND2_X1 MEM_stage_inst_dmem_U20271 ( .A1(MEM_stage_inst_dmem_ram_3982), .A2(MEM_stage_inst_dmem_n20653), .ZN(MEM_stage_inst_dmem_n20626) );
NAND2_X1 MEM_stage_inst_dmem_U20270 ( .A1(MEM_stage_inst_dmem_n20624), .A2(MEM_stage_inst_dmem_n20623), .ZN(MEM_stage_inst_dmem_n9162) );
NAND2_X1 MEM_stage_inst_dmem_U20269 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n20654), .ZN(MEM_stage_inst_dmem_n20623) );
INV_X1 MEM_stage_inst_dmem_U20268 ( .A(MEM_stage_inst_dmem_n20653), .ZN(MEM_stage_inst_dmem_n20654) );
NAND2_X1 MEM_stage_inst_dmem_U20267 ( .A1(MEM_stage_inst_dmem_ram_3983), .A2(MEM_stage_inst_dmem_n20653), .ZN(MEM_stage_inst_dmem_n20624) );
NAND2_X1 MEM_stage_inst_dmem_U20266 ( .A1(MEM_stage_inst_dmem_n21179), .A2(MEM_stage_inst_dmem_n20895), .ZN(MEM_stage_inst_dmem_n20653) );
NAND2_X1 MEM_stage_inst_dmem_U20265 ( .A1(MEM_stage_inst_dmem_n20622), .A2(MEM_stage_inst_dmem_n20621), .ZN(MEM_stage_inst_dmem_n9163) );
NAND2_X1 MEM_stage_inst_dmem_U20264 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n20620), .ZN(MEM_stage_inst_dmem_n20621) );
NAND2_X1 MEM_stage_inst_dmem_U20263 ( .A1(MEM_stage_inst_dmem_ram_3984), .A2(MEM_stage_inst_dmem_n20619), .ZN(MEM_stage_inst_dmem_n20622) );
NAND2_X1 MEM_stage_inst_dmem_U20262 ( .A1(MEM_stage_inst_dmem_n20618), .A2(MEM_stage_inst_dmem_n20617), .ZN(MEM_stage_inst_dmem_n9164) );
NAND2_X1 MEM_stage_inst_dmem_U20261 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n20620), .ZN(MEM_stage_inst_dmem_n20617) );
NAND2_X1 MEM_stage_inst_dmem_U20260 ( .A1(MEM_stage_inst_dmem_ram_3985), .A2(MEM_stage_inst_dmem_n20619), .ZN(MEM_stage_inst_dmem_n20618) );
NAND2_X1 MEM_stage_inst_dmem_U20259 ( .A1(MEM_stage_inst_dmem_n20616), .A2(MEM_stage_inst_dmem_n20615), .ZN(MEM_stage_inst_dmem_n9165) );
NAND2_X1 MEM_stage_inst_dmem_U20258 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n20620), .ZN(MEM_stage_inst_dmem_n20615) );
NAND2_X1 MEM_stage_inst_dmem_U20257 ( .A1(MEM_stage_inst_dmem_ram_3986), .A2(MEM_stage_inst_dmem_n20619), .ZN(MEM_stage_inst_dmem_n20616) );
NAND2_X1 MEM_stage_inst_dmem_U20256 ( .A1(MEM_stage_inst_dmem_n20614), .A2(MEM_stage_inst_dmem_n20613), .ZN(MEM_stage_inst_dmem_n9166) );
NAND2_X1 MEM_stage_inst_dmem_U20255 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n20620), .ZN(MEM_stage_inst_dmem_n20613) );
NAND2_X1 MEM_stage_inst_dmem_U20254 ( .A1(MEM_stage_inst_dmem_ram_3987), .A2(MEM_stage_inst_dmem_n20619), .ZN(MEM_stage_inst_dmem_n20614) );
NAND2_X1 MEM_stage_inst_dmem_U20253 ( .A1(MEM_stage_inst_dmem_n20612), .A2(MEM_stage_inst_dmem_n20611), .ZN(MEM_stage_inst_dmem_n9167) );
NAND2_X1 MEM_stage_inst_dmem_U20252 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n20620), .ZN(MEM_stage_inst_dmem_n20611) );
NAND2_X1 MEM_stage_inst_dmem_U20251 ( .A1(MEM_stage_inst_dmem_ram_3988), .A2(MEM_stage_inst_dmem_n20619), .ZN(MEM_stage_inst_dmem_n20612) );
NAND2_X1 MEM_stage_inst_dmem_U20250 ( .A1(MEM_stage_inst_dmem_n20610), .A2(MEM_stage_inst_dmem_n20609), .ZN(MEM_stage_inst_dmem_n9168) );
NAND2_X1 MEM_stage_inst_dmem_U20249 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n20620), .ZN(MEM_stage_inst_dmem_n20609) );
NAND2_X1 MEM_stage_inst_dmem_U20248 ( .A1(MEM_stage_inst_dmem_ram_3989), .A2(MEM_stage_inst_dmem_n20619), .ZN(MEM_stage_inst_dmem_n20610) );
NAND2_X1 MEM_stage_inst_dmem_U20247 ( .A1(MEM_stage_inst_dmem_n20608), .A2(MEM_stage_inst_dmem_n20607), .ZN(MEM_stage_inst_dmem_n9169) );
NAND2_X1 MEM_stage_inst_dmem_U20246 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n20620), .ZN(MEM_stage_inst_dmem_n20607) );
NAND2_X1 MEM_stage_inst_dmem_U20245 ( .A1(MEM_stage_inst_dmem_ram_3990), .A2(MEM_stage_inst_dmem_n20619), .ZN(MEM_stage_inst_dmem_n20608) );
NAND2_X1 MEM_stage_inst_dmem_U20244 ( .A1(MEM_stage_inst_dmem_n20606), .A2(MEM_stage_inst_dmem_n20605), .ZN(MEM_stage_inst_dmem_n9170) );
NAND2_X1 MEM_stage_inst_dmem_U20243 ( .A1(MEM_stage_inst_dmem_n112), .A2(MEM_stage_inst_dmem_n20620), .ZN(MEM_stage_inst_dmem_n20605) );
NAND2_X1 MEM_stage_inst_dmem_U20242 ( .A1(MEM_stage_inst_dmem_ram_3991), .A2(MEM_stage_inst_dmem_n20619), .ZN(MEM_stage_inst_dmem_n20606) );
NAND2_X1 MEM_stage_inst_dmem_U20241 ( .A1(MEM_stage_inst_dmem_n20604), .A2(MEM_stage_inst_dmem_n20603), .ZN(MEM_stage_inst_dmem_n9171) );
NAND2_X1 MEM_stage_inst_dmem_U20240 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n20620), .ZN(MEM_stage_inst_dmem_n20603) );
NAND2_X1 MEM_stage_inst_dmem_U20239 ( .A1(MEM_stage_inst_dmem_ram_3992), .A2(MEM_stage_inst_dmem_n20619), .ZN(MEM_stage_inst_dmem_n20604) );
NAND2_X1 MEM_stage_inst_dmem_U20238 ( .A1(MEM_stage_inst_dmem_n20602), .A2(MEM_stage_inst_dmem_n20601), .ZN(MEM_stage_inst_dmem_n9172) );
NAND2_X1 MEM_stage_inst_dmem_U20237 ( .A1(MEM_stage_inst_dmem_n96), .A2(MEM_stage_inst_dmem_n20620), .ZN(MEM_stage_inst_dmem_n20601) );
NAND2_X1 MEM_stage_inst_dmem_U20236 ( .A1(MEM_stage_inst_dmem_ram_3993), .A2(MEM_stage_inst_dmem_n20619), .ZN(MEM_stage_inst_dmem_n20602) );
NAND2_X1 MEM_stage_inst_dmem_U20235 ( .A1(MEM_stage_inst_dmem_n20600), .A2(MEM_stage_inst_dmem_n20599), .ZN(MEM_stage_inst_dmem_n9173) );
NAND2_X1 MEM_stage_inst_dmem_U20234 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n20620), .ZN(MEM_stage_inst_dmem_n20599) );
NAND2_X1 MEM_stage_inst_dmem_U20233 ( .A1(MEM_stage_inst_dmem_ram_3994), .A2(MEM_stage_inst_dmem_n20619), .ZN(MEM_stage_inst_dmem_n20600) );
NAND2_X1 MEM_stage_inst_dmem_U20232 ( .A1(MEM_stage_inst_dmem_n20598), .A2(MEM_stage_inst_dmem_n20597), .ZN(MEM_stage_inst_dmem_n9174) );
NAND2_X1 MEM_stage_inst_dmem_U20231 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n20620), .ZN(MEM_stage_inst_dmem_n20597) );
NAND2_X1 MEM_stage_inst_dmem_U20230 ( .A1(MEM_stage_inst_dmem_ram_3995), .A2(MEM_stage_inst_dmem_n20619), .ZN(MEM_stage_inst_dmem_n20598) );
NAND2_X1 MEM_stage_inst_dmem_U20229 ( .A1(MEM_stage_inst_dmem_n20596), .A2(MEM_stage_inst_dmem_n20595), .ZN(MEM_stage_inst_dmem_n9175) );
NAND2_X1 MEM_stage_inst_dmem_U20228 ( .A1(MEM_stage_inst_dmem_n21474), .A2(MEM_stage_inst_dmem_n20620), .ZN(MEM_stage_inst_dmem_n20595) );
NAND2_X1 MEM_stage_inst_dmem_U20227 ( .A1(MEM_stage_inst_dmem_ram_3996), .A2(MEM_stage_inst_dmem_n20619), .ZN(MEM_stage_inst_dmem_n20596) );
NAND2_X1 MEM_stage_inst_dmem_U20226 ( .A1(MEM_stage_inst_dmem_n20594), .A2(MEM_stage_inst_dmem_n20593), .ZN(MEM_stage_inst_dmem_n9176) );
NAND2_X1 MEM_stage_inst_dmem_U20225 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n20620), .ZN(MEM_stage_inst_dmem_n20593) );
NAND2_X1 MEM_stage_inst_dmem_U20224 ( .A1(MEM_stage_inst_dmem_ram_3997), .A2(MEM_stage_inst_dmem_n20619), .ZN(MEM_stage_inst_dmem_n20594) );
NAND2_X1 MEM_stage_inst_dmem_U20223 ( .A1(MEM_stage_inst_dmem_n20592), .A2(MEM_stage_inst_dmem_n20591), .ZN(MEM_stage_inst_dmem_n9177) );
NAND2_X1 MEM_stage_inst_dmem_U20222 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n20620), .ZN(MEM_stage_inst_dmem_n20591) );
NAND2_X1 MEM_stage_inst_dmem_U20221 ( .A1(MEM_stage_inst_dmem_ram_3998), .A2(MEM_stage_inst_dmem_n20619), .ZN(MEM_stage_inst_dmem_n20592) );
NAND2_X1 MEM_stage_inst_dmem_U20220 ( .A1(MEM_stage_inst_dmem_n20590), .A2(MEM_stage_inst_dmem_n20589), .ZN(MEM_stage_inst_dmem_n9178) );
NAND2_X1 MEM_stage_inst_dmem_U20219 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n20620), .ZN(MEM_stage_inst_dmem_n20589) );
NAND2_X1 MEM_stage_inst_dmem_U20218 ( .A1(MEM_stage_inst_dmem_ram_3999), .A2(MEM_stage_inst_dmem_n20619), .ZN(MEM_stage_inst_dmem_n20590) );
NAND2_X1 MEM_stage_inst_dmem_U20217 ( .A1(MEM_stage_inst_dmem_n21144), .A2(MEM_stage_inst_dmem_n20895), .ZN(MEM_stage_inst_dmem_n20619) );
NAND2_X1 MEM_stage_inst_dmem_U20216 ( .A1(MEM_stage_inst_dmem_n20588), .A2(MEM_stage_inst_dmem_n20587), .ZN(MEM_stage_inst_dmem_n9179) );
NAND2_X1 MEM_stage_inst_dmem_U20215 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n20586), .ZN(MEM_stage_inst_dmem_n20587) );
NAND2_X1 MEM_stage_inst_dmem_U20214 ( .A1(MEM_stage_inst_dmem_ram_4000), .A2(MEM_stage_inst_dmem_n20585), .ZN(MEM_stage_inst_dmem_n20588) );
NAND2_X1 MEM_stage_inst_dmem_U20213 ( .A1(MEM_stage_inst_dmem_n20584), .A2(MEM_stage_inst_dmem_n20583), .ZN(MEM_stage_inst_dmem_n9180) );
NAND2_X1 MEM_stage_inst_dmem_U20212 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n20586), .ZN(MEM_stage_inst_dmem_n20583) );
NAND2_X1 MEM_stage_inst_dmem_U20211 ( .A1(MEM_stage_inst_dmem_ram_4001), .A2(MEM_stage_inst_dmem_n20585), .ZN(MEM_stage_inst_dmem_n20584) );
NAND2_X1 MEM_stage_inst_dmem_U20210 ( .A1(MEM_stage_inst_dmem_n20582), .A2(MEM_stage_inst_dmem_n20581), .ZN(MEM_stage_inst_dmem_n9181) );
NAND2_X1 MEM_stage_inst_dmem_U20209 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n20586), .ZN(MEM_stage_inst_dmem_n20581) );
NAND2_X1 MEM_stage_inst_dmem_U20208 ( .A1(MEM_stage_inst_dmem_ram_4002), .A2(MEM_stage_inst_dmem_n20585), .ZN(MEM_stage_inst_dmem_n20582) );
NAND2_X1 MEM_stage_inst_dmem_U20207 ( .A1(MEM_stage_inst_dmem_n20580), .A2(MEM_stage_inst_dmem_n20579), .ZN(MEM_stage_inst_dmem_n9182) );
NAND2_X1 MEM_stage_inst_dmem_U20206 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n20586), .ZN(MEM_stage_inst_dmem_n20579) );
NAND2_X1 MEM_stage_inst_dmem_U20205 ( .A1(MEM_stage_inst_dmem_ram_4003), .A2(MEM_stage_inst_dmem_n20585), .ZN(MEM_stage_inst_dmem_n20580) );
NAND2_X1 MEM_stage_inst_dmem_U20204 ( .A1(MEM_stage_inst_dmem_n20578), .A2(MEM_stage_inst_dmem_n20577), .ZN(MEM_stage_inst_dmem_n9183) );
NAND2_X1 MEM_stage_inst_dmem_U20203 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n20586), .ZN(MEM_stage_inst_dmem_n20577) );
NAND2_X1 MEM_stage_inst_dmem_U20202 ( .A1(MEM_stage_inst_dmem_ram_4004), .A2(MEM_stage_inst_dmem_n20585), .ZN(MEM_stage_inst_dmem_n20578) );
NAND2_X1 MEM_stage_inst_dmem_U20201 ( .A1(MEM_stage_inst_dmem_n20576), .A2(MEM_stage_inst_dmem_n20575), .ZN(MEM_stage_inst_dmem_n9184) );
NAND2_X1 MEM_stage_inst_dmem_U20200 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n20586), .ZN(MEM_stage_inst_dmem_n20575) );
NAND2_X1 MEM_stage_inst_dmem_U20199 ( .A1(MEM_stage_inst_dmem_ram_4005), .A2(MEM_stage_inst_dmem_n20585), .ZN(MEM_stage_inst_dmem_n20576) );
NAND2_X1 MEM_stage_inst_dmem_U20198 ( .A1(MEM_stage_inst_dmem_n20574), .A2(MEM_stage_inst_dmem_n20573), .ZN(MEM_stage_inst_dmem_n9185) );
NAND2_X1 MEM_stage_inst_dmem_U20197 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n20586), .ZN(MEM_stage_inst_dmem_n20573) );
NAND2_X1 MEM_stage_inst_dmem_U20196 ( .A1(MEM_stage_inst_dmem_ram_4006), .A2(MEM_stage_inst_dmem_n20585), .ZN(MEM_stage_inst_dmem_n20574) );
NAND2_X1 MEM_stage_inst_dmem_U20195 ( .A1(MEM_stage_inst_dmem_n20572), .A2(MEM_stage_inst_dmem_n20571), .ZN(MEM_stage_inst_dmem_n9186) );
NAND2_X1 MEM_stage_inst_dmem_U20194 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n20586), .ZN(MEM_stage_inst_dmem_n20571) );
NAND2_X1 MEM_stage_inst_dmem_U20193 ( .A1(MEM_stage_inst_dmem_ram_4007), .A2(MEM_stage_inst_dmem_n20585), .ZN(MEM_stage_inst_dmem_n20572) );
NAND2_X1 MEM_stage_inst_dmem_U20192 ( .A1(MEM_stage_inst_dmem_n20570), .A2(MEM_stage_inst_dmem_n20569), .ZN(MEM_stage_inst_dmem_n9187) );
NAND2_X1 MEM_stage_inst_dmem_U20191 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n20586), .ZN(MEM_stage_inst_dmem_n20569) );
NAND2_X1 MEM_stage_inst_dmem_U20190 ( .A1(MEM_stage_inst_dmem_ram_4008), .A2(MEM_stage_inst_dmem_n20585), .ZN(MEM_stage_inst_dmem_n20570) );
NAND2_X1 MEM_stage_inst_dmem_U20189 ( .A1(MEM_stage_inst_dmem_n20568), .A2(MEM_stage_inst_dmem_n20567), .ZN(MEM_stage_inst_dmem_n9188) );
NAND2_X1 MEM_stage_inst_dmem_U20188 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n20586), .ZN(MEM_stage_inst_dmem_n20567) );
NAND2_X1 MEM_stage_inst_dmem_U20187 ( .A1(MEM_stage_inst_dmem_ram_4009), .A2(MEM_stage_inst_dmem_n20585), .ZN(MEM_stage_inst_dmem_n20568) );
NAND2_X1 MEM_stage_inst_dmem_U20186 ( .A1(MEM_stage_inst_dmem_n20566), .A2(MEM_stage_inst_dmem_n20565), .ZN(MEM_stage_inst_dmem_n9189) );
NAND2_X1 MEM_stage_inst_dmem_U20185 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n20586), .ZN(MEM_stage_inst_dmem_n20565) );
NAND2_X1 MEM_stage_inst_dmem_U20184 ( .A1(MEM_stage_inst_dmem_ram_4010), .A2(MEM_stage_inst_dmem_n20585), .ZN(MEM_stage_inst_dmem_n20566) );
NAND2_X1 MEM_stage_inst_dmem_U20183 ( .A1(MEM_stage_inst_dmem_n20564), .A2(MEM_stage_inst_dmem_n20563), .ZN(MEM_stage_inst_dmem_n9190) );
NAND2_X1 MEM_stage_inst_dmem_U20182 ( .A1(MEM_stage_inst_dmem_n14705), .A2(MEM_stage_inst_dmem_n20586), .ZN(MEM_stage_inst_dmem_n20563) );
NAND2_X1 MEM_stage_inst_dmem_U20181 ( .A1(MEM_stage_inst_dmem_ram_4011), .A2(MEM_stage_inst_dmem_n20585), .ZN(MEM_stage_inst_dmem_n20564) );
NAND2_X1 MEM_stage_inst_dmem_U20180 ( .A1(MEM_stage_inst_dmem_n20562), .A2(MEM_stage_inst_dmem_n20561), .ZN(MEM_stage_inst_dmem_n9191) );
NAND2_X1 MEM_stage_inst_dmem_U20179 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n20586), .ZN(MEM_stage_inst_dmem_n20561) );
NAND2_X1 MEM_stage_inst_dmem_U20178 ( .A1(MEM_stage_inst_dmem_ram_4012), .A2(MEM_stage_inst_dmem_n20585), .ZN(MEM_stage_inst_dmem_n20562) );
NAND2_X1 MEM_stage_inst_dmem_U20177 ( .A1(MEM_stage_inst_dmem_n20560), .A2(MEM_stage_inst_dmem_n20559), .ZN(MEM_stage_inst_dmem_n9192) );
NAND2_X1 MEM_stage_inst_dmem_U20176 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n20586), .ZN(MEM_stage_inst_dmem_n20559) );
NAND2_X1 MEM_stage_inst_dmem_U20175 ( .A1(MEM_stage_inst_dmem_ram_4013), .A2(MEM_stage_inst_dmem_n20585), .ZN(MEM_stage_inst_dmem_n20560) );
NAND2_X1 MEM_stage_inst_dmem_U20174 ( .A1(MEM_stage_inst_dmem_n20558), .A2(MEM_stage_inst_dmem_n20557), .ZN(MEM_stage_inst_dmem_n9193) );
NAND2_X1 MEM_stage_inst_dmem_U20173 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n20586), .ZN(MEM_stage_inst_dmem_n20557) );
NAND2_X1 MEM_stage_inst_dmem_U20172 ( .A1(MEM_stage_inst_dmem_ram_4014), .A2(MEM_stage_inst_dmem_n20585), .ZN(MEM_stage_inst_dmem_n20558) );
NAND2_X1 MEM_stage_inst_dmem_U20171 ( .A1(MEM_stage_inst_dmem_n20556), .A2(MEM_stage_inst_dmem_n20555), .ZN(MEM_stage_inst_dmem_n9194) );
NAND2_X1 MEM_stage_inst_dmem_U20170 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n20586), .ZN(MEM_stage_inst_dmem_n20555) );
INV_X1 MEM_stage_inst_dmem_U20169 ( .A(MEM_stage_inst_dmem_n20585), .ZN(MEM_stage_inst_dmem_n20586) );
NAND2_X1 MEM_stage_inst_dmem_U20168 ( .A1(MEM_stage_inst_dmem_ram_4015), .A2(MEM_stage_inst_dmem_n20585), .ZN(MEM_stage_inst_dmem_n20556) );
NAND2_X1 MEM_stage_inst_dmem_U20167 ( .A1(MEM_stage_inst_dmem_n21109), .A2(MEM_stage_inst_dmem_n20895), .ZN(MEM_stage_inst_dmem_n20585) );
NAND2_X1 MEM_stage_inst_dmem_U20166 ( .A1(MEM_stage_inst_dmem_n20554), .A2(MEM_stage_inst_dmem_n20553), .ZN(MEM_stage_inst_dmem_n9195) );
NAND2_X1 MEM_stage_inst_dmem_U20165 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n20552), .ZN(MEM_stage_inst_dmem_n20553) );
NAND2_X1 MEM_stage_inst_dmem_U20164 ( .A1(MEM_stage_inst_dmem_ram_4016), .A2(MEM_stage_inst_dmem_n20550), .ZN(MEM_stage_inst_dmem_n20554) );
NAND2_X1 MEM_stage_inst_dmem_U20163 ( .A1(MEM_stage_inst_dmem_n20549), .A2(MEM_stage_inst_dmem_n20548), .ZN(MEM_stage_inst_dmem_n9196) );
NAND2_X1 MEM_stage_inst_dmem_U20162 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n20552), .ZN(MEM_stage_inst_dmem_n20548) );
NAND2_X1 MEM_stage_inst_dmem_U20161 ( .A1(MEM_stage_inst_dmem_ram_4017), .A2(MEM_stage_inst_dmem_n20550), .ZN(MEM_stage_inst_dmem_n20549) );
NAND2_X1 MEM_stage_inst_dmem_U20160 ( .A1(MEM_stage_inst_dmem_n20546), .A2(MEM_stage_inst_dmem_n20545), .ZN(MEM_stage_inst_dmem_n9197) );
NAND2_X1 MEM_stage_inst_dmem_U20159 ( .A1(MEM_stage_inst_dmem_n18887), .A2(MEM_stage_inst_dmem_n20552), .ZN(MEM_stage_inst_dmem_n20545) );
NAND2_X1 MEM_stage_inst_dmem_U20158 ( .A1(MEM_stage_inst_dmem_ram_4018), .A2(MEM_stage_inst_dmem_n20550), .ZN(MEM_stage_inst_dmem_n20546) );
NAND2_X1 MEM_stage_inst_dmem_U20157 ( .A1(MEM_stage_inst_dmem_n20543), .A2(MEM_stage_inst_dmem_n20542), .ZN(MEM_stage_inst_dmem_n9198) );
NAND2_X1 MEM_stage_inst_dmem_U20156 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n20552), .ZN(MEM_stage_inst_dmem_n20542) );
NAND2_X1 MEM_stage_inst_dmem_U20155 ( .A1(MEM_stage_inst_dmem_ram_4019), .A2(MEM_stage_inst_dmem_n20550), .ZN(MEM_stage_inst_dmem_n20543) );
NAND2_X1 MEM_stage_inst_dmem_U20154 ( .A1(MEM_stage_inst_dmem_n20540), .A2(MEM_stage_inst_dmem_n20539), .ZN(MEM_stage_inst_dmem_n9199) );
NAND2_X1 MEM_stage_inst_dmem_U20153 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n20552), .ZN(MEM_stage_inst_dmem_n20539) );
NAND2_X1 MEM_stage_inst_dmem_U20152 ( .A1(MEM_stage_inst_dmem_ram_4020), .A2(MEM_stage_inst_dmem_n20550), .ZN(MEM_stage_inst_dmem_n20540) );
NAND2_X1 MEM_stage_inst_dmem_U20151 ( .A1(MEM_stage_inst_dmem_n20538), .A2(MEM_stage_inst_dmem_n20537), .ZN(MEM_stage_inst_dmem_n9200) );
NAND2_X1 MEM_stage_inst_dmem_U20150 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n20552), .ZN(MEM_stage_inst_dmem_n20537) );
NAND2_X1 MEM_stage_inst_dmem_U20149 ( .A1(MEM_stage_inst_dmem_ram_4021), .A2(MEM_stage_inst_dmem_n20550), .ZN(MEM_stage_inst_dmem_n20538) );
NAND2_X1 MEM_stage_inst_dmem_U20148 ( .A1(MEM_stage_inst_dmem_n20535), .A2(MEM_stage_inst_dmem_n20534), .ZN(MEM_stage_inst_dmem_n9201) );
NAND2_X1 MEM_stage_inst_dmem_U20147 ( .A1(MEM_stage_inst_dmem_n14717), .A2(MEM_stage_inst_dmem_n20552), .ZN(MEM_stage_inst_dmem_n20534) );
NAND2_X1 MEM_stage_inst_dmem_U20146 ( .A1(MEM_stage_inst_dmem_ram_4022), .A2(MEM_stage_inst_dmem_n20550), .ZN(MEM_stage_inst_dmem_n20535) );
NAND2_X1 MEM_stage_inst_dmem_U20145 ( .A1(MEM_stage_inst_dmem_n20532), .A2(MEM_stage_inst_dmem_n20531), .ZN(MEM_stage_inst_dmem_n9202) );
NAND2_X1 MEM_stage_inst_dmem_U20144 ( .A1(MEM_stage_inst_dmem_n16361), .A2(MEM_stage_inst_dmem_n20552), .ZN(MEM_stage_inst_dmem_n20531) );
NAND2_X1 MEM_stage_inst_dmem_U20143 ( .A1(MEM_stage_inst_dmem_ram_4023), .A2(MEM_stage_inst_dmem_n20550), .ZN(MEM_stage_inst_dmem_n20532) );
NAND2_X1 MEM_stage_inst_dmem_U20142 ( .A1(MEM_stage_inst_dmem_n20529), .A2(MEM_stage_inst_dmem_n20528), .ZN(MEM_stage_inst_dmem_n9203) );
NAND2_X1 MEM_stage_inst_dmem_U20141 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n20552), .ZN(MEM_stage_inst_dmem_n20528) );
NAND2_X1 MEM_stage_inst_dmem_U20140 ( .A1(MEM_stage_inst_dmem_ram_4024), .A2(MEM_stage_inst_dmem_n20550), .ZN(MEM_stage_inst_dmem_n20529) );
NAND2_X1 MEM_stage_inst_dmem_U20139 ( .A1(MEM_stage_inst_dmem_n20526), .A2(MEM_stage_inst_dmem_n20525), .ZN(MEM_stage_inst_dmem_n9204) );
NAND2_X1 MEM_stage_inst_dmem_U20138 ( .A1(MEM_stage_inst_dmem_n96), .A2(MEM_stage_inst_dmem_n20552), .ZN(MEM_stage_inst_dmem_n20525) );
NAND2_X1 MEM_stage_inst_dmem_U20137 ( .A1(MEM_stage_inst_dmem_ram_4025), .A2(MEM_stage_inst_dmem_n20550), .ZN(MEM_stage_inst_dmem_n20526) );
NAND2_X1 MEM_stage_inst_dmem_U20136 ( .A1(MEM_stage_inst_dmem_n20523), .A2(MEM_stage_inst_dmem_n20522), .ZN(MEM_stage_inst_dmem_n9205) );
NAND2_X1 MEM_stage_inst_dmem_U20135 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n20552), .ZN(MEM_stage_inst_dmem_n20522) );
NAND2_X1 MEM_stage_inst_dmem_U20134 ( .A1(MEM_stage_inst_dmem_ram_4026), .A2(MEM_stage_inst_dmem_n20550), .ZN(MEM_stage_inst_dmem_n20523) );
NAND2_X1 MEM_stage_inst_dmem_U20133 ( .A1(MEM_stage_inst_dmem_n20520), .A2(MEM_stage_inst_dmem_n20519), .ZN(MEM_stage_inst_dmem_n9206) );
NAND2_X1 MEM_stage_inst_dmem_U20132 ( .A1(MEM_stage_inst_dmem_n20904), .A2(MEM_stage_inst_dmem_n20552), .ZN(MEM_stage_inst_dmem_n20519) );
NAND2_X1 MEM_stage_inst_dmem_U20131 ( .A1(MEM_stage_inst_dmem_ram_4027), .A2(MEM_stage_inst_dmem_n20550), .ZN(MEM_stage_inst_dmem_n20520) );
NAND2_X1 MEM_stage_inst_dmem_U20130 ( .A1(MEM_stage_inst_dmem_n20517), .A2(MEM_stage_inst_dmem_n20516), .ZN(MEM_stage_inst_dmem_n9207) );
NAND2_X1 MEM_stage_inst_dmem_U20129 ( .A1(MEM_stage_inst_dmem_n21474), .A2(MEM_stage_inst_dmem_n20552), .ZN(MEM_stage_inst_dmem_n20516) );
NAND2_X1 MEM_stage_inst_dmem_U20128 ( .A1(MEM_stage_inst_dmem_ram_4028), .A2(MEM_stage_inst_dmem_n20550), .ZN(MEM_stage_inst_dmem_n20517) );
NAND2_X1 MEM_stage_inst_dmem_U20127 ( .A1(MEM_stage_inst_dmem_n20514), .A2(MEM_stage_inst_dmem_n20513), .ZN(MEM_stage_inst_dmem_n9208) );
NAND2_X1 MEM_stage_inst_dmem_U20126 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n20552), .ZN(MEM_stage_inst_dmem_n20513) );
NAND2_X1 MEM_stage_inst_dmem_U20125 ( .A1(MEM_stage_inst_dmem_ram_4029), .A2(MEM_stage_inst_dmem_n20550), .ZN(MEM_stage_inst_dmem_n20514) );
NAND2_X1 MEM_stage_inst_dmem_U20124 ( .A1(MEM_stage_inst_dmem_n20511), .A2(MEM_stage_inst_dmem_n20510), .ZN(MEM_stage_inst_dmem_n9209) );
NAND2_X1 MEM_stage_inst_dmem_U20123 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n20552), .ZN(MEM_stage_inst_dmem_n20510) );
NAND2_X1 MEM_stage_inst_dmem_U20122 ( .A1(MEM_stage_inst_dmem_ram_4030), .A2(MEM_stage_inst_dmem_n20550), .ZN(MEM_stage_inst_dmem_n20511) );
NAND2_X1 MEM_stage_inst_dmem_U20121 ( .A1(MEM_stage_inst_dmem_n20508), .A2(MEM_stage_inst_dmem_n20507), .ZN(MEM_stage_inst_dmem_n9210) );
NAND2_X1 MEM_stage_inst_dmem_U20120 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n20552), .ZN(MEM_stage_inst_dmem_n20507) );
INV_X1 MEM_stage_inst_dmem_U20119 ( .A(MEM_stage_inst_dmem_n20550), .ZN(MEM_stage_inst_dmem_n20552) );
NAND2_X1 MEM_stage_inst_dmem_U20118 ( .A1(MEM_stage_inst_dmem_ram_4031), .A2(MEM_stage_inst_dmem_n20550), .ZN(MEM_stage_inst_dmem_n20508) );
NAND2_X1 MEM_stage_inst_dmem_U20117 ( .A1(MEM_stage_inst_dmem_n21074), .A2(MEM_stage_inst_dmem_n20895), .ZN(MEM_stage_inst_dmem_n20550) );
NAND2_X1 MEM_stage_inst_dmem_U20116 ( .A1(MEM_stage_inst_dmem_n20505), .A2(MEM_stage_inst_dmem_n20504), .ZN(MEM_stage_inst_dmem_n9211) );
NAND2_X1 MEM_stage_inst_dmem_U20115 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n20503), .ZN(MEM_stage_inst_dmem_n20504) );
NAND2_X1 MEM_stage_inst_dmem_U20114 ( .A1(MEM_stage_inst_dmem_ram_4032), .A2(MEM_stage_inst_dmem_n20502), .ZN(MEM_stage_inst_dmem_n20505) );
NAND2_X1 MEM_stage_inst_dmem_U20113 ( .A1(MEM_stage_inst_dmem_n20501), .A2(MEM_stage_inst_dmem_n20500), .ZN(MEM_stage_inst_dmem_n9212) );
NAND2_X1 MEM_stage_inst_dmem_U20112 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n20503), .ZN(MEM_stage_inst_dmem_n20500) );
NAND2_X1 MEM_stage_inst_dmem_U20111 ( .A1(MEM_stage_inst_dmem_ram_4033), .A2(MEM_stage_inst_dmem_n20502), .ZN(MEM_stage_inst_dmem_n20501) );
NAND2_X1 MEM_stage_inst_dmem_U20110 ( .A1(MEM_stage_inst_dmem_n20499), .A2(MEM_stage_inst_dmem_n20498), .ZN(MEM_stage_inst_dmem_n9213) );
NAND2_X1 MEM_stage_inst_dmem_U20109 ( .A1(MEM_stage_inst_dmem_n20544), .A2(MEM_stage_inst_dmem_n20503), .ZN(MEM_stage_inst_dmem_n20498) );
NAND2_X1 MEM_stage_inst_dmem_U20108 ( .A1(MEM_stage_inst_dmem_ram_4034), .A2(MEM_stage_inst_dmem_n20502), .ZN(MEM_stage_inst_dmem_n20499) );
NAND2_X1 MEM_stage_inst_dmem_U20107 ( .A1(MEM_stage_inst_dmem_n20497), .A2(MEM_stage_inst_dmem_n20496), .ZN(MEM_stage_inst_dmem_n9214) );
NAND2_X1 MEM_stage_inst_dmem_U20106 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n20503), .ZN(MEM_stage_inst_dmem_n20496) );
NAND2_X1 MEM_stage_inst_dmem_U20105 ( .A1(MEM_stage_inst_dmem_ram_4035), .A2(MEM_stage_inst_dmem_n20502), .ZN(MEM_stage_inst_dmem_n20497) );
NAND2_X1 MEM_stage_inst_dmem_U20104 ( .A1(MEM_stage_inst_dmem_n20495), .A2(MEM_stage_inst_dmem_n20494), .ZN(MEM_stage_inst_dmem_n9215) );
NAND2_X1 MEM_stage_inst_dmem_U20103 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n20503), .ZN(MEM_stage_inst_dmem_n20494) );
NAND2_X1 MEM_stage_inst_dmem_U20102 ( .A1(MEM_stage_inst_dmem_ram_4036), .A2(MEM_stage_inst_dmem_n20502), .ZN(MEM_stage_inst_dmem_n20495) );
NAND2_X1 MEM_stage_inst_dmem_U20101 ( .A1(MEM_stage_inst_dmem_n20493), .A2(MEM_stage_inst_dmem_n20492), .ZN(MEM_stage_inst_dmem_n9216) );
NAND2_X1 MEM_stage_inst_dmem_U20100 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n20503), .ZN(MEM_stage_inst_dmem_n20492) );
NAND2_X1 MEM_stage_inst_dmem_U20099 ( .A1(MEM_stage_inst_dmem_ram_4037), .A2(MEM_stage_inst_dmem_n20502), .ZN(MEM_stage_inst_dmem_n20493) );
NAND2_X1 MEM_stage_inst_dmem_U20098 ( .A1(MEM_stage_inst_dmem_n20491), .A2(MEM_stage_inst_dmem_n20490), .ZN(MEM_stage_inst_dmem_n9217) );
NAND2_X1 MEM_stage_inst_dmem_U20097 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n20503), .ZN(MEM_stage_inst_dmem_n20490) );
NAND2_X1 MEM_stage_inst_dmem_U20096 ( .A1(MEM_stage_inst_dmem_ram_4038), .A2(MEM_stage_inst_dmem_n20502), .ZN(MEM_stage_inst_dmem_n20491) );
NAND2_X1 MEM_stage_inst_dmem_U20095 ( .A1(MEM_stage_inst_dmem_n20489), .A2(MEM_stage_inst_dmem_n20488), .ZN(MEM_stage_inst_dmem_n9218) );
NAND2_X1 MEM_stage_inst_dmem_U20094 ( .A1(MEM_stage_inst_dmem_n20530), .A2(MEM_stage_inst_dmem_n20503), .ZN(MEM_stage_inst_dmem_n20488) );
NAND2_X1 MEM_stage_inst_dmem_U20093 ( .A1(MEM_stage_inst_dmem_ram_4039), .A2(MEM_stage_inst_dmem_n20502), .ZN(MEM_stage_inst_dmem_n20489) );
NAND2_X1 MEM_stage_inst_dmem_U20092 ( .A1(MEM_stage_inst_dmem_n20487), .A2(MEM_stage_inst_dmem_n20486), .ZN(MEM_stage_inst_dmem_n9219) );
NAND2_X1 MEM_stage_inst_dmem_U20091 ( .A1(MEM_stage_inst_dmem_n18013), .A2(MEM_stage_inst_dmem_n20503), .ZN(MEM_stage_inst_dmem_n20486) );
NAND2_X1 MEM_stage_inst_dmem_U20090 ( .A1(MEM_stage_inst_dmem_ram_4040), .A2(MEM_stage_inst_dmem_n20502), .ZN(MEM_stage_inst_dmem_n20487) );
NAND2_X1 MEM_stage_inst_dmem_U20089 ( .A1(MEM_stage_inst_dmem_n20485), .A2(MEM_stage_inst_dmem_n20484), .ZN(MEM_stage_inst_dmem_n9220) );
NAND2_X1 MEM_stage_inst_dmem_U20088 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n20503), .ZN(MEM_stage_inst_dmem_n20484) );
NAND2_X1 MEM_stage_inst_dmem_U20087 ( .A1(MEM_stage_inst_dmem_ram_4041), .A2(MEM_stage_inst_dmem_n20502), .ZN(MEM_stage_inst_dmem_n20485) );
NAND2_X1 MEM_stage_inst_dmem_U20086 ( .A1(MEM_stage_inst_dmem_n20483), .A2(MEM_stage_inst_dmem_n20482), .ZN(MEM_stage_inst_dmem_n9221) );
NAND2_X1 MEM_stage_inst_dmem_U20085 ( .A1(MEM_stage_inst_dmem_n20521), .A2(MEM_stage_inst_dmem_n20503), .ZN(MEM_stage_inst_dmem_n20482) );
NAND2_X1 MEM_stage_inst_dmem_U20084 ( .A1(MEM_stage_inst_dmem_ram_4042), .A2(MEM_stage_inst_dmem_n20502), .ZN(MEM_stage_inst_dmem_n20483) );
NAND2_X1 MEM_stage_inst_dmem_U20083 ( .A1(MEM_stage_inst_dmem_n20481), .A2(MEM_stage_inst_dmem_n20480), .ZN(MEM_stage_inst_dmem_n9222) );
NAND2_X1 MEM_stage_inst_dmem_U20082 ( .A1(MEM_stage_inst_dmem_n14705), .A2(MEM_stage_inst_dmem_n20503), .ZN(MEM_stage_inst_dmem_n20480) );
NAND2_X1 MEM_stage_inst_dmem_U20081 ( .A1(MEM_stage_inst_dmem_ram_4043), .A2(MEM_stage_inst_dmem_n20502), .ZN(MEM_stage_inst_dmem_n20481) );
NAND2_X1 MEM_stage_inst_dmem_U20080 ( .A1(MEM_stage_inst_dmem_n20479), .A2(MEM_stage_inst_dmem_n20478), .ZN(MEM_stage_inst_dmem_n9223) );
NAND2_X1 MEM_stage_inst_dmem_U20079 ( .A1(MEM_stage_inst_dmem_n14702), .A2(MEM_stage_inst_dmem_n20503), .ZN(MEM_stage_inst_dmem_n20478) );
NAND2_X1 MEM_stage_inst_dmem_U20078 ( .A1(MEM_stage_inst_dmem_ram_4044), .A2(MEM_stage_inst_dmem_n20502), .ZN(MEM_stage_inst_dmem_n20479) );
NAND2_X1 MEM_stage_inst_dmem_U20077 ( .A1(MEM_stage_inst_dmem_n20477), .A2(MEM_stage_inst_dmem_n20476), .ZN(MEM_stage_inst_dmem_n9224) );
NAND2_X1 MEM_stage_inst_dmem_U20076 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n20503), .ZN(MEM_stage_inst_dmem_n20476) );
NAND2_X1 MEM_stage_inst_dmem_U20075 ( .A1(MEM_stage_inst_dmem_ram_4045), .A2(MEM_stage_inst_dmem_n20502), .ZN(MEM_stage_inst_dmem_n20477) );
NAND2_X1 MEM_stage_inst_dmem_U20074 ( .A1(MEM_stage_inst_dmem_n20475), .A2(MEM_stage_inst_dmem_n20474), .ZN(MEM_stage_inst_dmem_n9225) );
NAND2_X1 MEM_stage_inst_dmem_U20073 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n20503), .ZN(MEM_stage_inst_dmem_n20474) );
NAND2_X1 MEM_stage_inst_dmem_U20072 ( .A1(MEM_stage_inst_dmem_ram_4046), .A2(MEM_stage_inst_dmem_n20502), .ZN(MEM_stage_inst_dmem_n20475) );
NAND2_X1 MEM_stage_inst_dmem_U20071 ( .A1(MEM_stage_inst_dmem_n20473), .A2(MEM_stage_inst_dmem_n20472), .ZN(MEM_stage_inst_dmem_n9226) );
NAND2_X1 MEM_stage_inst_dmem_U20070 ( .A1(MEM_stage_inst_dmem_n15110), .A2(MEM_stage_inst_dmem_n20503), .ZN(MEM_stage_inst_dmem_n20472) );
INV_X1 MEM_stage_inst_dmem_U20069 ( .A(MEM_stage_inst_dmem_n20502), .ZN(MEM_stage_inst_dmem_n20503) );
NAND2_X1 MEM_stage_inst_dmem_U20068 ( .A1(MEM_stage_inst_dmem_ram_4047), .A2(MEM_stage_inst_dmem_n20502), .ZN(MEM_stage_inst_dmem_n20473) );
NAND2_X1 MEM_stage_inst_dmem_U20067 ( .A1(MEM_stage_inst_dmem_n21039), .A2(MEM_stage_inst_dmem_n20895), .ZN(MEM_stage_inst_dmem_n20502) );
NAND2_X1 MEM_stage_inst_dmem_U20066 ( .A1(MEM_stage_inst_dmem_n20471), .A2(MEM_stage_inst_dmem_n20470), .ZN(MEM_stage_inst_dmem_n9227) );
NAND2_X1 MEM_stage_inst_dmem_U20065 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n20469), .ZN(MEM_stage_inst_dmem_n20470) );
NAND2_X1 MEM_stage_inst_dmem_U20064 ( .A1(MEM_stage_inst_dmem_ram_4048), .A2(MEM_stage_inst_dmem_n20468), .ZN(MEM_stage_inst_dmem_n20471) );
NAND2_X1 MEM_stage_inst_dmem_U20063 ( .A1(MEM_stage_inst_dmem_n20467), .A2(MEM_stage_inst_dmem_n20466), .ZN(MEM_stage_inst_dmem_n9228) );
NAND2_X1 MEM_stage_inst_dmem_U20062 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n20469), .ZN(MEM_stage_inst_dmem_n20466) );
NAND2_X1 MEM_stage_inst_dmem_U20061 ( .A1(MEM_stage_inst_dmem_ram_4049), .A2(MEM_stage_inst_dmem_n20468), .ZN(MEM_stage_inst_dmem_n20467) );
NAND2_X1 MEM_stage_inst_dmem_U20060 ( .A1(MEM_stage_inst_dmem_n20465), .A2(MEM_stage_inst_dmem_n20464), .ZN(MEM_stage_inst_dmem_n9229) );
NAND2_X1 MEM_stage_inst_dmem_U20059 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n20469), .ZN(MEM_stage_inst_dmem_n20464) );
NAND2_X1 MEM_stage_inst_dmem_U20058 ( .A1(MEM_stage_inst_dmem_ram_4050), .A2(MEM_stage_inst_dmem_n20468), .ZN(MEM_stage_inst_dmem_n20465) );
NAND2_X1 MEM_stage_inst_dmem_U20057 ( .A1(MEM_stage_inst_dmem_n20463), .A2(MEM_stage_inst_dmem_n20462), .ZN(MEM_stage_inst_dmem_n9230) );
NAND2_X1 MEM_stage_inst_dmem_U20056 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n20469), .ZN(MEM_stage_inst_dmem_n20462) );
NAND2_X1 MEM_stage_inst_dmem_U20055 ( .A1(MEM_stage_inst_dmem_ram_4051), .A2(MEM_stage_inst_dmem_n20468), .ZN(MEM_stage_inst_dmem_n20463) );
NAND2_X1 MEM_stage_inst_dmem_U20054 ( .A1(MEM_stage_inst_dmem_n20461), .A2(MEM_stage_inst_dmem_n20460), .ZN(MEM_stage_inst_dmem_n9231) );
NAND2_X1 MEM_stage_inst_dmem_U20053 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n20469), .ZN(MEM_stage_inst_dmem_n20460) );
NAND2_X1 MEM_stage_inst_dmem_U20052 ( .A1(MEM_stage_inst_dmem_ram_4052), .A2(MEM_stage_inst_dmem_n20468), .ZN(MEM_stage_inst_dmem_n20461) );
NAND2_X1 MEM_stage_inst_dmem_U20051 ( .A1(MEM_stage_inst_dmem_n20459), .A2(MEM_stage_inst_dmem_n20458), .ZN(MEM_stage_inst_dmem_n9232) );
NAND2_X1 MEM_stage_inst_dmem_U20050 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n20469), .ZN(MEM_stage_inst_dmem_n20458) );
NAND2_X1 MEM_stage_inst_dmem_U20049 ( .A1(MEM_stage_inst_dmem_ram_4053), .A2(MEM_stage_inst_dmem_n20468), .ZN(MEM_stage_inst_dmem_n20459) );
NAND2_X1 MEM_stage_inst_dmem_U20048 ( .A1(MEM_stage_inst_dmem_n20457), .A2(MEM_stage_inst_dmem_n20456), .ZN(MEM_stage_inst_dmem_n9233) );
NAND2_X1 MEM_stage_inst_dmem_U20047 ( .A1(MEM_stage_inst_dmem_n14717), .A2(MEM_stage_inst_dmem_n20469), .ZN(MEM_stage_inst_dmem_n20456) );
NAND2_X1 MEM_stage_inst_dmem_U20046 ( .A1(MEM_stage_inst_dmem_ram_4054), .A2(MEM_stage_inst_dmem_n20468), .ZN(MEM_stage_inst_dmem_n20457) );
NAND2_X1 MEM_stage_inst_dmem_U20045 ( .A1(MEM_stage_inst_dmem_n20455), .A2(MEM_stage_inst_dmem_n20454), .ZN(MEM_stage_inst_dmem_n9234) );
NAND2_X1 MEM_stage_inst_dmem_U20044 ( .A1(MEM_stage_inst_dmem_n18), .A2(MEM_stage_inst_dmem_n20469), .ZN(MEM_stage_inst_dmem_n20454) );
NAND2_X1 MEM_stage_inst_dmem_U20043 ( .A1(MEM_stage_inst_dmem_ram_4055), .A2(MEM_stage_inst_dmem_n20468), .ZN(MEM_stage_inst_dmem_n20455) );
NAND2_X1 MEM_stage_inst_dmem_U20042 ( .A1(MEM_stage_inst_dmem_n20453), .A2(MEM_stage_inst_dmem_n20452), .ZN(MEM_stage_inst_dmem_n9235) );
NAND2_X1 MEM_stage_inst_dmem_U20041 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n20469), .ZN(MEM_stage_inst_dmem_n20452) );
NAND2_X1 MEM_stage_inst_dmem_U20040 ( .A1(MEM_stage_inst_dmem_ram_4056), .A2(MEM_stage_inst_dmem_n20468), .ZN(MEM_stage_inst_dmem_n20453) );
NAND2_X1 MEM_stage_inst_dmem_U20039 ( .A1(MEM_stage_inst_dmem_n20451), .A2(MEM_stage_inst_dmem_n20450), .ZN(MEM_stage_inst_dmem_n9236) );
NAND2_X1 MEM_stage_inst_dmem_U20038 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n20469), .ZN(MEM_stage_inst_dmem_n20450) );
NAND2_X1 MEM_stage_inst_dmem_U20037 ( .A1(MEM_stage_inst_dmem_ram_4057), .A2(MEM_stage_inst_dmem_n20468), .ZN(MEM_stage_inst_dmem_n20451) );
NAND2_X1 MEM_stage_inst_dmem_U20036 ( .A1(MEM_stage_inst_dmem_n20449), .A2(MEM_stage_inst_dmem_n20448), .ZN(MEM_stage_inst_dmem_n9237) );
NAND2_X1 MEM_stage_inst_dmem_U20035 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n20469), .ZN(MEM_stage_inst_dmem_n20448) );
NAND2_X1 MEM_stage_inst_dmem_U20034 ( .A1(MEM_stage_inst_dmem_ram_4058), .A2(MEM_stage_inst_dmem_n20468), .ZN(MEM_stage_inst_dmem_n20449) );
NAND2_X1 MEM_stage_inst_dmem_U20033 ( .A1(MEM_stage_inst_dmem_n20447), .A2(MEM_stage_inst_dmem_n20446), .ZN(MEM_stage_inst_dmem_n9238) );
NAND2_X1 MEM_stage_inst_dmem_U20032 ( .A1(MEM_stage_inst_dmem_n18004), .A2(MEM_stage_inst_dmem_n20469), .ZN(MEM_stage_inst_dmem_n20446) );
NAND2_X1 MEM_stage_inst_dmem_U20031 ( .A1(MEM_stage_inst_dmem_ram_4059), .A2(MEM_stage_inst_dmem_n20468), .ZN(MEM_stage_inst_dmem_n20447) );
NAND2_X1 MEM_stage_inst_dmem_U20030 ( .A1(MEM_stage_inst_dmem_n20445), .A2(MEM_stage_inst_dmem_n20444), .ZN(MEM_stage_inst_dmem_n9239) );
NAND2_X1 MEM_stage_inst_dmem_U20029 ( .A1(MEM_stage_inst_dmem_n18001), .A2(MEM_stage_inst_dmem_n20469), .ZN(MEM_stage_inst_dmem_n20444) );
NAND2_X1 MEM_stage_inst_dmem_U20028 ( .A1(MEM_stage_inst_dmem_ram_4060), .A2(MEM_stage_inst_dmem_n20468), .ZN(MEM_stage_inst_dmem_n20445) );
NAND2_X1 MEM_stage_inst_dmem_U20027 ( .A1(MEM_stage_inst_dmem_n20443), .A2(MEM_stage_inst_dmem_n20442), .ZN(MEM_stage_inst_dmem_n9240) );
NAND2_X1 MEM_stage_inst_dmem_U20026 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n20469), .ZN(MEM_stage_inst_dmem_n20442) );
NAND2_X1 MEM_stage_inst_dmem_U20025 ( .A1(MEM_stage_inst_dmem_ram_4061), .A2(MEM_stage_inst_dmem_n20468), .ZN(MEM_stage_inst_dmem_n20443) );
NAND2_X1 MEM_stage_inst_dmem_U20024 ( .A1(MEM_stage_inst_dmem_n20441), .A2(MEM_stage_inst_dmem_n20440), .ZN(MEM_stage_inst_dmem_n9241) );
NAND2_X1 MEM_stage_inst_dmem_U20023 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n20469), .ZN(MEM_stage_inst_dmem_n20440) );
NAND2_X1 MEM_stage_inst_dmem_U20022 ( .A1(MEM_stage_inst_dmem_ram_4062), .A2(MEM_stage_inst_dmem_n20468), .ZN(MEM_stage_inst_dmem_n20441) );
NAND2_X1 MEM_stage_inst_dmem_U20021 ( .A1(MEM_stage_inst_dmem_n20439), .A2(MEM_stage_inst_dmem_n20438), .ZN(MEM_stage_inst_dmem_n9242) );
NAND2_X1 MEM_stage_inst_dmem_U20020 ( .A1(MEM_stage_inst_dmem_n14693), .A2(MEM_stage_inst_dmem_n20469), .ZN(MEM_stage_inst_dmem_n20438) );
INV_X1 MEM_stage_inst_dmem_U20019 ( .A(MEM_stage_inst_dmem_n20468), .ZN(MEM_stage_inst_dmem_n20469) );
NAND2_X1 MEM_stage_inst_dmem_U20018 ( .A1(MEM_stage_inst_dmem_ram_4063), .A2(MEM_stage_inst_dmem_n20468), .ZN(MEM_stage_inst_dmem_n20439) );
NAND2_X1 MEM_stage_inst_dmem_U20017 ( .A1(MEM_stage_inst_dmem_n21004), .A2(MEM_stage_inst_dmem_n20895), .ZN(MEM_stage_inst_dmem_n20468) );
NAND2_X1 MEM_stage_inst_dmem_U20016 ( .A1(MEM_stage_inst_dmem_n20437), .A2(MEM_stage_inst_dmem_n20436), .ZN(MEM_stage_inst_dmem_n9243) );
NAND2_X1 MEM_stage_inst_dmem_U20015 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n20435), .ZN(MEM_stage_inst_dmem_n20436) );
NAND2_X1 MEM_stage_inst_dmem_U20014 ( .A1(MEM_stage_inst_dmem_ram_4064), .A2(MEM_stage_inst_dmem_n20434), .ZN(MEM_stage_inst_dmem_n20437) );
NAND2_X1 MEM_stage_inst_dmem_U20013 ( .A1(MEM_stage_inst_dmem_n20433), .A2(MEM_stage_inst_dmem_n20432), .ZN(MEM_stage_inst_dmem_n9244) );
NAND2_X1 MEM_stage_inst_dmem_U20012 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n20435), .ZN(MEM_stage_inst_dmem_n20432) );
NAND2_X1 MEM_stage_inst_dmem_U20011 ( .A1(MEM_stage_inst_dmem_ram_4065), .A2(MEM_stage_inst_dmem_n20434), .ZN(MEM_stage_inst_dmem_n20433) );
NAND2_X1 MEM_stage_inst_dmem_U20010 ( .A1(MEM_stage_inst_dmem_n20431), .A2(MEM_stage_inst_dmem_n20430), .ZN(MEM_stage_inst_dmem_n9245) );
NAND2_X1 MEM_stage_inst_dmem_U20009 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n20435), .ZN(MEM_stage_inst_dmem_n20430) );
NAND2_X1 MEM_stage_inst_dmem_U20008 ( .A1(MEM_stage_inst_dmem_ram_4066), .A2(MEM_stage_inst_dmem_n20434), .ZN(MEM_stage_inst_dmem_n20431) );
NAND2_X1 MEM_stage_inst_dmem_U20007 ( .A1(MEM_stage_inst_dmem_n20429), .A2(MEM_stage_inst_dmem_n20428), .ZN(MEM_stage_inst_dmem_n9246) );
NAND2_X1 MEM_stage_inst_dmem_U20006 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n20435), .ZN(MEM_stage_inst_dmem_n20428) );
NAND2_X1 MEM_stage_inst_dmem_U20005 ( .A1(MEM_stage_inst_dmem_ram_4067), .A2(MEM_stage_inst_dmem_n20434), .ZN(MEM_stage_inst_dmem_n20429) );
NAND2_X1 MEM_stage_inst_dmem_U20004 ( .A1(MEM_stage_inst_dmem_n20427), .A2(MEM_stage_inst_dmem_n20426), .ZN(MEM_stage_inst_dmem_n9247) );
NAND2_X1 MEM_stage_inst_dmem_U20003 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n20435), .ZN(MEM_stage_inst_dmem_n20426) );
NAND2_X1 MEM_stage_inst_dmem_U20002 ( .A1(MEM_stage_inst_dmem_ram_4068), .A2(MEM_stage_inst_dmem_n20434), .ZN(MEM_stage_inst_dmem_n20427) );
NAND2_X1 MEM_stage_inst_dmem_U20001 ( .A1(MEM_stage_inst_dmem_n20425), .A2(MEM_stage_inst_dmem_n20424), .ZN(MEM_stage_inst_dmem_n9248) );
NAND2_X1 MEM_stage_inst_dmem_U20000 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n20435), .ZN(MEM_stage_inst_dmem_n20424) );
NAND2_X1 MEM_stage_inst_dmem_U19999 ( .A1(MEM_stage_inst_dmem_ram_4069), .A2(MEM_stage_inst_dmem_n20434), .ZN(MEM_stage_inst_dmem_n20425) );
NAND2_X1 MEM_stage_inst_dmem_U19998 ( .A1(MEM_stage_inst_dmem_n20423), .A2(MEM_stage_inst_dmem_n20422), .ZN(MEM_stage_inst_dmem_n9249) );
NAND2_X1 MEM_stage_inst_dmem_U19997 ( .A1(MEM_stage_inst_dmem_n21340), .A2(MEM_stage_inst_dmem_n20435), .ZN(MEM_stage_inst_dmem_n20422) );
NAND2_X1 MEM_stage_inst_dmem_U19996 ( .A1(MEM_stage_inst_dmem_ram_4070), .A2(MEM_stage_inst_dmem_n20434), .ZN(MEM_stage_inst_dmem_n20423) );
NAND2_X1 MEM_stage_inst_dmem_U19995 ( .A1(MEM_stage_inst_dmem_n20421), .A2(MEM_stage_inst_dmem_n20420), .ZN(MEM_stage_inst_dmem_n9250) );
NAND2_X1 MEM_stage_inst_dmem_U19994 ( .A1(MEM_stage_inst_dmem_n18875), .A2(MEM_stage_inst_dmem_n20435), .ZN(MEM_stage_inst_dmem_n20420) );
NAND2_X1 MEM_stage_inst_dmem_U19993 ( .A1(MEM_stage_inst_dmem_ram_4071), .A2(MEM_stage_inst_dmem_n20434), .ZN(MEM_stage_inst_dmem_n20421) );
NAND2_X1 MEM_stage_inst_dmem_U19992 ( .A1(MEM_stage_inst_dmem_n20419), .A2(MEM_stage_inst_dmem_n20418), .ZN(MEM_stage_inst_dmem_n9251) );
NAND2_X1 MEM_stage_inst_dmem_U19991 ( .A1(MEM_stage_inst_dmem_n21335), .A2(MEM_stage_inst_dmem_n20435), .ZN(MEM_stage_inst_dmem_n20418) );
NAND2_X1 MEM_stage_inst_dmem_U19990 ( .A1(MEM_stage_inst_dmem_ram_4072), .A2(MEM_stage_inst_dmem_n20434), .ZN(MEM_stage_inst_dmem_n20419) );
NAND2_X1 MEM_stage_inst_dmem_U19989 ( .A1(MEM_stage_inst_dmem_n20417), .A2(MEM_stage_inst_dmem_n20416), .ZN(MEM_stage_inst_dmem_n9252) );
NAND2_X1 MEM_stage_inst_dmem_U19988 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n20435), .ZN(MEM_stage_inst_dmem_n20416) );
NAND2_X1 MEM_stage_inst_dmem_U19987 ( .A1(MEM_stage_inst_dmem_ram_4073), .A2(MEM_stage_inst_dmem_n20434), .ZN(MEM_stage_inst_dmem_n20417) );
NAND2_X1 MEM_stage_inst_dmem_U19986 ( .A1(MEM_stage_inst_dmem_n20415), .A2(MEM_stage_inst_dmem_n20414), .ZN(MEM_stage_inst_dmem_n9253) );
NAND2_X1 MEM_stage_inst_dmem_U19985 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n20435), .ZN(MEM_stage_inst_dmem_n20414) );
NAND2_X1 MEM_stage_inst_dmem_U19984 ( .A1(MEM_stage_inst_dmem_ram_4074), .A2(MEM_stage_inst_dmem_n20434), .ZN(MEM_stage_inst_dmem_n20415) );
NAND2_X1 MEM_stage_inst_dmem_U19983 ( .A1(MEM_stage_inst_dmem_n20413), .A2(MEM_stage_inst_dmem_n20412), .ZN(MEM_stage_inst_dmem_n9254) );
NAND2_X1 MEM_stage_inst_dmem_U19982 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n20435), .ZN(MEM_stage_inst_dmem_n20412) );
NAND2_X1 MEM_stage_inst_dmem_U19981 ( .A1(MEM_stage_inst_dmem_ram_4075), .A2(MEM_stage_inst_dmem_n20434), .ZN(MEM_stage_inst_dmem_n20413) );
NAND2_X1 MEM_stage_inst_dmem_U19980 ( .A1(MEM_stage_inst_dmem_n20411), .A2(MEM_stage_inst_dmem_n20410), .ZN(MEM_stage_inst_dmem_n9255) );
NAND2_X1 MEM_stage_inst_dmem_U19979 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n20435), .ZN(MEM_stage_inst_dmem_n20410) );
NAND2_X1 MEM_stage_inst_dmem_U19978 ( .A1(MEM_stage_inst_dmem_ram_4076), .A2(MEM_stage_inst_dmem_n20434), .ZN(MEM_stage_inst_dmem_n20411) );
NAND2_X1 MEM_stage_inst_dmem_U19977 ( .A1(MEM_stage_inst_dmem_n20409), .A2(MEM_stage_inst_dmem_n20408), .ZN(MEM_stage_inst_dmem_n9256) );
NAND2_X1 MEM_stage_inst_dmem_U19976 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n20435), .ZN(MEM_stage_inst_dmem_n20408) );
NAND2_X1 MEM_stage_inst_dmem_U19975 ( .A1(MEM_stage_inst_dmem_ram_4077), .A2(MEM_stage_inst_dmem_n20434), .ZN(MEM_stage_inst_dmem_n20409) );
NAND2_X1 MEM_stage_inst_dmem_U19974 ( .A1(MEM_stage_inst_dmem_n20407), .A2(MEM_stage_inst_dmem_n20406), .ZN(MEM_stage_inst_dmem_n9257) );
NAND2_X1 MEM_stage_inst_dmem_U19973 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n20435), .ZN(MEM_stage_inst_dmem_n20406) );
NAND2_X1 MEM_stage_inst_dmem_U19972 ( .A1(MEM_stage_inst_dmem_ram_4078), .A2(MEM_stage_inst_dmem_n20434), .ZN(MEM_stage_inst_dmem_n20407) );
NAND2_X1 MEM_stage_inst_dmem_U19971 ( .A1(MEM_stage_inst_dmem_n20405), .A2(MEM_stage_inst_dmem_n20404), .ZN(MEM_stage_inst_dmem_n9258) );
NAND2_X1 MEM_stage_inst_dmem_U19970 ( .A1(MEM_stage_inst_dmem_n16343), .A2(MEM_stage_inst_dmem_n20435), .ZN(MEM_stage_inst_dmem_n20404) );
INV_X1 MEM_stage_inst_dmem_U19969 ( .A(MEM_stage_inst_dmem_n20434), .ZN(MEM_stage_inst_dmem_n20435) );
NAND2_X1 MEM_stage_inst_dmem_U19968 ( .A1(MEM_stage_inst_dmem_ram_4079), .A2(MEM_stage_inst_dmem_n20434), .ZN(MEM_stage_inst_dmem_n20405) );
NAND2_X1 MEM_stage_inst_dmem_U19967 ( .A1(MEM_stage_inst_dmem_n20969), .A2(MEM_stage_inst_dmem_n20895), .ZN(MEM_stage_inst_dmem_n20434) );
NAND2_X1 MEM_stage_inst_dmem_U19966 ( .A1(MEM_stage_inst_dmem_n20403), .A2(MEM_stage_inst_dmem_n20402), .ZN(MEM_stage_inst_dmem_n9259) );
NAND2_X1 MEM_stage_inst_dmem_U19965 ( .A1(MEM_stage_inst_dmem_n20551), .A2(MEM_stage_inst_dmem_n20401), .ZN(MEM_stage_inst_dmem_n20402) );
NAND2_X1 MEM_stage_inst_dmem_U19964 ( .A1(MEM_stage_inst_dmem_ram_4080), .A2(MEM_stage_inst_dmem_n20400), .ZN(MEM_stage_inst_dmem_n20403) );
NAND2_X1 MEM_stage_inst_dmem_U19963 ( .A1(MEM_stage_inst_dmem_n20399), .A2(MEM_stage_inst_dmem_n20398), .ZN(MEM_stage_inst_dmem_n9260) );
NAND2_X1 MEM_stage_inst_dmem_U19962 ( .A1(MEM_stage_inst_dmem_n20547), .A2(MEM_stage_inst_dmem_n20401), .ZN(MEM_stage_inst_dmem_n20398) );
NAND2_X1 MEM_stage_inst_dmem_U19961 ( .A1(MEM_stage_inst_dmem_ram_4081), .A2(MEM_stage_inst_dmem_n20400), .ZN(MEM_stage_inst_dmem_n20399) );
NAND2_X1 MEM_stage_inst_dmem_U19960 ( .A1(MEM_stage_inst_dmem_n20397), .A2(MEM_stage_inst_dmem_n20396), .ZN(MEM_stage_inst_dmem_n9261) );
NAND2_X1 MEM_stage_inst_dmem_U19959 ( .A1(MEM_stage_inst_dmem_n20544), .A2(MEM_stage_inst_dmem_n20401), .ZN(MEM_stage_inst_dmem_n20396) );
NAND2_X1 MEM_stage_inst_dmem_U19958 ( .A1(MEM_stage_inst_dmem_ram_4082), .A2(MEM_stage_inst_dmem_n20400), .ZN(MEM_stage_inst_dmem_n20397) );
NAND2_X1 MEM_stage_inst_dmem_U19957 ( .A1(MEM_stage_inst_dmem_n20395), .A2(MEM_stage_inst_dmem_n20394), .ZN(MEM_stage_inst_dmem_n9262) );
NAND2_X1 MEM_stage_inst_dmem_U19956 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n20401), .ZN(MEM_stage_inst_dmem_n20394) );
NAND2_X1 MEM_stage_inst_dmem_U19955 ( .A1(MEM_stage_inst_dmem_ram_4083), .A2(MEM_stage_inst_dmem_n20400), .ZN(MEM_stage_inst_dmem_n20395) );
NAND2_X1 MEM_stage_inst_dmem_U19954 ( .A1(MEM_stage_inst_dmem_n20393), .A2(MEM_stage_inst_dmem_n20392), .ZN(MEM_stage_inst_dmem_n9263) );
NAND2_X1 MEM_stage_inst_dmem_U19953 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n20401), .ZN(MEM_stage_inst_dmem_n20392) );
NAND2_X1 MEM_stage_inst_dmem_U19952 ( .A1(MEM_stage_inst_dmem_ram_4084), .A2(MEM_stage_inst_dmem_n20400), .ZN(MEM_stage_inst_dmem_n20393) );
NAND2_X1 MEM_stage_inst_dmem_U19951 ( .A1(MEM_stage_inst_dmem_n20391), .A2(MEM_stage_inst_dmem_n20390), .ZN(MEM_stage_inst_dmem_n9264) );
NAND2_X1 MEM_stage_inst_dmem_U19950 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n20401), .ZN(MEM_stage_inst_dmem_n20390) );
NAND2_X1 MEM_stage_inst_dmem_U19949 ( .A1(MEM_stage_inst_dmem_ram_4085), .A2(MEM_stage_inst_dmem_n20400), .ZN(MEM_stage_inst_dmem_n20391) );
NAND2_X1 MEM_stage_inst_dmem_U19948 ( .A1(MEM_stage_inst_dmem_n20389), .A2(MEM_stage_inst_dmem_n20388), .ZN(MEM_stage_inst_dmem_n9265) );
NAND2_X1 MEM_stage_inst_dmem_U19947 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n20401), .ZN(MEM_stage_inst_dmem_n20388) );
NAND2_X1 MEM_stage_inst_dmem_U19946 ( .A1(MEM_stage_inst_dmem_ram_4086), .A2(MEM_stage_inst_dmem_n20400), .ZN(MEM_stage_inst_dmem_n20389) );
NAND2_X1 MEM_stage_inst_dmem_U19945 ( .A1(MEM_stage_inst_dmem_n20387), .A2(MEM_stage_inst_dmem_n20386), .ZN(MEM_stage_inst_dmem_n9266) );
NAND2_X1 MEM_stage_inst_dmem_U19944 ( .A1(MEM_stage_inst_dmem_n20530), .A2(MEM_stage_inst_dmem_n20401), .ZN(MEM_stage_inst_dmem_n20386) );
NAND2_X1 MEM_stage_inst_dmem_U19943 ( .A1(MEM_stage_inst_dmem_ram_4087), .A2(MEM_stage_inst_dmem_n20400), .ZN(MEM_stage_inst_dmem_n20387) );
NAND2_X1 MEM_stage_inst_dmem_U19942 ( .A1(MEM_stage_inst_dmem_n20385), .A2(MEM_stage_inst_dmem_n20384), .ZN(MEM_stage_inst_dmem_n9267) );
NAND2_X1 MEM_stage_inst_dmem_U19941 ( .A1(MEM_stage_inst_dmem_n20527), .A2(MEM_stage_inst_dmem_n20401), .ZN(MEM_stage_inst_dmem_n20384) );
NAND2_X1 MEM_stage_inst_dmem_U19940 ( .A1(MEM_stage_inst_dmem_ram_4088), .A2(MEM_stage_inst_dmem_n20400), .ZN(MEM_stage_inst_dmem_n20385) );
NAND2_X1 MEM_stage_inst_dmem_U19939 ( .A1(MEM_stage_inst_dmem_n20383), .A2(MEM_stage_inst_dmem_n20382), .ZN(MEM_stage_inst_dmem_n9268) );
NAND2_X1 MEM_stage_inst_dmem_U19938 ( .A1(MEM_stage_inst_dmem_n20524), .A2(MEM_stage_inst_dmem_n20401), .ZN(MEM_stage_inst_dmem_n20382) );
NAND2_X1 MEM_stage_inst_dmem_U19937 ( .A1(MEM_stage_inst_dmem_ram_4089), .A2(MEM_stage_inst_dmem_n20400), .ZN(MEM_stage_inst_dmem_n20383) );
NAND2_X1 MEM_stage_inst_dmem_U19936 ( .A1(MEM_stage_inst_dmem_n20381), .A2(MEM_stage_inst_dmem_n20380), .ZN(MEM_stage_inst_dmem_n9269) );
NAND2_X1 MEM_stage_inst_dmem_U19935 ( .A1(MEM_stage_inst_dmem_n20521), .A2(MEM_stage_inst_dmem_n20401), .ZN(MEM_stage_inst_dmem_n20380) );
NAND2_X1 MEM_stage_inst_dmem_U19934 ( .A1(MEM_stage_inst_dmem_ram_4090), .A2(MEM_stage_inst_dmem_n20400), .ZN(MEM_stage_inst_dmem_n20381) );
NAND2_X1 MEM_stage_inst_dmem_U19933 ( .A1(MEM_stage_inst_dmem_n20379), .A2(MEM_stage_inst_dmem_n20378), .ZN(MEM_stage_inst_dmem_n9270) );
NAND2_X1 MEM_stage_inst_dmem_U19932 ( .A1(MEM_stage_inst_dmem_n20518), .A2(MEM_stage_inst_dmem_n20401), .ZN(MEM_stage_inst_dmem_n20378) );
NAND2_X1 MEM_stage_inst_dmem_U19931 ( .A1(MEM_stage_inst_dmem_ram_4091), .A2(MEM_stage_inst_dmem_n20400), .ZN(MEM_stage_inst_dmem_n20379) );
NAND2_X1 MEM_stage_inst_dmem_U19930 ( .A1(MEM_stage_inst_dmem_n20377), .A2(MEM_stage_inst_dmem_n20376), .ZN(MEM_stage_inst_dmem_n9271) );
NAND2_X1 MEM_stage_inst_dmem_U19929 ( .A1(MEM_stage_inst_dmem_n20515), .A2(MEM_stage_inst_dmem_n20401), .ZN(MEM_stage_inst_dmem_n20376) );
NAND2_X1 MEM_stage_inst_dmem_U19928 ( .A1(MEM_stage_inst_dmem_ram_4092), .A2(MEM_stage_inst_dmem_n20400), .ZN(MEM_stage_inst_dmem_n20377) );
NAND2_X1 MEM_stage_inst_dmem_U19927 ( .A1(MEM_stage_inst_dmem_n20375), .A2(MEM_stage_inst_dmem_n20374), .ZN(MEM_stage_inst_dmem_n9272) );
NAND2_X1 MEM_stage_inst_dmem_U19926 ( .A1(MEM_stage_inst_dmem_n20512), .A2(MEM_stage_inst_dmem_n20401), .ZN(MEM_stage_inst_dmem_n20374) );
NAND2_X1 MEM_stage_inst_dmem_U19925 ( .A1(MEM_stage_inst_dmem_ram_4093), .A2(MEM_stage_inst_dmem_n20400), .ZN(MEM_stage_inst_dmem_n20375) );
NAND2_X1 MEM_stage_inst_dmem_U19924 ( .A1(MEM_stage_inst_dmem_n20373), .A2(MEM_stage_inst_dmem_n20372), .ZN(MEM_stage_inst_dmem_n9273) );
NAND2_X1 MEM_stage_inst_dmem_U19923 ( .A1(MEM_stage_inst_dmem_n20509), .A2(MEM_stage_inst_dmem_n20401), .ZN(MEM_stage_inst_dmem_n20372) );
NAND2_X1 MEM_stage_inst_dmem_U19922 ( .A1(MEM_stage_inst_dmem_ram_4094), .A2(MEM_stage_inst_dmem_n20400), .ZN(MEM_stage_inst_dmem_n20373) );
NAND2_X1 MEM_stage_inst_dmem_U19921 ( .A1(MEM_stage_inst_dmem_n20371), .A2(MEM_stage_inst_dmem_n20370), .ZN(MEM_stage_inst_dmem_n9274) );
NAND2_X1 MEM_stage_inst_dmem_U19920 ( .A1(MEM_stage_inst_dmem_n20506), .A2(MEM_stage_inst_dmem_n20401), .ZN(MEM_stage_inst_dmem_n20370) );
INV_X1 MEM_stage_inst_dmem_U19919 ( .A(MEM_stage_inst_dmem_n20400), .ZN(MEM_stage_inst_dmem_n20401) );
NAND2_X1 MEM_stage_inst_dmem_U19918 ( .A1(MEM_stage_inst_dmem_ram_4095), .A2(MEM_stage_inst_dmem_n20400), .ZN(MEM_stage_inst_dmem_n20371) );
NAND2_X1 MEM_stage_inst_dmem_U19917 ( .A1(MEM_stage_inst_dmem_n20934), .A2(MEM_stage_inst_dmem_n20895), .ZN(MEM_stage_inst_dmem_n20400) );
NOR2_X2 MEM_stage_inst_dmem_U19916 ( .A1(MEM_stage_inst_dmem_n20933), .A2(MEM_stage_inst_dmem_n20369), .ZN(MEM_stage_inst_dmem_n20895) );
NAND2_X1 MEM_stage_inst_dmem_U19915 ( .A1(MEM_stage_inst_dmem_n20368), .A2(MEM_stage_inst_dmem_n20367), .ZN(MEM_stage_inst_dmem_n9275) );
NAND2_X1 MEM_stage_inst_dmem_U19914 ( .A1(MEM_stage_inst_dmem_n20551), .A2(MEM_stage_inst_dmem_n20366), .ZN(MEM_stage_inst_dmem_n20367) );
NAND2_X1 MEM_stage_inst_dmem_U19913 ( .A1(MEM_stage_inst_dmem_ram_3072), .A2(MEM_stage_inst_dmem_n20365), .ZN(MEM_stage_inst_dmem_n20368) );
NAND2_X1 MEM_stage_inst_dmem_U19912 ( .A1(MEM_stage_inst_dmem_n20364), .A2(MEM_stage_inst_dmem_n20363), .ZN(MEM_stage_inst_dmem_n9276) );
NAND2_X1 MEM_stage_inst_dmem_U19911 ( .A1(MEM_stage_inst_dmem_n20547), .A2(MEM_stage_inst_dmem_n20366), .ZN(MEM_stage_inst_dmem_n20363) );
NAND2_X1 MEM_stage_inst_dmem_U19910 ( .A1(MEM_stage_inst_dmem_ram_3073), .A2(MEM_stage_inst_dmem_n20365), .ZN(MEM_stage_inst_dmem_n20364) );
NAND2_X1 MEM_stage_inst_dmem_U19909 ( .A1(MEM_stage_inst_dmem_n20362), .A2(MEM_stage_inst_dmem_n20361), .ZN(MEM_stage_inst_dmem_n9277) );
NAND2_X1 MEM_stage_inst_dmem_U19908 ( .A1(MEM_stage_inst_dmem_n20544), .A2(MEM_stage_inst_dmem_n20366), .ZN(MEM_stage_inst_dmem_n20361) );
NAND2_X1 MEM_stage_inst_dmem_U19907 ( .A1(MEM_stage_inst_dmem_ram_3074), .A2(MEM_stage_inst_dmem_n20365), .ZN(MEM_stage_inst_dmem_n20362) );
NAND2_X1 MEM_stage_inst_dmem_U19906 ( .A1(MEM_stage_inst_dmem_n20360), .A2(MEM_stage_inst_dmem_n20359), .ZN(MEM_stage_inst_dmem_n9278) );
NAND2_X1 MEM_stage_inst_dmem_U19905 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n20366), .ZN(MEM_stage_inst_dmem_n20359) );
NAND2_X1 MEM_stage_inst_dmem_U19904 ( .A1(MEM_stage_inst_dmem_ram_3075), .A2(MEM_stage_inst_dmem_n20365), .ZN(MEM_stage_inst_dmem_n20360) );
NAND2_X1 MEM_stage_inst_dmem_U19903 ( .A1(MEM_stage_inst_dmem_n20358), .A2(MEM_stage_inst_dmem_n20357), .ZN(MEM_stage_inst_dmem_n9279) );
NAND2_X1 MEM_stage_inst_dmem_U19902 ( .A1(EX_pipeline_reg_out_9), .A2(MEM_stage_inst_dmem_n20366), .ZN(MEM_stage_inst_dmem_n20357) );
NAND2_X1 MEM_stage_inst_dmem_U19901 ( .A1(MEM_stage_inst_dmem_ram_3076), .A2(MEM_stage_inst_dmem_n20365), .ZN(MEM_stage_inst_dmem_n20358) );
NAND2_X1 MEM_stage_inst_dmem_U19900 ( .A1(MEM_stage_inst_dmem_n20356), .A2(MEM_stage_inst_dmem_n20355), .ZN(MEM_stage_inst_dmem_n9280) );
NAND2_X1 MEM_stage_inst_dmem_U19899 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n20366), .ZN(MEM_stage_inst_dmem_n20355) );
NAND2_X1 MEM_stage_inst_dmem_U19898 ( .A1(MEM_stage_inst_dmem_ram_3077), .A2(MEM_stage_inst_dmem_n20365), .ZN(MEM_stage_inst_dmem_n20356) );
NAND2_X1 MEM_stage_inst_dmem_U19897 ( .A1(MEM_stage_inst_dmem_n20354), .A2(MEM_stage_inst_dmem_n20353), .ZN(MEM_stage_inst_dmem_n9281) );
NAND2_X1 MEM_stage_inst_dmem_U19896 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n20366), .ZN(MEM_stage_inst_dmem_n20353) );
NAND2_X1 MEM_stage_inst_dmem_U19895 ( .A1(MEM_stage_inst_dmem_ram_3078), .A2(MEM_stage_inst_dmem_n20365), .ZN(MEM_stage_inst_dmem_n20354) );
NAND2_X1 MEM_stage_inst_dmem_U19894 ( .A1(MEM_stage_inst_dmem_n20352), .A2(MEM_stage_inst_dmem_n20351), .ZN(MEM_stage_inst_dmem_n9282) );
NAND2_X1 MEM_stage_inst_dmem_U19893 ( .A1(MEM_stage_inst_dmem_n20530), .A2(MEM_stage_inst_dmem_n20366), .ZN(MEM_stage_inst_dmem_n20351) );
NAND2_X1 MEM_stage_inst_dmem_U19892 ( .A1(MEM_stage_inst_dmem_ram_3079), .A2(MEM_stage_inst_dmem_n20365), .ZN(MEM_stage_inst_dmem_n20352) );
NAND2_X1 MEM_stage_inst_dmem_U19891 ( .A1(MEM_stage_inst_dmem_n20350), .A2(MEM_stage_inst_dmem_n20349), .ZN(MEM_stage_inst_dmem_n9283) );
NAND2_X1 MEM_stage_inst_dmem_U19890 ( .A1(MEM_stage_inst_dmem_n20527), .A2(MEM_stage_inst_dmem_n20366), .ZN(MEM_stage_inst_dmem_n20349) );
NAND2_X1 MEM_stage_inst_dmem_U19889 ( .A1(MEM_stage_inst_dmem_ram_3080), .A2(MEM_stage_inst_dmem_n20365), .ZN(MEM_stage_inst_dmem_n20350) );
NAND2_X1 MEM_stage_inst_dmem_U19888 ( .A1(MEM_stage_inst_dmem_n20348), .A2(MEM_stage_inst_dmem_n20347), .ZN(MEM_stage_inst_dmem_n9284) );
NAND2_X1 MEM_stage_inst_dmem_U19887 ( .A1(MEM_stage_inst_dmem_n20524), .A2(MEM_stage_inst_dmem_n20366), .ZN(MEM_stage_inst_dmem_n20347) );
NAND2_X1 MEM_stage_inst_dmem_U19886 ( .A1(MEM_stage_inst_dmem_ram_3081), .A2(MEM_stage_inst_dmem_n20365), .ZN(MEM_stage_inst_dmem_n20348) );
NAND2_X1 MEM_stage_inst_dmem_U19885 ( .A1(MEM_stage_inst_dmem_n20346), .A2(MEM_stage_inst_dmem_n20345), .ZN(MEM_stage_inst_dmem_n9285) );
NAND2_X1 MEM_stage_inst_dmem_U19884 ( .A1(MEM_stage_inst_dmem_n20521), .A2(MEM_stage_inst_dmem_n20366), .ZN(MEM_stage_inst_dmem_n20345) );
NAND2_X1 MEM_stage_inst_dmem_U19883 ( .A1(MEM_stage_inst_dmem_ram_3082), .A2(MEM_stage_inst_dmem_n20365), .ZN(MEM_stage_inst_dmem_n20346) );
NAND2_X1 MEM_stage_inst_dmem_U19882 ( .A1(MEM_stage_inst_dmem_n20344), .A2(MEM_stage_inst_dmem_n20343), .ZN(MEM_stage_inst_dmem_n9286) );
NAND2_X1 MEM_stage_inst_dmem_U19881 ( .A1(MEM_stage_inst_dmem_n20518), .A2(MEM_stage_inst_dmem_n20366), .ZN(MEM_stage_inst_dmem_n20343) );
NAND2_X1 MEM_stage_inst_dmem_U19880 ( .A1(MEM_stage_inst_dmem_ram_3083), .A2(MEM_stage_inst_dmem_n20365), .ZN(MEM_stage_inst_dmem_n20344) );
NAND2_X1 MEM_stage_inst_dmem_U19879 ( .A1(MEM_stage_inst_dmem_n20342), .A2(MEM_stage_inst_dmem_n20341), .ZN(MEM_stage_inst_dmem_n9287) );
NAND2_X1 MEM_stage_inst_dmem_U19878 ( .A1(MEM_stage_inst_dmem_n20515), .A2(MEM_stage_inst_dmem_n20366), .ZN(MEM_stage_inst_dmem_n20341) );
NAND2_X1 MEM_stage_inst_dmem_U19877 ( .A1(MEM_stage_inst_dmem_ram_3084), .A2(MEM_stage_inst_dmem_n20365), .ZN(MEM_stage_inst_dmem_n20342) );
NAND2_X1 MEM_stage_inst_dmem_U19876 ( .A1(MEM_stage_inst_dmem_n20340), .A2(MEM_stage_inst_dmem_n20339), .ZN(MEM_stage_inst_dmem_n9288) );
NAND2_X1 MEM_stage_inst_dmem_U19875 ( .A1(MEM_stage_inst_dmem_n20512), .A2(MEM_stage_inst_dmem_n20366), .ZN(MEM_stage_inst_dmem_n20339) );
NAND2_X1 MEM_stage_inst_dmem_U19874 ( .A1(MEM_stage_inst_dmem_ram_3085), .A2(MEM_stage_inst_dmem_n20365), .ZN(MEM_stage_inst_dmem_n20340) );
NAND2_X1 MEM_stage_inst_dmem_U19873 ( .A1(MEM_stage_inst_dmem_n20338), .A2(MEM_stage_inst_dmem_n20337), .ZN(MEM_stage_inst_dmem_n9289) );
NAND2_X1 MEM_stage_inst_dmem_U19872 ( .A1(MEM_stage_inst_dmem_n20509), .A2(MEM_stage_inst_dmem_n20366), .ZN(MEM_stage_inst_dmem_n20337) );
NAND2_X1 MEM_stage_inst_dmem_U19871 ( .A1(MEM_stage_inst_dmem_ram_3086), .A2(MEM_stage_inst_dmem_n20365), .ZN(MEM_stage_inst_dmem_n20338) );
NAND2_X1 MEM_stage_inst_dmem_U19870 ( .A1(MEM_stage_inst_dmem_n20336), .A2(MEM_stage_inst_dmem_n20335), .ZN(MEM_stage_inst_dmem_n9290) );
NAND2_X1 MEM_stage_inst_dmem_U19869 ( .A1(MEM_stage_inst_dmem_n20506), .A2(MEM_stage_inst_dmem_n20366), .ZN(MEM_stage_inst_dmem_n20335) );
NAND2_X1 MEM_stage_inst_dmem_U19868 ( .A1(MEM_stage_inst_dmem_ram_3087), .A2(MEM_stage_inst_dmem_n20365), .ZN(MEM_stage_inst_dmem_n20336) );
NAND2_X1 MEM_stage_inst_dmem_U19867 ( .A1(MEM_stage_inst_dmem_n21465), .A2(MEM_stage_inst_dmem_n20334), .ZN(MEM_stage_inst_dmem_n20365) );
NAND2_X1 MEM_stage_inst_dmem_U19866 ( .A1(MEM_stage_inst_dmem_n20333), .A2(MEM_stage_inst_dmem_n20332), .ZN(MEM_stage_inst_dmem_n9291) );
NAND2_X1 MEM_stage_inst_dmem_U19865 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n20331), .ZN(MEM_stage_inst_dmem_n20332) );
NAND2_X1 MEM_stage_inst_dmem_U19864 ( .A1(MEM_stage_inst_dmem_ram_3088), .A2(MEM_stage_inst_dmem_n20330), .ZN(MEM_stage_inst_dmem_n20333) );
NAND2_X1 MEM_stage_inst_dmem_U19863 ( .A1(MEM_stage_inst_dmem_n20329), .A2(MEM_stage_inst_dmem_n20328), .ZN(MEM_stage_inst_dmem_n9292) );
NAND2_X1 MEM_stage_inst_dmem_U19862 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n20331), .ZN(MEM_stage_inst_dmem_n20328) );
NAND2_X1 MEM_stage_inst_dmem_U19861 ( .A1(MEM_stage_inst_dmem_ram_3089), .A2(MEM_stage_inst_dmem_n20330), .ZN(MEM_stage_inst_dmem_n20329) );
NAND2_X1 MEM_stage_inst_dmem_U19860 ( .A1(MEM_stage_inst_dmem_n20327), .A2(MEM_stage_inst_dmem_n20326), .ZN(MEM_stage_inst_dmem_n9293) );
NAND2_X1 MEM_stage_inst_dmem_U19859 ( .A1(MEM_stage_inst_dmem_n20544), .A2(MEM_stage_inst_dmem_n20331), .ZN(MEM_stage_inst_dmem_n20326) );
NAND2_X1 MEM_stage_inst_dmem_U19858 ( .A1(MEM_stage_inst_dmem_ram_3090), .A2(MEM_stage_inst_dmem_n20330), .ZN(MEM_stage_inst_dmem_n20327) );
NAND2_X1 MEM_stage_inst_dmem_U19857 ( .A1(MEM_stage_inst_dmem_n20325), .A2(MEM_stage_inst_dmem_n20324), .ZN(MEM_stage_inst_dmem_n9294) );
NAND2_X1 MEM_stage_inst_dmem_U19856 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n20331), .ZN(MEM_stage_inst_dmem_n20324) );
NAND2_X1 MEM_stage_inst_dmem_U19855 ( .A1(MEM_stage_inst_dmem_ram_3091), .A2(MEM_stage_inst_dmem_n20330), .ZN(MEM_stage_inst_dmem_n20325) );
NAND2_X1 MEM_stage_inst_dmem_U19854 ( .A1(MEM_stage_inst_dmem_n20323), .A2(MEM_stage_inst_dmem_n20322), .ZN(MEM_stage_inst_dmem_n9295) );
NAND2_X1 MEM_stage_inst_dmem_U19853 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n20331), .ZN(MEM_stage_inst_dmem_n20322) );
NAND2_X1 MEM_stage_inst_dmem_U19852 ( .A1(MEM_stage_inst_dmem_ram_3092), .A2(MEM_stage_inst_dmem_n20330), .ZN(MEM_stage_inst_dmem_n20323) );
NAND2_X1 MEM_stage_inst_dmem_U19851 ( .A1(MEM_stage_inst_dmem_n20321), .A2(MEM_stage_inst_dmem_n20320), .ZN(MEM_stage_inst_dmem_n9296) );
NAND2_X1 MEM_stage_inst_dmem_U19850 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n20331), .ZN(MEM_stage_inst_dmem_n20320) );
NAND2_X1 MEM_stage_inst_dmem_U19849 ( .A1(MEM_stage_inst_dmem_ram_3093), .A2(MEM_stage_inst_dmem_n20330), .ZN(MEM_stage_inst_dmem_n20321) );
NAND2_X1 MEM_stage_inst_dmem_U19848 ( .A1(MEM_stage_inst_dmem_n20319), .A2(MEM_stage_inst_dmem_n20318), .ZN(MEM_stage_inst_dmem_n9297) );
NAND2_X1 MEM_stage_inst_dmem_U19847 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n20331), .ZN(MEM_stage_inst_dmem_n20318) );
NAND2_X1 MEM_stage_inst_dmem_U19846 ( .A1(MEM_stage_inst_dmem_ram_3094), .A2(MEM_stage_inst_dmem_n20330), .ZN(MEM_stage_inst_dmem_n20319) );
NAND2_X1 MEM_stage_inst_dmem_U19845 ( .A1(MEM_stage_inst_dmem_n20317), .A2(MEM_stage_inst_dmem_n20316), .ZN(MEM_stage_inst_dmem_n9298) );
NAND2_X1 MEM_stage_inst_dmem_U19844 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n20331), .ZN(MEM_stage_inst_dmem_n20316) );
NAND2_X1 MEM_stage_inst_dmem_U19843 ( .A1(MEM_stage_inst_dmem_ram_3095), .A2(MEM_stage_inst_dmem_n20330), .ZN(MEM_stage_inst_dmem_n20317) );
NAND2_X1 MEM_stage_inst_dmem_U19842 ( .A1(MEM_stage_inst_dmem_n20315), .A2(MEM_stage_inst_dmem_n20314), .ZN(MEM_stage_inst_dmem_n9299) );
NAND2_X1 MEM_stage_inst_dmem_U19841 ( .A1(MEM_stage_inst_dmem_n13051), .A2(MEM_stage_inst_dmem_n20331), .ZN(MEM_stage_inst_dmem_n20314) );
NAND2_X1 MEM_stage_inst_dmem_U19840 ( .A1(MEM_stage_inst_dmem_ram_3096), .A2(MEM_stage_inst_dmem_n20330), .ZN(MEM_stage_inst_dmem_n20315) );
NAND2_X1 MEM_stage_inst_dmem_U19839 ( .A1(MEM_stage_inst_dmem_n20313), .A2(MEM_stage_inst_dmem_n20312), .ZN(MEM_stage_inst_dmem_n9300) );
NAND2_X1 MEM_stage_inst_dmem_U19838 ( .A1(MEM_stage_inst_dmem_n19251), .A2(MEM_stage_inst_dmem_n20331), .ZN(MEM_stage_inst_dmem_n20312) );
NAND2_X1 MEM_stage_inst_dmem_U19837 ( .A1(MEM_stage_inst_dmem_ram_3097), .A2(MEM_stage_inst_dmem_n20330), .ZN(MEM_stage_inst_dmem_n20313) );
NAND2_X1 MEM_stage_inst_dmem_U19836 ( .A1(MEM_stage_inst_dmem_n20311), .A2(MEM_stage_inst_dmem_n20310), .ZN(MEM_stage_inst_dmem_n9301) );
NAND2_X1 MEM_stage_inst_dmem_U19835 ( .A1(MEM_stage_inst_dmem_n20521), .A2(MEM_stage_inst_dmem_n20331), .ZN(MEM_stage_inst_dmem_n20310) );
NAND2_X1 MEM_stage_inst_dmem_U19834 ( .A1(MEM_stage_inst_dmem_ram_3098), .A2(MEM_stage_inst_dmem_n20330), .ZN(MEM_stage_inst_dmem_n20311) );
NAND2_X1 MEM_stage_inst_dmem_U19833 ( .A1(MEM_stage_inst_dmem_n20309), .A2(MEM_stage_inst_dmem_n20308), .ZN(MEM_stage_inst_dmem_n9302) );
NAND2_X1 MEM_stage_inst_dmem_U19832 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n20331), .ZN(MEM_stage_inst_dmem_n20308) );
NAND2_X1 MEM_stage_inst_dmem_U19831 ( .A1(MEM_stage_inst_dmem_ram_3099), .A2(MEM_stage_inst_dmem_n20330), .ZN(MEM_stage_inst_dmem_n20309) );
NAND2_X1 MEM_stage_inst_dmem_U19830 ( .A1(MEM_stage_inst_dmem_n20307), .A2(MEM_stage_inst_dmem_n20306), .ZN(MEM_stage_inst_dmem_n9303) );
NAND2_X1 MEM_stage_inst_dmem_U19829 ( .A1(MEM_stage_inst_dmem_n14702), .A2(MEM_stage_inst_dmem_n20331), .ZN(MEM_stage_inst_dmem_n20306) );
NAND2_X1 MEM_stage_inst_dmem_U19828 ( .A1(MEM_stage_inst_dmem_ram_3100), .A2(MEM_stage_inst_dmem_n20330), .ZN(MEM_stage_inst_dmem_n20307) );
NAND2_X1 MEM_stage_inst_dmem_U19827 ( .A1(MEM_stage_inst_dmem_n20305), .A2(MEM_stage_inst_dmem_n20304), .ZN(MEM_stage_inst_dmem_n9304) );
NAND2_X1 MEM_stage_inst_dmem_U19826 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n20331), .ZN(MEM_stage_inst_dmem_n20304) );
NAND2_X1 MEM_stage_inst_dmem_U19825 ( .A1(MEM_stage_inst_dmem_ram_3101), .A2(MEM_stage_inst_dmem_n20330), .ZN(MEM_stage_inst_dmem_n20305) );
NAND2_X1 MEM_stage_inst_dmem_U19824 ( .A1(MEM_stage_inst_dmem_n20303), .A2(MEM_stage_inst_dmem_n20302), .ZN(MEM_stage_inst_dmem_n9305) );
NAND2_X1 MEM_stage_inst_dmem_U19823 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n20331), .ZN(MEM_stage_inst_dmem_n20302) );
NAND2_X1 MEM_stage_inst_dmem_U19822 ( .A1(MEM_stage_inst_dmem_ram_3102), .A2(MEM_stage_inst_dmem_n20330), .ZN(MEM_stage_inst_dmem_n20303) );
NAND2_X1 MEM_stage_inst_dmem_U19821 ( .A1(MEM_stage_inst_dmem_n20301), .A2(MEM_stage_inst_dmem_n20300), .ZN(MEM_stage_inst_dmem_n9306) );
NAND2_X1 MEM_stage_inst_dmem_U19820 ( .A1(MEM_stage_inst_dmem_n21320), .A2(MEM_stage_inst_dmem_n20331), .ZN(MEM_stage_inst_dmem_n20300) );
INV_X1 MEM_stage_inst_dmem_U19819 ( .A(MEM_stage_inst_dmem_n20330), .ZN(MEM_stage_inst_dmem_n20331) );
NAND2_X1 MEM_stage_inst_dmem_U19818 ( .A1(MEM_stage_inst_dmem_ram_3103), .A2(MEM_stage_inst_dmem_n20330), .ZN(MEM_stage_inst_dmem_n20301) );
NAND2_X1 MEM_stage_inst_dmem_U19817 ( .A1(MEM_stage_inst_dmem_n21429), .A2(MEM_stage_inst_dmem_n20334), .ZN(MEM_stage_inst_dmem_n20330) );
NAND2_X1 MEM_stage_inst_dmem_U19816 ( .A1(MEM_stage_inst_dmem_n20299), .A2(MEM_stage_inst_dmem_n20298), .ZN(MEM_stage_inst_dmem_n9307) );
NAND2_X1 MEM_stage_inst_dmem_U19815 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n20297), .ZN(MEM_stage_inst_dmem_n20298) );
NAND2_X1 MEM_stage_inst_dmem_U19814 ( .A1(MEM_stage_inst_dmem_ram_3104), .A2(MEM_stage_inst_dmem_n20296), .ZN(MEM_stage_inst_dmem_n20299) );
NAND2_X1 MEM_stage_inst_dmem_U19813 ( .A1(MEM_stage_inst_dmem_n20295), .A2(MEM_stage_inst_dmem_n20294), .ZN(MEM_stage_inst_dmem_n9308) );
NAND2_X1 MEM_stage_inst_dmem_U19812 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n20297), .ZN(MEM_stage_inst_dmem_n20294) );
NAND2_X1 MEM_stage_inst_dmem_U19811 ( .A1(MEM_stage_inst_dmem_ram_3105), .A2(MEM_stage_inst_dmem_n20296), .ZN(MEM_stage_inst_dmem_n20295) );
NAND2_X1 MEM_stage_inst_dmem_U19810 ( .A1(MEM_stage_inst_dmem_n20293), .A2(MEM_stage_inst_dmem_n20292), .ZN(MEM_stage_inst_dmem_n9309) );
NAND2_X1 MEM_stage_inst_dmem_U19809 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n20297), .ZN(MEM_stage_inst_dmem_n20292) );
NAND2_X1 MEM_stage_inst_dmem_U19808 ( .A1(MEM_stage_inst_dmem_ram_3106), .A2(MEM_stage_inst_dmem_n20296), .ZN(MEM_stage_inst_dmem_n20293) );
NAND2_X1 MEM_stage_inst_dmem_U19807 ( .A1(MEM_stage_inst_dmem_n20291), .A2(MEM_stage_inst_dmem_n20290), .ZN(MEM_stage_inst_dmem_n9310) );
NAND2_X1 MEM_stage_inst_dmem_U19806 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n20297), .ZN(MEM_stage_inst_dmem_n20290) );
NAND2_X1 MEM_stage_inst_dmem_U19805 ( .A1(MEM_stage_inst_dmem_ram_3107), .A2(MEM_stage_inst_dmem_n20296), .ZN(MEM_stage_inst_dmem_n20291) );
NAND2_X1 MEM_stage_inst_dmem_U19804 ( .A1(MEM_stage_inst_dmem_n20289), .A2(MEM_stage_inst_dmem_n20288), .ZN(MEM_stage_inst_dmem_n9311) );
NAND2_X1 MEM_stage_inst_dmem_U19803 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n20297), .ZN(MEM_stage_inst_dmem_n20288) );
NAND2_X1 MEM_stage_inst_dmem_U19802 ( .A1(MEM_stage_inst_dmem_ram_3108), .A2(MEM_stage_inst_dmem_n20296), .ZN(MEM_stage_inst_dmem_n20289) );
NAND2_X1 MEM_stage_inst_dmem_U19801 ( .A1(MEM_stage_inst_dmem_n20287), .A2(MEM_stage_inst_dmem_n20286), .ZN(MEM_stage_inst_dmem_n9312) );
NAND2_X1 MEM_stage_inst_dmem_U19800 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n20297), .ZN(MEM_stage_inst_dmem_n20286) );
NAND2_X1 MEM_stage_inst_dmem_U19799 ( .A1(MEM_stage_inst_dmem_ram_3109), .A2(MEM_stage_inst_dmem_n20296), .ZN(MEM_stage_inst_dmem_n20287) );
NAND2_X1 MEM_stage_inst_dmem_U19798 ( .A1(MEM_stage_inst_dmem_n20285), .A2(MEM_stage_inst_dmem_n20284), .ZN(MEM_stage_inst_dmem_n9313) );
NAND2_X1 MEM_stage_inst_dmem_U19797 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n20297), .ZN(MEM_stage_inst_dmem_n20284) );
NAND2_X1 MEM_stage_inst_dmem_U19796 ( .A1(MEM_stage_inst_dmem_ram_3110), .A2(MEM_stage_inst_dmem_n20296), .ZN(MEM_stage_inst_dmem_n20285) );
NAND2_X1 MEM_stage_inst_dmem_U19795 ( .A1(MEM_stage_inst_dmem_n20283), .A2(MEM_stage_inst_dmem_n20282), .ZN(MEM_stage_inst_dmem_n9314) );
NAND2_X1 MEM_stage_inst_dmem_U19794 ( .A1(MEM_stage_inst_dmem_n112), .A2(MEM_stage_inst_dmem_n20297), .ZN(MEM_stage_inst_dmem_n20282) );
NAND2_X1 MEM_stage_inst_dmem_U19793 ( .A1(MEM_stage_inst_dmem_ram_3111), .A2(MEM_stage_inst_dmem_n20296), .ZN(MEM_stage_inst_dmem_n20283) );
NAND2_X1 MEM_stage_inst_dmem_U19792 ( .A1(MEM_stage_inst_dmem_n20281), .A2(MEM_stage_inst_dmem_n20280), .ZN(MEM_stage_inst_dmem_n9315) );
NAND2_X1 MEM_stage_inst_dmem_U19791 ( .A1(MEM_stage_inst_dmem_n111), .A2(MEM_stage_inst_dmem_n20297), .ZN(MEM_stage_inst_dmem_n20280) );
NAND2_X1 MEM_stage_inst_dmem_U19790 ( .A1(MEM_stage_inst_dmem_ram_3112), .A2(MEM_stage_inst_dmem_n20296), .ZN(MEM_stage_inst_dmem_n20281) );
NAND2_X1 MEM_stage_inst_dmem_U19789 ( .A1(MEM_stage_inst_dmem_n20279), .A2(MEM_stage_inst_dmem_n20278), .ZN(MEM_stage_inst_dmem_n9316) );
NAND2_X1 MEM_stage_inst_dmem_U19788 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n20297), .ZN(MEM_stage_inst_dmem_n20278) );
NAND2_X1 MEM_stage_inst_dmem_U19787 ( .A1(MEM_stage_inst_dmem_ram_3113), .A2(MEM_stage_inst_dmem_n20296), .ZN(MEM_stage_inst_dmem_n20279) );
NAND2_X1 MEM_stage_inst_dmem_U19786 ( .A1(MEM_stage_inst_dmem_n20277), .A2(MEM_stage_inst_dmem_n20276), .ZN(MEM_stage_inst_dmem_n9317) );
NAND2_X1 MEM_stage_inst_dmem_U19785 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n20297), .ZN(MEM_stage_inst_dmem_n20276) );
NAND2_X1 MEM_stage_inst_dmem_U19784 ( .A1(MEM_stage_inst_dmem_ram_3114), .A2(MEM_stage_inst_dmem_n20296), .ZN(MEM_stage_inst_dmem_n20277) );
NAND2_X1 MEM_stage_inst_dmem_U19783 ( .A1(MEM_stage_inst_dmem_n20275), .A2(MEM_stage_inst_dmem_n20274), .ZN(MEM_stage_inst_dmem_n9318) );
NAND2_X1 MEM_stage_inst_dmem_U19782 ( .A1(MEM_stage_inst_dmem_n18864), .A2(MEM_stage_inst_dmem_n20297), .ZN(MEM_stage_inst_dmem_n20274) );
NAND2_X1 MEM_stage_inst_dmem_U19781 ( .A1(MEM_stage_inst_dmem_ram_3115), .A2(MEM_stage_inst_dmem_n20296), .ZN(MEM_stage_inst_dmem_n20275) );
NAND2_X1 MEM_stage_inst_dmem_U19780 ( .A1(MEM_stage_inst_dmem_n20273), .A2(MEM_stage_inst_dmem_n20272), .ZN(MEM_stage_inst_dmem_n9319) );
NAND2_X1 MEM_stage_inst_dmem_U19779 ( .A1(MEM_stage_inst_dmem_n18861), .A2(MEM_stage_inst_dmem_n20297), .ZN(MEM_stage_inst_dmem_n20272) );
NAND2_X1 MEM_stage_inst_dmem_U19778 ( .A1(MEM_stage_inst_dmem_ram_3116), .A2(MEM_stage_inst_dmem_n20296), .ZN(MEM_stage_inst_dmem_n20273) );
NAND2_X1 MEM_stage_inst_dmem_U19777 ( .A1(MEM_stage_inst_dmem_n20271), .A2(MEM_stage_inst_dmem_n20270), .ZN(MEM_stage_inst_dmem_n9320) );
NAND2_X1 MEM_stage_inst_dmem_U19776 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n20297), .ZN(MEM_stage_inst_dmem_n20270) );
NAND2_X1 MEM_stage_inst_dmem_U19775 ( .A1(MEM_stage_inst_dmem_ram_3117), .A2(MEM_stage_inst_dmem_n20296), .ZN(MEM_stage_inst_dmem_n20271) );
NAND2_X1 MEM_stage_inst_dmem_U19774 ( .A1(MEM_stage_inst_dmem_n20269), .A2(MEM_stage_inst_dmem_n20268), .ZN(MEM_stage_inst_dmem_n9321) );
NAND2_X1 MEM_stage_inst_dmem_U19773 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n20297), .ZN(MEM_stage_inst_dmem_n20268) );
NAND2_X1 MEM_stage_inst_dmem_U19772 ( .A1(MEM_stage_inst_dmem_ram_3118), .A2(MEM_stage_inst_dmem_n20296), .ZN(MEM_stage_inst_dmem_n20269) );
NAND2_X1 MEM_stage_inst_dmem_U19771 ( .A1(MEM_stage_inst_dmem_n20267), .A2(MEM_stage_inst_dmem_n20266), .ZN(MEM_stage_inst_dmem_n9322) );
NAND2_X1 MEM_stage_inst_dmem_U19770 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n20297), .ZN(MEM_stage_inst_dmem_n20266) );
INV_X1 MEM_stage_inst_dmem_U19769 ( .A(MEM_stage_inst_dmem_n20296), .ZN(MEM_stage_inst_dmem_n20297) );
NAND2_X1 MEM_stage_inst_dmem_U19768 ( .A1(MEM_stage_inst_dmem_ram_3119), .A2(MEM_stage_inst_dmem_n20296), .ZN(MEM_stage_inst_dmem_n20267) );
NAND2_X1 MEM_stage_inst_dmem_U19767 ( .A1(MEM_stage_inst_dmem_n21394), .A2(MEM_stage_inst_dmem_n20334), .ZN(MEM_stage_inst_dmem_n20296) );
NAND2_X1 MEM_stage_inst_dmem_U19766 ( .A1(MEM_stage_inst_dmem_n20265), .A2(MEM_stage_inst_dmem_n20264), .ZN(MEM_stage_inst_dmem_n9323) );
NAND2_X1 MEM_stage_inst_dmem_U19765 ( .A1(MEM_stage_inst_dmem_n20551), .A2(MEM_stage_inst_dmem_n20263), .ZN(MEM_stage_inst_dmem_n20264) );
NAND2_X1 MEM_stage_inst_dmem_U19764 ( .A1(MEM_stage_inst_dmem_ram_3120), .A2(MEM_stage_inst_dmem_n20262), .ZN(MEM_stage_inst_dmem_n20265) );
NAND2_X1 MEM_stage_inst_dmem_U19763 ( .A1(MEM_stage_inst_dmem_n20261), .A2(MEM_stage_inst_dmem_n20260), .ZN(MEM_stage_inst_dmem_n9324) );
NAND2_X1 MEM_stage_inst_dmem_U19762 ( .A1(MEM_stage_inst_dmem_n20547), .A2(MEM_stage_inst_dmem_n20263), .ZN(MEM_stage_inst_dmem_n20260) );
NAND2_X1 MEM_stage_inst_dmem_U19761 ( .A1(MEM_stage_inst_dmem_ram_3121), .A2(MEM_stage_inst_dmem_n20262), .ZN(MEM_stage_inst_dmem_n20261) );
NAND2_X1 MEM_stage_inst_dmem_U19760 ( .A1(MEM_stage_inst_dmem_n20259), .A2(MEM_stage_inst_dmem_n20258), .ZN(MEM_stage_inst_dmem_n9325) );
NAND2_X1 MEM_stage_inst_dmem_U19759 ( .A1(MEM_stage_inst_dmem_n20544), .A2(MEM_stage_inst_dmem_n20263), .ZN(MEM_stage_inst_dmem_n20258) );
NAND2_X1 MEM_stage_inst_dmem_U19758 ( .A1(MEM_stage_inst_dmem_ram_3122), .A2(MEM_stage_inst_dmem_n20262), .ZN(MEM_stage_inst_dmem_n20259) );
NAND2_X1 MEM_stage_inst_dmem_U19757 ( .A1(MEM_stage_inst_dmem_n20257), .A2(MEM_stage_inst_dmem_n20256), .ZN(MEM_stage_inst_dmem_n9326) );
NAND2_X1 MEM_stage_inst_dmem_U19756 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n20263), .ZN(MEM_stage_inst_dmem_n20256) );
NAND2_X1 MEM_stage_inst_dmem_U19755 ( .A1(MEM_stage_inst_dmem_ram_3123), .A2(MEM_stage_inst_dmem_n20262), .ZN(MEM_stage_inst_dmem_n20257) );
NAND2_X1 MEM_stage_inst_dmem_U19754 ( .A1(MEM_stage_inst_dmem_n20255), .A2(MEM_stage_inst_dmem_n20254), .ZN(MEM_stage_inst_dmem_n9327) );
NAND2_X1 MEM_stage_inst_dmem_U19753 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n20263), .ZN(MEM_stage_inst_dmem_n20254) );
NAND2_X1 MEM_stage_inst_dmem_U19752 ( .A1(MEM_stage_inst_dmem_ram_3124), .A2(MEM_stage_inst_dmem_n20262), .ZN(MEM_stage_inst_dmem_n20255) );
NAND2_X1 MEM_stage_inst_dmem_U19751 ( .A1(MEM_stage_inst_dmem_n20253), .A2(MEM_stage_inst_dmem_n20252), .ZN(MEM_stage_inst_dmem_n9328) );
NAND2_X1 MEM_stage_inst_dmem_U19750 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n20263), .ZN(MEM_stage_inst_dmem_n20252) );
NAND2_X1 MEM_stage_inst_dmem_U19749 ( .A1(MEM_stage_inst_dmem_ram_3125), .A2(MEM_stage_inst_dmem_n20262), .ZN(MEM_stage_inst_dmem_n20253) );
NAND2_X1 MEM_stage_inst_dmem_U19748 ( .A1(MEM_stage_inst_dmem_n20251), .A2(MEM_stage_inst_dmem_n20250), .ZN(MEM_stage_inst_dmem_n9329) );
NAND2_X1 MEM_stage_inst_dmem_U19747 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n20263), .ZN(MEM_stage_inst_dmem_n20250) );
NAND2_X1 MEM_stage_inst_dmem_U19746 ( .A1(MEM_stage_inst_dmem_ram_3126), .A2(MEM_stage_inst_dmem_n20262), .ZN(MEM_stage_inst_dmem_n20251) );
NAND2_X1 MEM_stage_inst_dmem_U19745 ( .A1(MEM_stage_inst_dmem_n20249), .A2(MEM_stage_inst_dmem_n20248), .ZN(MEM_stage_inst_dmem_n9330) );
NAND2_X1 MEM_stage_inst_dmem_U19744 ( .A1(MEM_stage_inst_dmem_n20530), .A2(MEM_stage_inst_dmem_n20263), .ZN(MEM_stage_inst_dmem_n20248) );
NAND2_X1 MEM_stage_inst_dmem_U19743 ( .A1(MEM_stage_inst_dmem_ram_3127), .A2(MEM_stage_inst_dmem_n20262), .ZN(MEM_stage_inst_dmem_n20249) );
NAND2_X1 MEM_stage_inst_dmem_U19742 ( .A1(MEM_stage_inst_dmem_n20247), .A2(MEM_stage_inst_dmem_n20246), .ZN(MEM_stage_inst_dmem_n9331) );
NAND2_X1 MEM_stage_inst_dmem_U19741 ( .A1(MEM_stage_inst_dmem_n20527), .A2(MEM_stage_inst_dmem_n20263), .ZN(MEM_stage_inst_dmem_n20246) );
NAND2_X1 MEM_stage_inst_dmem_U19740 ( .A1(MEM_stage_inst_dmem_ram_3128), .A2(MEM_stage_inst_dmem_n20262), .ZN(MEM_stage_inst_dmem_n20247) );
NAND2_X1 MEM_stage_inst_dmem_U19739 ( .A1(MEM_stage_inst_dmem_n20245), .A2(MEM_stage_inst_dmem_n20244), .ZN(MEM_stage_inst_dmem_n9332) );
NAND2_X1 MEM_stage_inst_dmem_U19738 ( .A1(MEM_stage_inst_dmem_n20524), .A2(MEM_stage_inst_dmem_n20263), .ZN(MEM_stage_inst_dmem_n20244) );
NAND2_X1 MEM_stage_inst_dmem_U19737 ( .A1(MEM_stage_inst_dmem_ram_3129), .A2(MEM_stage_inst_dmem_n20262), .ZN(MEM_stage_inst_dmem_n20245) );
NAND2_X1 MEM_stage_inst_dmem_U19736 ( .A1(MEM_stage_inst_dmem_n20243), .A2(MEM_stage_inst_dmem_n20242), .ZN(MEM_stage_inst_dmem_n9333) );
NAND2_X1 MEM_stage_inst_dmem_U19735 ( .A1(MEM_stage_inst_dmem_n20521), .A2(MEM_stage_inst_dmem_n20263), .ZN(MEM_stage_inst_dmem_n20242) );
NAND2_X1 MEM_stage_inst_dmem_U19734 ( .A1(MEM_stage_inst_dmem_ram_3130), .A2(MEM_stage_inst_dmem_n20262), .ZN(MEM_stage_inst_dmem_n20243) );
NAND2_X1 MEM_stage_inst_dmem_U19733 ( .A1(MEM_stage_inst_dmem_n20241), .A2(MEM_stage_inst_dmem_n20240), .ZN(MEM_stage_inst_dmem_n9334) );
NAND2_X1 MEM_stage_inst_dmem_U19732 ( .A1(MEM_stage_inst_dmem_n20518), .A2(MEM_stage_inst_dmem_n20263), .ZN(MEM_stage_inst_dmem_n20240) );
NAND2_X1 MEM_stage_inst_dmem_U19731 ( .A1(MEM_stage_inst_dmem_ram_3131), .A2(MEM_stage_inst_dmem_n20262), .ZN(MEM_stage_inst_dmem_n20241) );
NAND2_X1 MEM_stage_inst_dmem_U19730 ( .A1(MEM_stage_inst_dmem_n20239), .A2(MEM_stage_inst_dmem_n20238), .ZN(MEM_stage_inst_dmem_n9335) );
NAND2_X1 MEM_stage_inst_dmem_U19729 ( .A1(MEM_stage_inst_dmem_n20515), .A2(MEM_stage_inst_dmem_n20263), .ZN(MEM_stage_inst_dmem_n20238) );
NAND2_X1 MEM_stage_inst_dmem_U19728 ( .A1(MEM_stage_inst_dmem_ram_3132), .A2(MEM_stage_inst_dmem_n20262), .ZN(MEM_stage_inst_dmem_n20239) );
NAND2_X1 MEM_stage_inst_dmem_U19727 ( .A1(MEM_stage_inst_dmem_n20237), .A2(MEM_stage_inst_dmem_n20236), .ZN(MEM_stage_inst_dmem_n9336) );
NAND2_X1 MEM_stage_inst_dmem_U19726 ( .A1(MEM_stage_inst_dmem_n20512), .A2(MEM_stage_inst_dmem_n20263), .ZN(MEM_stage_inst_dmem_n20236) );
NAND2_X1 MEM_stage_inst_dmem_U19725 ( .A1(MEM_stage_inst_dmem_ram_3133), .A2(MEM_stage_inst_dmem_n20262), .ZN(MEM_stage_inst_dmem_n20237) );
NAND2_X1 MEM_stage_inst_dmem_U19724 ( .A1(MEM_stage_inst_dmem_n20235), .A2(MEM_stage_inst_dmem_n20234), .ZN(MEM_stage_inst_dmem_n9337) );
NAND2_X1 MEM_stage_inst_dmem_U19723 ( .A1(MEM_stage_inst_dmem_n20509), .A2(MEM_stage_inst_dmem_n20263), .ZN(MEM_stage_inst_dmem_n20234) );
NAND2_X1 MEM_stage_inst_dmem_U19722 ( .A1(MEM_stage_inst_dmem_ram_3134), .A2(MEM_stage_inst_dmem_n20262), .ZN(MEM_stage_inst_dmem_n20235) );
NAND2_X1 MEM_stage_inst_dmem_U19721 ( .A1(MEM_stage_inst_dmem_n20233), .A2(MEM_stage_inst_dmem_n20232), .ZN(MEM_stage_inst_dmem_n9338) );
NAND2_X1 MEM_stage_inst_dmem_U19720 ( .A1(MEM_stage_inst_dmem_n20506), .A2(MEM_stage_inst_dmem_n20263), .ZN(MEM_stage_inst_dmem_n20232) );
INV_X1 MEM_stage_inst_dmem_U19719 ( .A(MEM_stage_inst_dmem_n20262), .ZN(MEM_stage_inst_dmem_n20263) );
NAND2_X1 MEM_stage_inst_dmem_U19718 ( .A1(MEM_stage_inst_dmem_ram_3135), .A2(MEM_stage_inst_dmem_n20262), .ZN(MEM_stage_inst_dmem_n20233) );
NAND2_X1 MEM_stage_inst_dmem_U19717 ( .A1(MEM_stage_inst_dmem_n21359), .A2(MEM_stage_inst_dmem_n20334), .ZN(MEM_stage_inst_dmem_n20262) );
NAND2_X1 MEM_stage_inst_dmem_U19716 ( .A1(MEM_stage_inst_dmem_n20231), .A2(MEM_stage_inst_dmem_n20230), .ZN(MEM_stage_inst_dmem_n9339) );
NAND2_X1 MEM_stage_inst_dmem_U19715 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n20229), .ZN(MEM_stage_inst_dmem_n20230) );
NAND2_X1 MEM_stage_inst_dmem_U19714 ( .A1(MEM_stage_inst_dmem_ram_3136), .A2(MEM_stage_inst_dmem_n20228), .ZN(MEM_stage_inst_dmem_n20231) );
NAND2_X1 MEM_stage_inst_dmem_U19713 ( .A1(MEM_stage_inst_dmem_n20227), .A2(MEM_stage_inst_dmem_n20226), .ZN(MEM_stage_inst_dmem_n9340) );
NAND2_X1 MEM_stage_inst_dmem_U19712 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n20229), .ZN(MEM_stage_inst_dmem_n20226) );
NAND2_X1 MEM_stage_inst_dmem_U19711 ( .A1(MEM_stage_inst_dmem_ram_3137), .A2(MEM_stage_inst_dmem_n20228), .ZN(MEM_stage_inst_dmem_n20227) );
NAND2_X1 MEM_stage_inst_dmem_U19710 ( .A1(MEM_stage_inst_dmem_n20225), .A2(MEM_stage_inst_dmem_n20224), .ZN(MEM_stage_inst_dmem_n9341) );
NAND2_X1 MEM_stage_inst_dmem_U19709 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n20229), .ZN(MEM_stage_inst_dmem_n20224) );
NAND2_X1 MEM_stage_inst_dmem_U19708 ( .A1(MEM_stage_inst_dmem_ram_3138), .A2(MEM_stage_inst_dmem_n20228), .ZN(MEM_stage_inst_dmem_n20225) );
NAND2_X1 MEM_stage_inst_dmem_U19707 ( .A1(MEM_stage_inst_dmem_n20223), .A2(MEM_stage_inst_dmem_n20222), .ZN(MEM_stage_inst_dmem_n9342) );
NAND2_X1 MEM_stage_inst_dmem_U19706 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n20229), .ZN(MEM_stage_inst_dmem_n20222) );
NAND2_X1 MEM_stage_inst_dmem_U19705 ( .A1(MEM_stage_inst_dmem_ram_3139), .A2(MEM_stage_inst_dmem_n20228), .ZN(MEM_stage_inst_dmem_n20223) );
NAND2_X1 MEM_stage_inst_dmem_U19704 ( .A1(MEM_stage_inst_dmem_n20221), .A2(MEM_stage_inst_dmem_n20220), .ZN(MEM_stage_inst_dmem_n9343) );
NAND2_X1 MEM_stage_inst_dmem_U19703 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n20229), .ZN(MEM_stage_inst_dmem_n20220) );
NAND2_X1 MEM_stage_inst_dmem_U19702 ( .A1(MEM_stage_inst_dmem_ram_3140), .A2(MEM_stage_inst_dmem_n20228), .ZN(MEM_stage_inst_dmem_n20221) );
NAND2_X1 MEM_stage_inst_dmem_U19701 ( .A1(MEM_stage_inst_dmem_n20219), .A2(MEM_stage_inst_dmem_n20218), .ZN(MEM_stage_inst_dmem_n9344) );
NAND2_X1 MEM_stage_inst_dmem_U19700 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n20229), .ZN(MEM_stage_inst_dmem_n20218) );
NAND2_X1 MEM_stage_inst_dmem_U19699 ( .A1(MEM_stage_inst_dmem_ram_3141), .A2(MEM_stage_inst_dmem_n20228), .ZN(MEM_stage_inst_dmem_n20219) );
NAND2_X1 MEM_stage_inst_dmem_U19698 ( .A1(MEM_stage_inst_dmem_n20217), .A2(MEM_stage_inst_dmem_n20216), .ZN(MEM_stage_inst_dmem_n9345) );
NAND2_X1 MEM_stage_inst_dmem_U19697 ( .A1(MEM_stage_inst_dmem_n21340), .A2(MEM_stage_inst_dmem_n20229), .ZN(MEM_stage_inst_dmem_n20216) );
NAND2_X1 MEM_stage_inst_dmem_U19696 ( .A1(MEM_stage_inst_dmem_ram_3142), .A2(MEM_stage_inst_dmem_n20228), .ZN(MEM_stage_inst_dmem_n20217) );
NAND2_X1 MEM_stage_inst_dmem_U19695 ( .A1(MEM_stage_inst_dmem_n20215), .A2(MEM_stage_inst_dmem_n20214), .ZN(MEM_stage_inst_dmem_n9346) );
NAND2_X1 MEM_stage_inst_dmem_U19694 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n20229), .ZN(MEM_stage_inst_dmem_n20214) );
NAND2_X1 MEM_stage_inst_dmem_U19693 ( .A1(MEM_stage_inst_dmem_ram_3143), .A2(MEM_stage_inst_dmem_n20228), .ZN(MEM_stage_inst_dmem_n20215) );
NAND2_X1 MEM_stage_inst_dmem_U19692 ( .A1(MEM_stage_inst_dmem_n20213), .A2(MEM_stage_inst_dmem_n20212), .ZN(MEM_stage_inst_dmem_n9347) );
NAND2_X1 MEM_stage_inst_dmem_U19691 ( .A1(MEM_stage_inst_dmem_n13051), .A2(MEM_stage_inst_dmem_n20229), .ZN(MEM_stage_inst_dmem_n20212) );
NAND2_X1 MEM_stage_inst_dmem_U19690 ( .A1(MEM_stage_inst_dmem_ram_3144), .A2(MEM_stage_inst_dmem_n20228), .ZN(MEM_stage_inst_dmem_n20213) );
NAND2_X1 MEM_stage_inst_dmem_U19689 ( .A1(MEM_stage_inst_dmem_n20211), .A2(MEM_stage_inst_dmem_n20210), .ZN(MEM_stage_inst_dmem_n9348) );
NAND2_X1 MEM_stage_inst_dmem_U19688 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n20229), .ZN(MEM_stage_inst_dmem_n20210) );
NAND2_X1 MEM_stage_inst_dmem_U19687 ( .A1(MEM_stage_inst_dmem_ram_3145), .A2(MEM_stage_inst_dmem_n20228), .ZN(MEM_stage_inst_dmem_n20211) );
NAND2_X1 MEM_stage_inst_dmem_U19686 ( .A1(MEM_stage_inst_dmem_n20209), .A2(MEM_stage_inst_dmem_n20208), .ZN(MEM_stage_inst_dmem_n9349) );
NAND2_X1 MEM_stage_inst_dmem_U19685 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n20229), .ZN(MEM_stage_inst_dmem_n20208) );
NAND2_X1 MEM_stage_inst_dmem_U19684 ( .A1(MEM_stage_inst_dmem_ram_3146), .A2(MEM_stage_inst_dmem_n20228), .ZN(MEM_stage_inst_dmem_n20209) );
NAND2_X1 MEM_stage_inst_dmem_U19683 ( .A1(MEM_stage_inst_dmem_n20207), .A2(MEM_stage_inst_dmem_n20206), .ZN(MEM_stage_inst_dmem_n9350) );
NAND2_X1 MEM_stage_inst_dmem_U19682 ( .A1(EX_pipeline_reg_out_16), .A2(MEM_stage_inst_dmem_n20229), .ZN(MEM_stage_inst_dmem_n20206) );
NAND2_X1 MEM_stage_inst_dmem_U19681 ( .A1(MEM_stage_inst_dmem_ram_3147), .A2(MEM_stage_inst_dmem_n20228), .ZN(MEM_stage_inst_dmem_n20207) );
NAND2_X1 MEM_stage_inst_dmem_U19680 ( .A1(MEM_stage_inst_dmem_n20205), .A2(MEM_stage_inst_dmem_n20204), .ZN(MEM_stage_inst_dmem_n9351) );
NAND2_X1 MEM_stage_inst_dmem_U19679 ( .A1(EX_pipeline_reg_out_17), .A2(MEM_stage_inst_dmem_n20229), .ZN(MEM_stage_inst_dmem_n20204) );
NAND2_X1 MEM_stage_inst_dmem_U19678 ( .A1(MEM_stage_inst_dmem_ram_3148), .A2(MEM_stage_inst_dmem_n20228), .ZN(MEM_stage_inst_dmem_n20205) );
NAND2_X1 MEM_stage_inst_dmem_U19677 ( .A1(MEM_stage_inst_dmem_n20203), .A2(MEM_stage_inst_dmem_n20202), .ZN(MEM_stage_inst_dmem_n9352) );
NAND2_X1 MEM_stage_inst_dmem_U19676 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n20229), .ZN(MEM_stage_inst_dmem_n20202) );
NAND2_X1 MEM_stage_inst_dmem_U19675 ( .A1(MEM_stage_inst_dmem_ram_3149), .A2(MEM_stage_inst_dmem_n20228), .ZN(MEM_stage_inst_dmem_n20203) );
NAND2_X1 MEM_stage_inst_dmem_U19674 ( .A1(MEM_stage_inst_dmem_n20201), .A2(MEM_stage_inst_dmem_n20200), .ZN(MEM_stage_inst_dmem_n9353) );
NAND2_X1 MEM_stage_inst_dmem_U19673 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n20229), .ZN(MEM_stage_inst_dmem_n20200) );
NAND2_X1 MEM_stage_inst_dmem_U19672 ( .A1(MEM_stage_inst_dmem_ram_3150), .A2(MEM_stage_inst_dmem_n20228), .ZN(MEM_stage_inst_dmem_n20201) );
NAND2_X1 MEM_stage_inst_dmem_U19671 ( .A1(MEM_stage_inst_dmem_n20199), .A2(MEM_stage_inst_dmem_n20198), .ZN(MEM_stage_inst_dmem_n9354) );
NAND2_X1 MEM_stage_inst_dmem_U19670 ( .A1(MEM_stage_inst_dmem_n15110), .A2(MEM_stage_inst_dmem_n20229), .ZN(MEM_stage_inst_dmem_n20198) );
INV_X1 MEM_stage_inst_dmem_U19669 ( .A(MEM_stage_inst_dmem_n20228), .ZN(MEM_stage_inst_dmem_n20229) );
NAND2_X1 MEM_stage_inst_dmem_U19668 ( .A1(MEM_stage_inst_dmem_ram_3151), .A2(MEM_stage_inst_dmem_n20228), .ZN(MEM_stage_inst_dmem_n20199) );
NAND2_X1 MEM_stage_inst_dmem_U19667 ( .A1(MEM_stage_inst_dmem_n21319), .A2(MEM_stage_inst_dmem_n20334), .ZN(MEM_stage_inst_dmem_n20228) );
NAND2_X1 MEM_stage_inst_dmem_U19666 ( .A1(MEM_stage_inst_dmem_n20197), .A2(MEM_stage_inst_dmem_n20196), .ZN(MEM_stage_inst_dmem_n9355) );
NAND2_X1 MEM_stage_inst_dmem_U19665 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n20195), .ZN(MEM_stage_inst_dmem_n20196) );
NAND2_X1 MEM_stage_inst_dmem_U19664 ( .A1(MEM_stage_inst_dmem_ram_3152), .A2(MEM_stage_inst_dmem_n20194), .ZN(MEM_stage_inst_dmem_n20197) );
NAND2_X1 MEM_stage_inst_dmem_U19663 ( .A1(MEM_stage_inst_dmem_n20193), .A2(MEM_stage_inst_dmem_n20192), .ZN(MEM_stage_inst_dmem_n9356) );
NAND2_X1 MEM_stage_inst_dmem_U19662 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n20195), .ZN(MEM_stage_inst_dmem_n20192) );
NAND2_X1 MEM_stage_inst_dmem_U19661 ( .A1(MEM_stage_inst_dmem_ram_3153), .A2(MEM_stage_inst_dmem_n20194), .ZN(MEM_stage_inst_dmem_n20193) );
NAND2_X1 MEM_stage_inst_dmem_U19660 ( .A1(MEM_stage_inst_dmem_n20191), .A2(MEM_stage_inst_dmem_n20190), .ZN(MEM_stage_inst_dmem_n9357) );
NAND2_X1 MEM_stage_inst_dmem_U19659 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n20195), .ZN(MEM_stage_inst_dmem_n20190) );
NAND2_X1 MEM_stage_inst_dmem_U19658 ( .A1(MEM_stage_inst_dmem_ram_3154), .A2(MEM_stage_inst_dmem_n20194), .ZN(MEM_stage_inst_dmem_n20191) );
NAND2_X1 MEM_stage_inst_dmem_U19657 ( .A1(MEM_stage_inst_dmem_n20189), .A2(MEM_stage_inst_dmem_n20188), .ZN(MEM_stage_inst_dmem_n9358) );
NAND2_X1 MEM_stage_inst_dmem_U19656 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n20195), .ZN(MEM_stage_inst_dmem_n20188) );
NAND2_X1 MEM_stage_inst_dmem_U19655 ( .A1(MEM_stage_inst_dmem_ram_3155), .A2(MEM_stage_inst_dmem_n20194), .ZN(MEM_stage_inst_dmem_n20189) );
NAND2_X1 MEM_stage_inst_dmem_U19654 ( .A1(MEM_stage_inst_dmem_n20187), .A2(MEM_stage_inst_dmem_n20186), .ZN(MEM_stage_inst_dmem_n9359) );
NAND2_X1 MEM_stage_inst_dmem_U19653 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n20195), .ZN(MEM_stage_inst_dmem_n20186) );
NAND2_X1 MEM_stage_inst_dmem_U19652 ( .A1(MEM_stage_inst_dmem_ram_3156), .A2(MEM_stage_inst_dmem_n20194), .ZN(MEM_stage_inst_dmem_n20187) );
NAND2_X1 MEM_stage_inst_dmem_U19651 ( .A1(MEM_stage_inst_dmem_n20185), .A2(MEM_stage_inst_dmem_n20184), .ZN(MEM_stage_inst_dmem_n9360) );
NAND2_X1 MEM_stage_inst_dmem_U19650 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n20195), .ZN(MEM_stage_inst_dmem_n20184) );
NAND2_X1 MEM_stage_inst_dmem_U19649 ( .A1(MEM_stage_inst_dmem_ram_3157), .A2(MEM_stage_inst_dmem_n20194), .ZN(MEM_stage_inst_dmem_n20185) );
NAND2_X1 MEM_stage_inst_dmem_U19648 ( .A1(MEM_stage_inst_dmem_n20183), .A2(MEM_stage_inst_dmem_n20182), .ZN(MEM_stage_inst_dmem_n9361) );
NAND2_X1 MEM_stage_inst_dmem_U19647 ( .A1(MEM_stage_inst_dmem_n14717), .A2(MEM_stage_inst_dmem_n20195), .ZN(MEM_stage_inst_dmem_n20182) );
NAND2_X1 MEM_stage_inst_dmem_U19646 ( .A1(MEM_stage_inst_dmem_ram_3158), .A2(MEM_stage_inst_dmem_n20194), .ZN(MEM_stage_inst_dmem_n20183) );
NAND2_X1 MEM_stage_inst_dmem_U19645 ( .A1(MEM_stage_inst_dmem_n20181), .A2(MEM_stage_inst_dmem_n20180), .ZN(MEM_stage_inst_dmem_n9362) );
NAND2_X1 MEM_stage_inst_dmem_U19644 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n20195), .ZN(MEM_stage_inst_dmem_n20180) );
NAND2_X1 MEM_stage_inst_dmem_U19643 ( .A1(MEM_stage_inst_dmem_ram_3159), .A2(MEM_stage_inst_dmem_n20194), .ZN(MEM_stage_inst_dmem_n20181) );
NAND2_X1 MEM_stage_inst_dmem_U19642 ( .A1(MEM_stage_inst_dmem_n20179), .A2(MEM_stage_inst_dmem_n20178), .ZN(MEM_stage_inst_dmem_n9363) );
NAND2_X1 MEM_stage_inst_dmem_U19641 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n20195), .ZN(MEM_stage_inst_dmem_n20178) );
NAND2_X1 MEM_stage_inst_dmem_U19640 ( .A1(MEM_stage_inst_dmem_ram_3160), .A2(MEM_stage_inst_dmem_n20194), .ZN(MEM_stage_inst_dmem_n20179) );
NAND2_X1 MEM_stage_inst_dmem_U19639 ( .A1(MEM_stage_inst_dmem_n20177), .A2(MEM_stage_inst_dmem_n20176), .ZN(MEM_stage_inst_dmem_n9364) );
NAND2_X1 MEM_stage_inst_dmem_U19638 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n20195), .ZN(MEM_stage_inst_dmem_n20176) );
NAND2_X1 MEM_stage_inst_dmem_U19637 ( .A1(MEM_stage_inst_dmem_ram_3161), .A2(MEM_stage_inst_dmem_n20194), .ZN(MEM_stage_inst_dmem_n20177) );
NAND2_X1 MEM_stage_inst_dmem_U19636 ( .A1(MEM_stage_inst_dmem_n20175), .A2(MEM_stage_inst_dmem_n20174), .ZN(MEM_stage_inst_dmem_n9365) );
NAND2_X1 MEM_stage_inst_dmem_U19635 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n20195), .ZN(MEM_stage_inst_dmem_n20174) );
NAND2_X1 MEM_stage_inst_dmem_U19634 ( .A1(MEM_stage_inst_dmem_ram_3162), .A2(MEM_stage_inst_dmem_n20194), .ZN(MEM_stage_inst_dmem_n20175) );
NAND2_X1 MEM_stage_inst_dmem_U19633 ( .A1(MEM_stage_inst_dmem_n20173), .A2(MEM_stage_inst_dmem_n20172), .ZN(MEM_stage_inst_dmem_n9366) );
NAND2_X1 MEM_stage_inst_dmem_U19632 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n20195), .ZN(MEM_stage_inst_dmem_n20172) );
NAND2_X1 MEM_stage_inst_dmem_U19631 ( .A1(MEM_stage_inst_dmem_ram_3163), .A2(MEM_stage_inst_dmem_n20194), .ZN(MEM_stage_inst_dmem_n20173) );
NAND2_X1 MEM_stage_inst_dmem_U19630 ( .A1(MEM_stage_inst_dmem_n20171), .A2(MEM_stage_inst_dmem_n20170), .ZN(MEM_stage_inst_dmem_n9367) );
NAND2_X1 MEM_stage_inst_dmem_U19629 ( .A1(MEM_stage_inst_dmem_n21474), .A2(MEM_stage_inst_dmem_n20195), .ZN(MEM_stage_inst_dmem_n20170) );
NAND2_X1 MEM_stage_inst_dmem_U19628 ( .A1(MEM_stage_inst_dmem_ram_3164), .A2(MEM_stage_inst_dmem_n20194), .ZN(MEM_stage_inst_dmem_n20171) );
NAND2_X1 MEM_stage_inst_dmem_U19627 ( .A1(MEM_stage_inst_dmem_n20169), .A2(MEM_stage_inst_dmem_n20168), .ZN(MEM_stage_inst_dmem_n9368) );
NAND2_X1 MEM_stage_inst_dmem_U19626 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n20195), .ZN(MEM_stage_inst_dmem_n20168) );
NAND2_X1 MEM_stage_inst_dmem_U19625 ( .A1(MEM_stage_inst_dmem_ram_3165), .A2(MEM_stage_inst_dmem_n20194), .ZN(MEM_stage_inst_dmem_n20169) );
NAND2_X1 MEM_stage_inst_dmem_U19624 ( .A1(MEM_stage_inst_dmem_n20167), .A2(MEM_stage_inst_dmem_n20166), .ZN(MEM_stage_inst_dmem_n9369) );
NAND2_X1 MEM_stage_inst_dmem_U19623 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n20195), .ZN(MEM_stage_inst_dmem_n20166) );
NAND2_X1 MEM_stage_inst_dmem_U19622 ( .A1(MEM_stage_inst_dmem_ram_3166), .A2(MEM_stage_inst_dmem_n20194), .ZN(MEM_stage_inst_dmem_n20167) );
NAND2_X1 MEM_stage_inst_dmem_U19621 ( .A1(MEM_stage_inst_dmem_n20165), .A2(MEM_stage_inst_dmem_n20164), .ZN(MEM_stage_inst_dmem_n9370) );
NAND2_X1 MEM_stage_inst_dmem_U19620 ( .A1(MEM_stage_inst_dmem_n16758), .A2(MEM_stage_inst_dmem_n20195), .ZN(MEM_stage_inst_dmem_n20164) );
INV_X1 MEM_stage_inst_dmem_U19619 ( .A(MEM_stage_inst_dmem_n20194), .ZN(MEM_stage_inst_dmem_n20195) );
NAND2_X1 MEM_stage_inst_dmem_U19618 ( .A1(MEM_stage_inst_dmem_ram_3167), .A2(MEM_stage_inst_dmem_n20194), .ZN(MEM_stage_inst_dmem_n20165) );
NAND2_X1 MEM_stage_inst_dmem_U19617 ( .A1(MEM_stage_inst_dmem_n21284), .A2(MEM_stage_inst_dmem_n20334), .ZN(MEM_stage_inst_dmem_n20194) );
NAND2_X1 MEM_stage_inst_dmem_U19616 ( .A1(MEM_stage_inst_dmem_n20163), .A2(MEM_stage_inst_dmem_n20162), .ZN(MEM_stage_inst_dmem_n9371) );
NAND2_X1 MEM_stage_inst_dmem_U19615 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n20161), .ZN(MEM_stage_inst_dmem_n20162) );
NAND2_X1 MEM_stage_inst_dmem_U19614 ( .A1(MEM_stage_inst_dmem_ram_3168), .A2(MEM_stage_inst_dmem_n20160), .ZN(MEM_stage_inst_dmem_n20163) );
NAND2_X1 MEM_stage_inst_dmem_U19613 ( .A1(MEM_stage_inst_dmem_n20159), .A2(MEM_stage_inst_dmem_n20158), .ZN(MEM_stage_inst_dmem_n9372) );
NAND2_X1 MEM_stage_inst_dmem_U19612 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n20161), .ZN(MEM_stage_inst_dmem_n20158) );
NAND2_X1 MEM_stage_inst_dmem_U19611 ( .A1(MEM_stage_inst_dmem_ram_3169), .A2(MEM_stage_inst_dmem_n20160), .ZN(MEM_stage_inst_dmem_n20159) );
NAND2_X1 MEM_stage_inst_dmem_U19610 ( .A1(MEM_stage_inst_dmem_n20157), .A2(MEM_stage_inst_dmem_n20156), .ZN(MEM_stage_inst_dmem_n9373) );
NAND2_X1 MEM_stage_inst_dmem_U19609 ( .A1(MEM_stage_inst_dmem_n18887), .A2(MEM_stage_inst_dmem_n20161), .ZN(MEM_stage_inst_dmem_n20156) );
NAND2_X1 MEM_stage_inst_dmem_U19608 ( .A1(MEM_stage_inst_dmem_ram_3170), .A2(MEM_stage_inst_dmem_n20160), .ZN(MEM_stage_inst_dmem_n20157) );
NAND2_X1 MEM_stage_inst_dmem_U19607 ( .A1(MEM_stage_inst_dmem_n20155), .A2(MEM_stage_inst_dmem_n20154), .ZN(MEM_stage_inst_dmem_n9374) );
NAND2_X1 MEM_stage_inst_dmem_U19606 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n20161), .ZN(MEM_stage_inst_dmem_n20154) );
NAND2_X1 MEM_stage_inst_dmem_U19605 ( .A1(MEM_stage_inst_dmem_ram_3171), .A2(MEM_stage_inst_dmem_n20160), .ZN(MEM_stage_inst_dmem_n20155) );
NAND2_X1 MEM_stage_inst_dmem_U19604 ( .A1(MEM_stage_inst_dmem_n20153), .A2(MEM_stage_inst_dmem_n20152), .ZN(MEM_stage_inst_dmem_n9375) );
NAND2_X1 MEM_stage_inst_dmem_U19603 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n20161), .ZN(MEM_stage_inst_dmem_n20152) );
NAND2_X1 MEM_stage_inst_dmem_U19602 ( .A1(MEM_stage_inst_dmem_ram_3172), .A2(MEM_stage_inst_dmem_n20160), .ZN(MEM_stage_inst_dmem_n20153) );
NAND2_X1 MEM_stage_inst_dmem_U19601 ( .A1(MEM_stage_inst_dmem_n20151), .A2(MEM_stage_inst_dmem_n20150), .ZN(MEM_stage_inst_dmem_n9376) );
NAND2_X1 MEM_stage_inst_dmem_U19600 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n20161), .ZN(MEM_stage_inst_dmem_n20150) );
NAND2_X1 MEM_stage_inst_dmem_U19599 ( .A1(MEM_stage_inst_dmem_ram_3173), .A2(MEM_stage_inst_dmem_n20160), .ZN(MEM_stage_inst_dmem_n20151) );
NAND2_X1 MEM_stage_inst_dmem_U19598 ( .A1(MEM_stage_inst_dmem_n20149), .A2(MEM_stage_inst_dmem_n20148), .ZN(MEM_stage_inst_dmem_n9377) );
NAND2_X1 MEM_stage_inst_dmem_U19597 ( .A1(EX_pipeline_reg_out_11), .A2(MEM_stage_inst_dmem_n20161), .ZN(MEM_stage_inst_dmem_n20148) );
NAND2_X1 MEM_stage_inst_dmem_U19596 ( .A1(MEM_stage_inst_dmem_ram_3174), .A2(MEM_stage_inst_dmem_n20160), .ZN(MEM_stage_inst_dmem_n20149) );
NAND2_X1 MEM_stage_inst_dmem_U19595 ( .A1(MEM_stage_inst_dmem_n20147), .A2(MEM_stage_inst_dmem_n20146), .ZN(MEM_stage_inst_dmem_n9378) );
NAND2_X1 MEM_stage_inst_dmem_U19594 ( .A1(MEM_stage_inst_dmem_n112), .A2(MEM_stage_inst_dmem_n20161), .ZN(MEM_stage_inst_dmem_n20146) );
NAND2_X1 MEM_stage_inst_dmem_U19593 ( .A1(MEM_stage_inst_dmem_ram_3175), .A2(MEM_stage_inst_dmem_n20160), .ZN(MEM_stage_inst_dmem_n20147) );
NAND2_X1 MEM_stage_inst_dmem_U19592 ( .A1(MEM_stage_inst_dmem_n20145), .A2(MEM_stage_inst_dmem_n20144), .ZN(MEM_stage_inst_dmem_n9379) );
NAND2_X1 MEM_stage_inst_dmem_U19591 ( .A1(MEM_stage_inst_dmem_n20527), .A2(MEM_stage_inst_dmem_n20161), .ZN(MEM_stage_inst_dmem_n20144) );
NAND2_X1 MEM_stage_inst_dmem_U19590 ( .A1(MEM_stage_inst_dmem_ram_3176), .A2(MEM_stage_inst_dmem_n20160), .ZN(MEM_stage_inst_dmem_n20145) );
NAND2_X1 MEM_stage_inst_dmem_U19589 ( .A1(MEM_stage_inst_dmem_n20143), .A2(MEM_stage_inst_dmem_n20142), .ZN(MEM_stage_inst_dmem_n9380) );
NAND2_X1 MEM_stage_inst_dmem_U19588 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n20161), .ZN(MEM_stage_inst_dmem_n20142) );
NAND2_X1 MEM_stage_inst_dmem_U19587 ( .A1(MEM_stage_inst_dmem_ram_3177), .A2(MEM_stage_inst_dmem_n20160), .ZN(MEM_stage_inst_dmem_n20143) );
NAND2_X1 MEM_stage_inst_dmem_U19586 ( .A1(MEM_stage_inst_dmem_n20141), .A2(MEM_stage_inst_dmem_n20140), .ZN(MEM_stage_inst_dmem_n9381) );
NAND2_X1 MEM_stage_inst_dmem_U19585 ( .A1(MEM_stage_inst_dmem_n18867), .A2(MEM_stage_inst_dmem_n20161), .ZN(MEM_stage_inst_dmem_n20140) );
NAND2_X1 MEM_stage_inst_dmem_U19584 ( .A1(MEM_stage_inst_dmem_ram_3178), .A2(MEM_stage_inst_dmem_n20160), .ZN(MEM_stage_inst_dmem_n20141) );
NAND2_X1 MEM_stage_inst_dmem_U19583 ( .A1(MEM_stage_inst_dmem_n20139), .A2(MEM_stage_inst_dmem_n20138), .ZN(MEM_stage_inst_dmem_n9382) );
NAND2_X1 MEM_stage_inst_dmem_U19582 ( .A1(MEM_stage_inst_dmem_n20518), .A2(MEM_stage_inst_dmem_n20161), .ZN(MEM_stage_inst_dmem_n20138) );
NAND2_X1 MEM_stage_inst_dmem_U19581 ( .A1(MEM_stage_inst_dmem_ram_3179), .A2(MEM_stage_inst_dmem_n20160), .ZN(MEM_stage_inst_dmem_n20139) );
NAND2_X1 MEM_stage_inst_dmem_U19580 ( .A1(MEM_stage_inst_dmem_n20137), .A2(MEM_stage_inst_dmem_n20136), .ZN(MEM_stage_inst_dmem_n9383) );
NAND2_X1 MEM_stage_inst_dmem_U19579 ( .A1(MEM_stage_inst_dmem_n20515), .A2(MEM_stage_inst_dmem_n20161), .ZN(MEM_stage_inst_dmem_n20136) );
NAND2_X1 MEM_stage_inst_dmem_U19578 ( .A1(MEM_stage_inst_dmem_ram_3180), .A2(MEM_stage_inst_dmem_n20160), .ZN(MEM_stage_inst_dmem_n20137) );
NAND2_X1 MEM_stage_inst_dmem_U19577 ( .A1(MEM_stage_inst_dmem_n20135), .A2(MEM_stage_inst_dmem_n20134), .ZN(MEM_stage_inst_dmem_n9384) );
NAND2_X1 MEM_stage_inst_dmem_U19576 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n20161), .ZN(MEM_stage_inst_dmem_n20134) );
NAND2_X1 MEM_stage_inst_dmem_U19575 ( .A1(MEM_stage_inst_dmem_ram_3181), .A2(MEM_stage_inst_dmem_n20160), .ZN(MEM_stage_inst_dmem_n20135) );
NAND2_X1 MEM_stage_inst_dmem_U19574 ( .A1(MEM_stage_inst_dmem_n20133), .A2(MEM_stage_inst_dmem_n20132), .ZN(MEM_stage_inst_dmem_n9385) );
NAND2_X1 MEM_stage_inst_dmem_U19573 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n20161), .ZN(MEM_stage_inst_dmem_n20132) );
NAND2_X1 MEM_stage_inst_dmem_U19572 ( .A1(MEM_stage_inst_dmem_ram_3182), .A2(MEM_stage_inst_dmem_n20160), .ZN(MEM_stage_inst_dmem_n20133) );
NAND2_X1 MEM_stage_inst_dmem_U19571 ( .A1(MEM_stage_inst_dmem_n20131), .A2(MEM_stage_inst_dmem_n20130), .ZN(MEM_stage_inst_dmem_n9386) );
NAND2_X1 MEM_stage_inst_dmem_U19570 ( .A1(MEM_stage_inst_dmem_n14693), .A2(MEM_stage_inst_dmem_n20161), .ZN(MEM_stage_inst_dmem_n20130) );
INV_X1 MEM_stage_inst_dmem_U19569 ( .A(MEM_stage_inst_dmem_n20160), .ZN(MEM_stage_inst_dmem_n20161) );
NAND2_X1 MEM_stage_inst_dmem_U19568 ( .A1(MEM_stage_inst_dmem_ram_3183), .A2(MEM_stage_inst_dmem_n20160), .ZN(MEM_stage_inst_dmem_n20131) );
NAND2_X1 MEM_stage_inst_dmem_U19567 ( .A1(MEM_stage_inst_dmem_n21249), .A2(MEM_stage_inst_dmem_n20334), .ZN(MEM_stage_inst_dmem_n20160) );
NAND2_X1 MEM_stage_inst_dmem_U19566 ( .A1(MEM_stage_inst_dmem_n20129), .A2(MEM_stage_inst_dmem_n20128), .ZN(MEM_stage_inst_dmem_n9387) );
NAND2_X1 MEM_stage_inst_dmem_U19565 ( .A1(MEM_stage_inst_dmem_n20551), .A2(MEM_stage_inst_dmem_n20127), .ZN(MEM_stage_inst_dmem_n20128) );
NAND2_X1 MEM_stage_inst_dmem_U19564 ( .A1(MEM_stage_inst_dmem_ram_3184), .A2(MEM_stage_inst_dmem_n20126), .ZN(MEM_stage_inst_dmem_n20129) );
NAND2_X1 MEM_stage_inst_dmem_U19563 ( .A1(MEM_stage_inst_dmem_n20125), .A2(MEM_stage_inst_dmem_n20124), .ZN(MEM_stage_inst_dmem_n9388) );
NAND2_X1 MEM_stage_inst_dmem_U19562 ( .A1(MEM_stage_inst_dmem_n20547), .A2(MEM_stage_inst_dmem_n20127), .ZN(MEM_stage_inst_dmem_n20124) );
NAND2_X1 MEM_stage_inst_dmem_U19561 ( .A1(MEM_stage_inst_dmem_ram_3185), .A2(MEM_stage_inst_dmem_n20126), .ZN(MEM_stage_inst_dmem_n20125) );
NAND2_X1 MEM_stage_inst_dmem_U19560 ( .A1(MEM_stage_inst_dmem_n20123), .A2(MEM_stage_inst_dmem_n20122), .ZN(MEM_stage_inst_dmem_n9389) );
NAND2_X1 MEM_stage_inst_dmem_U19559 ( .A1(MEM_stage_inst_dmem_n20544), .A2(MEM_stage_inst_dmem_n20127), .ZN(MEM_stage_inst_dmem_n20122) );
NAND2_X1 MEM_stage_inst_dmem_U19558 ( .A1(MEM_stage_inst_dmem_ram_3186), .A2(MEM_stage_inst_dmem_n20126), .ZN(MEM_stage_inst_dmem_n20123) );
NAND2_X1 MEM_stage_inst_dmem_U19557 ( .A1(MEM_stage_inst_dmem_n20121), .A2(MEM_stage_inst_dmem_n20120), .ZN(MEM_stage_inst_dmem_n9390) );
NAND2_X1 MEM_stage_inst_dmem_U19556 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n20127), .ZN(MEM_stage_inst_dmem_n20120) );
NAND2_X1 MEM_stage_inst_dmem_U19555 ( .A1(MEM_stage_inst_dmem_ram_3187), .A2(MEM_stage_inst_dmem_n20126), .ZN(MEM_stage_inst_dmem_n20121) );
NAND2_X1 MEM_stage_inst_dmem_U19554 ( .A1(MEM_stage_inst_dmem_n20119), .A2(MEM_stage_inst_dmem_n20118), .ZN(MEM_stage_inst_dmem_n9391) );
NAND2_X1 MEM_stage_inst_dmem_U19553 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n20127), .ZN(MEM_stage_inst_dmem_n20118) );
NAND2_X1 MEM_stage_inst_dmem_U19552 ( .A1(MEM_stage_inst_dmem_ram_3188), .A2(MEM_stage_inst_dmem_n20126), .ZN(MEM_stage_inst_dmem_n20119) );
NAND2_X1 MEM_stage_inst_dmem_U19551 ( .A1(MEM_stage_inst_dmem_n20117), .A2(MEM_stage_inst_dmem_n20116), .ZN(MEM_stage_inst_dmem_n9392) );
NAND2_X1 MEM_stage_inst_dmem_U19550 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n20127), .ZN(MEM_stage_inst_dmem_n20116) );
NAND2_X1 MEM_stage_inst_dmem_U19549 ( .A1(MEM_stage_inst_dmem_ram_3189), .A2(MEM_stage_inst_dmem_n20126), .ZN(MEM_stage_inst_dmem_n20117) );
NAND2_X1 MEM_stage_inst_dmem_U19548 ( .A1(MEM_stage_inst_dmem_n20115), .A2(MEM_stage_inst_dmem_n20114), .ZN(MEM_stage_inst_dmem_n9393) );
NAND2_X1 MEM_stage_inst_dmem_U19547 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n20127), .ZN(MEM_stage_inst_dmem_n20114) );
NAND2_X1 MEM_stage_inst_dmem_U19546 ( .A1(MEM_stage_inst_dmem_ram_3190), .A2(MEM_stage_inst_dmem_n20126), .ZN(MEM_stage_inst_dmem_n20115) );
NAND2_X1 MEM_stage_inst_dmem_U19545 ( .A1(MEM_stage_inst_dmem_n20113), .A2(MEM_stage_inst_dmem_n20112), .ZN(MEM_stage_inst_dmem_n9394) );
NAND2_X1 MEM_stage_inst_dmem_U19544 ( .A1(MEM_stage_inst_dmem_n20530), .A2(MEM_stage_inst_dmem_n20127), .ZN(MEM_stage_inst_dmem_n20112) );
NAND2_X1 MEM_stage_inst_dmem_U19543 ( .A1(MEM_stage_inst_dmem_ram_3191), .A2(MEM_stage_inst_dmem_n20126), .ZN(MEM_stage_inst_dmem_n20113) );
NAND2_X1 MEM_stage_inst_dmem_U19542 ( .A1(MEM_stage_inst_dmem_n20111), .A2(MEM_stage_inst_dmem_n20110), .ZN(MEM_stage_inst_dmem_n9395) );
NAND2_X1 MEM_stage_inst_dmem_U19541 ( .A1(MEM_stage_inst_dmem_n20527), .A2(MEM_stage_inst_dmem_n20127), .ZN(MEM_stage_inst_dmem_n20110) );
NAND2_X1 MEM_stage_inst_dmem_U19540 ( .A1(MEM_stage_inst_dmem_ram_3192), .A2(MEM_stage_inst_dmem_n20126), .ZN(MEM_stage_inst_dmem_n20111) );
NAND2_X1 MEM_stage_inst_dmem_U19539 ( .A1(MEM_stage_inst_dmem_n20109), .A2(MEM_stage_inst_dmem_n20108), .ZN(MEM_stage_inst_dmem_n9396) );
NAND2_X1 MEM_stage_inst_dmem_U19538 ( .A1(MEM_stage_inst_dmem_n20524), .A2(MEM_stage_inst_dmem_n20127), .ZN(MEM_stage_inst_dmem_n20108) );
NAND2_X1 MEM_stage_inst_dmem_U19537 ( .A1(MEM_stage_inst_dmem_ram_3193), .A2(MEM_stage_inst_dmem_n20126), .ZN(MEM_stage_inst_dmem_n20109) );
NAND2_X1 MEM_stage_inst_dmem_U19536 ( .A1(MEM_stage_inst_dmem_n20107), .A2(MEM_stage_inst_dmem_n20106), .ZN(MEM_stage_inst_dmem_n9397) );
NAND2_X1 MEM_stage_inst_dmem_U19535 ( .A1(MEM_stage_inst_dmem_n20521), .A2(MEM_stage_inst_dmem_n20127), .ZN(MEM_stage_inst_dmem_n20106) );
NAND2_X1 MEM_stage_inst_dmem_U19534 ( .A1(MEM_stage_inst_dmem_ram_3194), .A2(MEM_stage_inst_dmem_n20126), .ZN(MEM_stage_inst_dmem_n20107) );
NAND2_X1 MEM_stage_inst_dmem_U19533 ( .A1(MEM_stage_inst_dmem_n20105), .A2(MEM_stage_inst_dmem_n20104), .ZN(MEM_stage_inst_dmem_n9398) );
NAND2_X1 MEM_stage_inst_dmem_U19532 ( .A1(MEM_stage_inst_dmem_n20518), .A2(MEM_stage_inst_dmem_n20127), .ZN(MEM_stage_inst_dmem_n20104) );
NAND2_X1 MEM_stage_inst_dmem_U19531 ( .A1(MEM_stage_inst_dmem_ram_3195), .A2(MEM_stage_inst_dmem_n20126), .ZN(MEM_stage_inst_dmem_n20105) );
NAND2_X1 MEM_stage_inst_dmem_U19530 ( .A1(MEM_stage_inst_dmem_n20103), .A2(MEM_stage_inst_dmem_n20102), .ZN(MEM_stage_inst_dmem_n9399) );
NAND2_X1 MEM_stage_inst_dmem_U19529 ( .A1(MEM_stage_inst_dmem_n20515), .A2(MEM_stage_inst_dmem_n20127), .ZN(MEM_stage_inst_dmem_n20102) );
NAND2_X1 MEM_stage_inst_dmem_U19528 ( .A1(MEM_stage_inst_dmem_ram_3196), .A2(MEM_stage_inst_dmem_n20126), .ZN(MEM_stage_inst_dmem_n20103) );
NAND2_X1 MEM_stage_inst_dmem_U19527 ( .A1(MEM_stage_inst_dmem_n20101), .A2(MEM_stage_inst_dmem_n20100), .ZN(MEM_stage_inst_dmem_n9400) );
NAND2_X1 MEM_stage_inst_dmem_U19526 ( .A1(MEM_stage_inst_dmem_n20512), .A2(MEM_stage_inst_dmem_n20127), .ZN(MEM_stage_inst_dmem_n20100) );
NAND2_X1 MEM_stage_inst_dmem_U19525 ( .A1(MEM_stage_inst_dmem_ram_3197), .A2(MEM_stage_inst_dmem_n20126), .ZN(MEM_stage_inst_dmem_n20101) );
NAND2_X1 MEM_stage_inst_dmem_U19524 ( .A1(MEM_stage_inst_dmem_n20099), .A2(MEM_stage_inst_dmem_n20098), .ZN(MEM_stage_inst_dmem_n9401) );
NAND2_X1 MEM_stage_inst_dmem_U19523 ( .A1(MEM_stage_inst_dmem_n20509), .A2(MEM_stage_inst_dmem_n20127), .ZN(MEM_stage_inst_dmem_n20098) );
NAND2_X1 MEM_stage_inst_dmem_U19522 ( .A1(MEM_stage_inst_dmem_ram_3198), .A2(MEM_stage_inst_dmem_n20126), .ZN(MEM_stage_inst_dmem_n20099) );
NAND2_X1 MEM_stage_inst_dmem_U19521 ( .A1(MEM_stage_inst_dmem_n20097), .A2(MEM_stage_inst_dmem_n20096), .ZN(MEM_stage_inst_dmem_n9402) );
NAND2_X1 MEM_stage_inst_dmem_U19520 ( .A1(MEM_stage_inst_dmem_n20506), .A2(MEM_stage_inst_dmem_n20127), .ZN(MEM_stage_inst_dmem_n20096) );
INV_X1 MEM_stage_inst_dmem_U19519 ( .A(MEM_stage_inst_dmem_n20126), .ZN(MEM_stage_inst_dmem_n20127) );
NAND2_X1 MEM_stage_inst_dmem_U19518 ( .A1(MEM_stage_inst_dmem_ram_3199), .A2(MEM_stage_inst_dmem_n20126), .ZN(MEM_stage_inst_dmem_n20097) );
NAND2_X1 MEM_stage_inst_dmem_U19517 ( .A1(MEM_stage_inst_dmem_n21214), .A2(MEM_stage_inst_dmem_n20334), .ZN(MEM_stage_inst_dmem_n20126) );
NAND2_X1 MEM_stage_inst_dmem_U19516 ( .A1(MEM_stage_inst_dmem_n20095), .A2(MEM_stage_inst_dmem_n20094), .ZN(MEM_stage_inst_dmem_n9403) );
NAND2_X1 MEM_stage_inst_dmem_U19515 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n20093), .ZN(MEM_stage_inst_dmem_n20094) );
NAND2_X1 MEM_stage_inst_dmem_U19514 ( .A1(MEM_stage_inst_dmem_ram_3200), .A2(MEM_stage_inst_dmem_n20092), .ZN(MEM_stage_inst_dmem_n20095) );
NAND2_X1 MEM_stage_inst_dmem_U19513 ( .A1(MEM_stage_inst_dmem_n20091), .A2(MEM_stage_inst_dmem_n20090), .ZN(MEM_stage_inst_dmem_n9404) );
NAND2_X1 MEM_stage_inst_dmem_U19512 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n20093), .ZN(MEM_stage_inst_dmem_n20090) );
NAND2_X1 MEM_stage_inst_dmem_U19511 ( .A1(MEM_stage_inst_dmem_ram_3201), .A2(MEM_stage_inst_dmem_n20092), .ZN(MEM_stage_inst_dmem_n20091) );
NAND2_X1 MEM_stage_inst_dmem_U19510 ( .A1(MEM_stage_inst_dmem_n20089), .A2(MEM_stage_inst_dmem_n20088), .ZN(MEM_stage_inst_dmem_n9405) );
NAND2_X1 MEM_stage_inst_dmem_U19509 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n20093), .ZN(MEM_stage_inst_dmem_n20088) );
NAND2_X1 MEM_stage_inst_dmem_U19508 ( .A1(MEM_stage_inst_dmem_ram_3202), .A2(MEM_stage_inst_dmem_n20092), .ZN(MEM_stage_inst_dmem_n20089) );
NAND2_X1 MEM_stage_inst_dmem_U19507 ( .A1(MEM_stage_inst_dmem_n20087), .A2(MEM_stage_inst_dmem_n20086), .ZN(MEM_stage_inst_dmem_n9406) );
NAND2_X1 MEM_stage_inst_dmem_U19506 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n20093), .ZN(MEM_stage_inst_dmem_n20086) );
NAND2_X1 MEM_stage_inst_dmem_U19505 ( .A1(MEM_stage_inst_dmem_ram_3203), .A2(MEM_stage_inst_dmem_n20092), .ZN(MEM_stage_inst_dmem_n20087) );
NAND2_X1 MEM_stage_inst_dmem_U19504 ( .A1(MEM_stage_inst_dmem_n20085), .A2(MEM_stage_inst_dmem_n20084), .ZN(MEM_stage_inst_dmem_n9407) );
NAND2_X1 MEM_stage_inst_dmem_U19503 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n20093), .ZN(MEM_stage_inst_dmem_n20084) );
NAND2_X1 MEM_stage_inst_dmem_U19502 ( .A1(MEM_stage_inst_dmem_ram_3204), .A2(MEM_stage_inst_dmem_n20092), .ZN(MEM_stage_inst_dmem_n20085) );
NAND2_X1 MEM_stage_inst_dmem_U19501 ( .A1(MEM_stage_inst_dmem_n20083), .A2(MEM_stage_inst_dmem_n20082), .ZN(MEM_stage_inst_dmem_n9408) );
NAND2_X1 MEM_stage_inst_dmem_U19500 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n20093), .ZN(MEM_stage_inst_dmem_n20082) );
NAND2_X1 MEM_stage_inst_dmem_U19499 ( .A1(MEM_stage_inst_dmem_ram_3205), .A2(MEM_stage_inst_dmem_n20092), .ZN(MEM_stage_inst_dmem_n20083) );
NAND2_X1 MEM_stage_inst_dmem_U19498 ( .A1(MEM_stage_inst_dmem_n20081), .A2(MEM_stage_inst_dmem_n20080), .ZN(MEM_stage_inst_dmem_n9409) );
NAND2_X1 MEM_stage_inst_dmem_U19497 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n20093), .ZN(MEM_stage_inst_dmem_n20080) );
NAND2_X1 MEM_stage_inst_dmem_U19496 ( .A1(MEM_stage_inst_dmem_ram_3206), .A2(MEM_stage_inst_dmem_n20092), .ZN(MEM_stage_inst_dmem_n20081) );
NAND2_X1 MEM_stage_inst_dmem_U19495 ( .A1(MEM_stage_inst_dmem_n20079), .A2(MEM_stage_inst_dmem_n20078), .ZN(MEM_stage_inst_dmem_n9410) );
NAND2_X1 MEM_stage_inst_dmem_U19494 ( .A1(MEM_stage_inst_dmem_n16361), .A2(MEM_stage_inst_dmem_n20093), .ZN(MEM_stage_inst_dmem_n20078) );
NAND2_X1 MEM_stage_inst_dmem_U19493 ( .A1(MEM_stage_inst_dmem_ram_3207), .A2(MEM_stage_inst_dmem_n20092), .ZN(MEM_stage_inst_dmem_n20079) );
NAND2_X1 MEM_stage_inst_dmem_U19492 ( .A1(MEM_stage_inst_dmem_n20077), .A2(MEM_stage_inst_dmem_n20076), .ZN(MEM_stage_inst_dmem_n9411) );
NAND2_X1 MEM_stage_inst_dmem_U19491 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n20093), .ZN(MEM_stage_inst_dmem_n20076) );
NAND2_X1 MEM_stage_inst_dmem_U19490 ( .A1(MEM_stage_inst_dmem_ram_3208), .A2(MEM_stage_inst_dmem_n20092), .ZN(MEM_stage_inst_dmem_n20077) );
NAND2_X1 MEM_stage_inst_dmem_U19489 ( .A1(MEM_stage_inst_dmem_n20075), .A2(MEM_stage_inst_dmem_n20074), .ZN(MEM_stage_inst_dmem_n9412) );
NAND2_X1 MEM_stage_inst_dmem_U19488 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n20093), .ZN(MEM_stage_inst_dmem_n20074) );
NAND2_X1 MEM_stage_inst_dmem_U19487 ( .A1(MEM_stage_inst_dmem_ram_3209), .A2(MEM_stage_inst_dmem_n20092), .ZN(MEM_stage_inst_dmem_n20075) );
NAND2_X1 MEM_stage_inst_dmem_U19486 ( .A1(MEM_stage_inst_dmem_n20073), .A2(MEM_stage_inst_dmem_n20072), .ZN(MEM_stage_inst_dmem_n9413) );
NAND2_X1 MEM_stage_inst_dmem_U19485 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n20093), .ZN(MEM_stage_inst_dmem_n20072) );
NAND2_X1 MEM_stage_inst_dmem_U19484 ( .A1(MEM_stage_inst_dmem_ram_3210), .A2(MEM_stage_inst_dmem_n20092), .ZN(MEM_stage_inst_dmem_n20073) );
NAND2_X1 MEM_stage_inst_dmem_U19483 ( .A1(MEM_stage_inst_dmem_n20071), .A2(MEM_stage_inst_dmem_n20070), .ZN(MEM_stage_inst_dmem_n9414) );
NAND2_X1 MEM_stage_inst_dmem_U19482 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n20093), .ZN(MEM_stage_inst_dmem_n20070) );
NAND2_X1 MEM_stage_inst_dmem_U19481 ( .A1(MEM_stage_inst_dmem_ram_3211), .A2(MEM_stage_inst_dmem_n20092), .ZN(MEM_stage_inst_dmem_n20071) );
NAND2_X1 MEM_stage_inst_dmem_U19480 ( .A1(MEM_stage_inst_dmem_n20069), .A2(MEM_stage_inst_dmem_n20068), .ZN(MEM_stage_inst_dmem_n9415) );
NAND2_X1 MEM_stage_inst_dmem_U19479 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n20093), .ZN(MEM_stage_inst_dmem_n20068) );
NAND2_X1 MEM_stage_inst_dmem_U19478 ( .A1(MEM_stage_inst_dmem_ram_3212), .A2(MEM_stage_inst_dmem_n20092), .ZN(MEM_stage_inst_dmem_n20069) );
NAND2_X1 MEM_stage_inst_dmem_U19477 ( .A1(MEM_stage_inst_dmem_n20067), .A2(MEM_stage_inst_dmem_n20066), .ZN(MEM_stage_inst_dmem_n9416) );
NAND2_X1 MEM_stage_inst_dmem_U19476 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n20093), .ZN(MEM_stage_inst_dmem_n20066) );
NAND2_X1 MEM_stage_inst_dmem_U19475 ( .A1(MEM_stage_inst_dmem_ram_3213), .A2(MEM_stage_inst_dmem_n20092), .ZN(MEM_stage_inst_dmem_n20067) );
NAND2_X1 MEM_stage_inst_dmem_U19474 ( .A1(MEM_stage_inst_dmem_n20065), .A2(MEM_stage_inst_dmem_n20064), .ZN(MEM_stage_inst_dmem_n9417) );
NAND2_X1 MEM_stage_inst_dmem_U19473 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n20093), .ZN(MEM_stage_inst_dmem_n20064) );
NAND2_X1 MEM_stage_inst_dmem_U19472 ( .A1(MEM_stage_inst_dmem_ram_3214), .A2(MEM_stage_inst_dmem_n20092), .ZN(MEM_stage_inst_dmem_n20065) );
NAND2_X1 MEM_stage_inst_dmem_U19471 ( .A1(MEM_stage_inst_dmem_n20063), .A2(MEM_stage_inst_dmem_n20062), .ZN(MEM_stage_inst_dmem_n9418) );
NAND2_X1 MEM_stage_inst_dmem_U19470 ( .A1(MEM_stage_inst_dmem_n16343), .A2(MEM_stage_inst_dmem_n20093), .ZN(MEM_stage_inst_dmem_n20062) );
NAND2_X1 MEM_stage_inst_dmem_U19469 ( .A1(MEM_stage_inst_dmem_ram_3215), .A2(MEM_stage_inst_dmem_n20092), .ZN(MEM_stage_inst_dmem_n20063) );
NAND2_X1 MEM_stage_inst_dmem_U19468 ( .A1(MEM_stage_inst_dmem_n21179), .A2(MEM_stage_inst_dmem_n20334), .ZN(MEM_stage_inst_dmem_n20092) );
NAND2_X1 MEM_stage_inst_dmem_U19467 ( .A1(MEM_stage_inst_dmem_n20061), .A2(MEM_stage_inst_dmem_n20060), .ZN(MEM_stage_inst_dmem_n9419) );
NAND2_X1 MEM_stage_inst_dmem_U19466 ( .A1(MEM_stage_inst_dmem_n20551), .A2(MEM_stage_inst_dmem_n20059), .ZN(MEM_stage_inst_dmem_n20060) );
NAND2_X1 MEM_stage_inst_dmem_U19465 ( .A1(MEM_stage_inst_dmem_ram_3216), .A2(MEM_stage_inst_dmem_n20058), .ZN(MEM_stage_inst_dmem_n20061) );
NAND2_X1 MEM_stage_inst_dmem_U19464 ( .A1(MEM_stage_inst_dmem_n20057), .A2(MEM_stage_inst_dmem_n20056), .ZN(MEM_stage_inst_dmem_n9420) );
NAND2_X1 MEM_stage_inst_dmem_U19463 ( .A1(MEM_stage_inst_dmem_n20547), .A2(MEM_stage_inst_dmem_n20059), .ZN(MEM_stage_inst_dmem_n20056) );
NAND2_X1 MEM_stage_inst_dmem_U19462 ( .A1(MEM_stage_inst_dmem_ram_3217), .A2(MEM_stage_inst_dmem_n20058), .ZN(MEM_stage_inst_dmem_n20057) );
NAND2_X1 MEM_stage_inst_dmem_U19461 ( .A1(MEM_stage_inst_dmem_n20055), .A2(MEM_stage_inst_dmem_n20054), .ZN(MEM_stage_inst_dmem_n9421) );
NAND2_X1 MEM_stage_inst_dmem_U19460 ( .A1(MEM_stage_inst_dmem_n20544), .A2(MEM_stage_inst_dmem_n20059), .ZN(MEM_stage_inst_dmem_n20054) );
NAND2_X1 MEM_stage_inst_dmem_U19459 ( .A1(MEM_stage_inst_dmem_ram_3218), .A2(MEM_stage_inst_dmem_n20058), .ZN(MEM_stage_inst_dmem_n20055) );
NAND2_X1 MEM_stage_inst_dmem_U19458 ( .A1(MEM_stage_inst_dmem_n20053), .A2(MEM_stage_inst_dmem_n20052), .ZN(MEM_stage_inst_dmem_n9422) );
NAND2_X1 MEM_stage_inst_dmem_U19457 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n20059), .ZN(MEM_stage_inst_dmem_n20052) );
NAND2_X1 MEM_stage_inst_dmem_U19456 ( .A1(MEM_stage_inst_dmem_ram_3219), .A2(MEM_stage_inst_dmem_n20058), .ZN(MEM_stage_inst_dmem_n20053) );
NAND2_X1 MEM_stage_inst_dmem_U19455 ( .A1(MEM_stage_inst_dmem_n20051), .A2(MEM_stage_inst_dmem_n20050), .ZN(MEM_stage_inst_dmem_n9423) );
NAND2_X1 MEM_stage_inst_dmem_U19454 ( .A1(MEM_stage_inst_dmem_n16784), .A2(MEM_stage_inst_dmem_n20059), .ZN(MEM_stage_inst_dmem_n20050) );
NAND2_X1 MEM_stage_inst_dmem_U19453 ( .A1(MEM_stage_inst_dmem_ram_3220), .A2(MEM_stage_inst_dmem_n20058), .ZN(MEM_stage_inst_dmem_n20051) );
NAND2_X1 MEM_stage_inst_dmem_U19452 ( .A1(MEM_stage_inst_dmem_n20049), .A2(MEM_stage_inst_dmem_n20048), .ZN(MEM_stage_inst_dmem_n9424) );
NAND2_X1 MEM_stage_inst_dmem_U19451 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n20059), .ZN(MEM_stage_inst_dmem_n20048) );
NAND2_X1 MEM_stage_inst_dmem_U19450 ( .A1(MEM_stage_inst_dmem_ram_3221), .A2(MEM_stage_inst_dmem_n20058), .ZN(MEM_stage_inst_dmem_n20049) );
NAND2_X1 MEM_stage_inst_dmem_U19449 ( .A1(MEM_stage_inst_dmem_n20047), .A2(MEM_stage_inst_dmem_n20046), .ZN(MEM_stage_inst_dmem_n9425) );
NAND2_X1 MEM_stage_inst_dmem_U19448 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n20059), .ZN(MEM_stage_inst_dmem_n20046) );
NAND2_X1 MEM_stage_inst_dmem_U19447 ( .A1(MEM_stage_inst_dmem_ram_3222), .A2(MEM_stage_inst_dmem_n20058), .ZN(MEM_stage_inst_dmem_n20047) );
NAND2_X1 MEM_stage_inst_dmem_U19446 ( .A1(MEM_stage_inst_dmem_n20045), .A2(MEM_stage_inst_dmem_n20044), .ZN(MEM_stage_inst_dmem_n9426) );
NAND2_X1 MEM_stage_inst_dmem_U19445 ( .A1(MEM_stage_inst_dmem_n20530), .A2(MEM_stage_inst_dmem_n20059), .ZN(MEM_stage_inst_dmem_n20044) );
NAND2_X1 MEM_stage_inst_dmem_U19444 ( .A1(MEM_stage_inst_dmem_ram_3223), .A2(MEM_stage_inst_dmem_n20058), .ZN(MEM_stage_inst_dmem_n20045) );
NAND2_X1 MEM_stage_inst_dmem_U19443 ( .A1(MEM_stage_inst_dmem_n20043), .A2(MEM_stage_inst_dmem_n20042), .ZN(MEM_stage_inst_dmem_n9427) );
NAND2_X1 MEM_stage_inst_dmem_U19442 ( .A1(MEM_stage_inst_dmem_n20527), .A2(MEM_stage_inst_dmem_n20059), .ZN(MEM_stage_inst_dmem_n20042) );
NAND2_X1 MEM_stage_inst_dmem_U19441 ( .A1(MEM_stage_inst_dmem_ram_3224), .A2(MEM_stage_inst_dmem_n20058), .ZN(MEM_stage_inst_dmem_n20043) );
NAND2_X1 MEM_stage_inst_dmem_U19440 ( .A1(MEM_stage_inst_dmem_n20041), .A2(MEM_stage_inst_dmem_n20040), .ZN(MEM_stage_inst_dmem_n9428) );
NAND2_X1 MEM_stage_inst_dmem_U19439 ( .A1(MEM_stage_inst_dmem_n20524), .A2(MEM_stage_inst_dmem_n20059), .ZN(MEM_stage_inst_dmem_n20040) );
NAND2_X1 MEM_stage_inst_dmem_U19438 ( .A1(MEM_stage_inst_dmem_ram_3225), .A2(MEM_stage_inst_dmem_n20058), .ZN(MEM_stage_inst_dmem_n20041) );
NAND2_X1 MEM_stage_inst_dmem_U19437 ( .A1(MEM_stage_inst_dmem_n20039), .A2(MEM_stage_inst_dmem_n20038), .ZN(MEM_stage_inst_dmem_n9429) );
NAND2_X1 MEM_stage_inst_dmem_U19436 ( .A1(MEM_stage_inst_dmem_n20521), .A2(MEM_stage_inst_dmem_n20059), .ZN(MEM_stage_inst_dmem_n20038) );
NAND2_X1 MEM_stage_inst_dmem_U19435 ( .A1(MEM_stage_inst_dmem_ram_3226), .A2(MEM_stage_inst_dmem_n20058), .ZN(MEM_stage_inst_dmem_n20039) );
NAND2_X1 MEM_stage_inst_dmem_U19434 ( .A1(MEM_stage_inst_dmem_n20037), .A2(MEM_stage_inst_dmem_n20036), .ZN(MEM_stage_inst_dmem_n9430) );
NAND2_X1 MEM_stage_inst_dmem_U19433 ( .A1(MEM_stage_inst_dmem_n20518), .A2(MEM_stage_inst_dmem_n20059), .ZN(MEM_stage_inst_dmem_n20036) );
NAND2_X1 MEM_stage_inst_dmem_U19432 ( .A1(MEM_stage_inst_dmem_ram_3227), .A2(MEM_stage_inst_dmem_n20058), .ZN(MEM_stage_inst_dmem_n20037) );
NAND2_X1 MEM_stage_inst_dmem_U19431 ( .A1(MEM_stage_inst_dmem_n20035), .A2(MEM_stage_inst_dmem_n20034), .ZN(MEM_stage_inst_dmem_n9431) );
NAND2_X1 MEM_stage_inst_dmem_U19430 ( .A1(MEM_stage_inst_dmem_n20515), .A2(MEM_stage_inst_dmem_n20059), .ZN(MEM_stage_inst_dmem_n20034) );
NAND2_X1 MEM_stage_inst_dmem_U19429 ( .A1(MEM_stage_inst_dmem_ram_3228), .A2(MEM_stage_inst_dmem_n20058), .ZN(MEM_stage_inst_dmem_n20035) );
NAND2_X1 MEM_stage_inst_dmem_U19428 ( .A1(MEM_stage_inst_dmem_n20033), .A2(MEM_stage_inst_dmem_n20032), .ZN(MEM_stage_inst_dmem_n9432) );
NAND2_X1 MEM_stage_inst_dmem_U19427 ( .A1(MEM_stage_inst_dmem_n20512), .A2(MEM_stage_inst_dmem_n20059), .ZN(MEM_stage_inst_dmem_n20032) );
NAND2_X1 MEM_stage_inst_dmem_U19426 ( .A1(MEM_stage_inst_dmem_ram_3229), .A2(MEM_stage_inst_dmem_n20058), .ZN(MEM_stage_inst_dmem_n20033) );
NAND2_X1 MEM_stage_inst_dmem_U19425 ( .A1(MEM_stage_inst_dmem_n20031), .A2(MEM_stage_inst_dmem_n20030), .ZN(MEM_stage_inst_dmem_n9433) );
NAND2_X1 MEM_stage_inst_dmem_U19424 ( .A1(MEM_stage_inst_dmem_n20509), .A2(MEM_stage_inst_dmem_n20059), .ZN(MEM_stage_inst_dmem_n20030) );
NAND2_X1 MEM_stage_inst_dmem_U19423 ( .A1(MEM_stage_inst_dmem_ram_3230), .A2(MEM_stage_inst_dmem_n20058), .ZN(MEM_stage_inst_dmem_n20031) );
NAND2_X1 MEM_stage_inst_dmem_U19422 ( .A1(MEM_stage_inst_dmem_n20029), .A2(MEM_stage_inst_dmem_n20028), .ZN(MEM_stage_inst_dmem_n9434) );
NAND2_X1 MEM_stage_inst_dmem_U19421 ( .A1(MEM_stage_inst_dmem_n20506), .A2(MEM_stage_inst_dmem_n20059), .ZN(MEM_stage_inst_dmem_n20028) );
INV_X1 MEM_stage_inst_dmem_U19420 ( .A(MEM_stage_inst_dmem_n20058), .ZN(MEM_stage_inst_dmem_n20059) );
NAND2_X1 MEM_stage_inst_dmem_U19419 ( .A1(MEM_stage_inst_dmem_ram_3231), .A2(MEM_stage_inst_dmem_n20058), .ZN(MEM_stage_inst_dmem_n20029) );
NAND2_X1 MEM_stage_inst_dmem_U19418 ( .A1(MEM_stage_inst_dmem_n21144), .A2(MEM_stage_inst_dmem_n20334), .ZN(MEM_stage_inst_dmem_n20058) );
NAND2_X1 MEM_stage_inst_dmem_U19417 ( .A1(MEM_stage_inst_dmem_n20027), .A2(MEM_stage_inst_dmem_n20026), .ZN(MEM_stage_inst_dmem_n9435) );
NAND2_X1 MEM_stage_inst_dmem_U19416 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n20025), .ZN(MEM_stage_inst_dmem_n20026) );
NAND2_X1 MEM_stage_inst_dmem_U19415 ( .A1(MEM_stage_inst_dmem_ram_3232), .A2(MEM_stage_inst_dmem_n20024), .ZN(MEM_stage_inst_dmem_n20027) );
NAND2_X1 MEM_stage_inst_dmem_U19414 ( .A1(MEM_stage_inst_dmem_n20023), .A2(MEM_stage_inst_dmem_n20022), .ZN(MEM_stage_inst_dmem_n9436) );
NAND2_X1 MEM_stage_inst_dmem_U19413 ( .A1(MEM_stage_inst_dmem_n109), .A2(MEM_stage_inst_dmem_n20025), .ZN(MEM_stage_inst_dmem_n20022) );
NAND2_X1 MEM_stage_inst_dmem_U19412 ( .A1(MEM_stage_inst_dmem_ram_3233), .A2(MEM_stage_inst_dmem_n20024), .ZN(MEM_stage_inst_dmem_n20023) );
NAND2_X1 MEM_stage_inst_dmem_U19411 ( .A1(MEM_stage_inst_dmem_n20021), .A2(MEM_stage_inst_dmem_n20020), .ZN(MEM_stage_inst_dmem_n9437) );
NAND2_X1 MEM_stage_inst_dmem_U19410 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n20025), .ZN(MEM_stage_inst_dmem_n20020) );
NAND2_X1 MEM_stage_inst_dmem_U19409 ( .A1(MEM_stage_inst_dmem_ram_3234), .A2(MEM_stage_inst_dmem_n20024), .ZN(MEM_stage_inst_dmem_n20021) );
NAND2_X1 MEM_stage_inst_dmem_U19408 ( .A1(MEM_stage_inst_dmem_n20019), .A2(MEM_stage_inst_dmem_n20018), .ZN(MEM_stage_inst_dmem_n9438) );
NAND2_X1 MEM_stage_inst_dmem_U19407 ( .A1(MEM_stage_inst_dmem_n13064), .A2(MEM_stage_inst_dmem_n20025), .ZN(MEM_stage_inst_dmem_n20018) );
NAND2_X1 MEM_stage_inst_dmem_U19406 ( .A1(MEM_stage_inst_dmem_ram_3235), .A2(MEM_stage_inst_dmem_n20024), .ZN(MEM_stage_inst_dmem_n20019) );
NAND2_X1 MEM_stage_inst_dmem_U19405 ( .A1(MEM_stage_inst_dmem_n20017), .A2(MEM_stage_inst_dmem_n20016), .ZN(MEM_stage_inst_dmem_n9439) );
NAND2_X1 MEM_stage_inst_dmem_U19404 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n20025), .ZN(MEM_stage_inst_dmem_n20016) );
NAND2_X1 MEM_stage_inst_dmem_U19403 ( .A1(MEM_stage_inst_dmem_ram_3236), .A2(MEM_stage_inst_dmem_n20024), .ZN(MEM_stage_inst_dmem_n20017) );
NAND2_X1 MEM_stage_inst_dmem_U19402 ( .A1(MEM_stage_inst_dmem_n20015), .A2(MEM_stage_inst_dmem_n20014), .ZN(MEM_stage_inst_dmem_n9440) );
NAND2_X1 MEM_stage_inst_dmem_U19401 ( .A1(MEM_stage_inst_dmem_n13059), .A2(MEM_stage_inst_dmem_n20025), .ZN(MEM_stage_inst_dmem_n20014) );
NAND2_X1 MEM_stage_inst_dmem_U19400 ( .A1(MEM_stage_inst_dmem_ram_3237), .A2(MEM_stage_inst_dmem_n20024), .ZN(MEM_stage_inst_dmem_n20015) );
NAND2_X1 MEM_stage_inst_dmem_U19399 ( .A1(MEM_stage_inst_dmem_n20013), .A2(MEM_stage_inst_dmem_n20012), .ZN(MEM_stage_inst_dmem_n9441) );
NAND2_X1 MEM_stage_inst_dmem_U19398 ( .A1(MEM_stage_inst_dmem_n13056), .A2(MEM_stage_inst_dmem_n20025), .ZN(MEM_stage_inst_dmem_n20012) );
NAND2_X1 MEM_stage_inst_dmem_U19397 ( .A1(MEM_stage_inst_dmem_ram_3238), .A2(MEM_stage_inst_dmem_n20024), .ZN(MEM_stage_inst_dmem_n20013) );
NAND2_X1 MEM_stage_inst_dmem_U19396 ( .A1(MEM_stage_inst_dmem_n20011), .A2(MEM_stage_inst_dmem_n20010), .ZN(MEM_stage_inst_dmem_n9442) );
NAND2_X1 MEM_stage_inst_dmem_U19395 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n20025), .ZN(MEM_stage_inst_dmem_n20010) );
NAND2_X1 MEM_stage_inst_dmem_U19394 ( .A1(MEM_stage_inst_dmem_ram_3239), .A2(MEM_stage_inst_dmem_n20024), .ZN(MEM_stage_inst_dmem_n20011) );
NAND2_X1 MEM_stage_inst_dmem_U19393 ( .A1(MEM_stage_inst_dmem_n20009), .A2(MEM_stage_inst_dmem_n20008), .ZN(MEM_stage_inst_dmem_n9443) );
NAND2_X1 MEM_stage_inst_dmem_U19392 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n20025), .ZN(MEM_stage_inst_dmem_n20008) );
NAND2_X1 MEM_stage_inst_dmem_U19391 ( .A1(MEM_stage_inst_dmem_ram_3240), .A2(MEM_stage_inst_dmem_n20024), .ZN(MEM_stage_inst_dmem_n20009) );
NAND2_X1 MEM_stage_inst_dmem_U19390 ( .A1(MEM_stage_inst_dmem_n20007), .A2(MEM_stage_inst_dmem_n20006), .ZN(MEM_stage_inst_dmem_n9444) );
NAND2_X1 MEM_stage_inst_dmem_U19389 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n20025), .ZN(MEM_stage_inst_dmem_n20006) );
NAND2_X1 MEM_stage_inst_dmem_U19388 ( .A1(MEM_stage_inst_dmem_ram_3241), .A2(MEM_stage_inst_dmem_n20024), .ZN(MEM_stage_inst_dmem_n20007) );
NAND2_X1 MEM_stage_inst_dmem_U19387 ( .A1(MEM_stage_inst_dmem_n20005), .A2(MEM_stage_inst_dmem_n20004), .ZN(MEM_stage_inst_dmem_n9445) );
NAND2_X1 MEM_stage_inst_dmem_U19386 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n20025), .ZN(MEM_stage_inst_dmem_n20004) );
NAND2_X1 MEM_stage_inst_dmem_U19385 ( .A1(MEM_stage_inst_dmem_ram_3242), .A2(MEM_stage_inst_dmem_n20024), .ZN(MEM_stage_inst_dmem_n20005) );
NAND2_X1 MEM_stage_inst_dmem_U19384 ( .A1(MEM_stage_inst_dmem_n20003), .A2(MEM_stage_inst_dmem_n20002), .ZN(MEM_stage_inst_dmem_n9446) );
NAND2_X1 MEM_stage_inst_dmem_U19383 ( .A1(MEM_stage_inst_dmem_n20904), .A2(MEM_stage_inst_dmem_n20025), .ZN(MEM_stage_inst_dmem_n20002) );
NAND2_X1 MEM_stage_inst_dmem_U19382 ( .A1(MEM_stage_inst_dmem_ram_3243), .A2(MEM_stage_inst_dmem_n20024), .ZN(MEM_stage_inst_dmem_n20003) );
NAND2_X1 MEM_stage_inst_dmem_U19381 ( .A1(MEM_stage_inst_dmem_n20001), .A2(MEM_stage_inst_dmem_n20000), .ZN(MEM_stage_inst_dmem_n9447) );
NAND2_X1 MEM_stage_inst_dmem_U19380 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n20025), .ZN(MEM_stage_inst_dmem_n20000) );
NAND2_X1 MEM_stage_inst_dmem_U19379 ( .A1(MEM_stage_inst_dmem_ram_3244), .A2(MEM_stage_inst_dmem_n20024), .ZN(MEM_stage_inst_dmem_n20001) );
NAND2_X1 MEM_stage_inst_dmem_U19378 ( .A1(MEM_stage_inst_dmem_n19999), .A2(MEM_stage_inst_dmem_n19998), .ZN(MEM_stage_inst_dmem_n9448) );
NAND2_X1 MEM_stage_inst_dmem_U19377 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n20025), .ZN(MEM_stage_inst_dmem_n19998) );
NAND2_X1 MEM_stage_inst_dmem_U19376 ( .A1(MEM_stage_inst_dmem_ram_3245), .A2(MEM_stage_inst_dmem_n20024), .ZN(MEM_stage_inst_dmem_n19999) );
NAND2_X1 MEM_stage_inst_dmem_U19375 ( .A1(MEM_stage_inst_dmem_n19997), .A2(MEM_stage_inst_dmem_n19996), .ZN(MEM_stage_inst_dmem_n9449) );
NAND2_X1 MEM_stage_inst_dmem_U19374 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n20025), .ZN(MEM_stage_inst_dmem_n19996) );
NAND2_X1 MEM_stage_inst_dmem_U19373 ( .A1(MEM_stage_inst_dmem_ram_3246), .A2(MEM_stage_inst_dmem_n20024), .ZN(MEM_stage_inst_dmem_n19997) );
NAND2_X1 MEM_stage_inst_dmem_U19372 ( .A1(MEM_stage_inst_dmem_n19995), .A2(MEM_stage_inst_dmem_n19994), .ZN(MEM_stage_inst_dmem_n9450) );
NAND2_X1 MEM_stage_inst_dmem_U19371 ( .A1(MEM_stage_inst_dmem_n15110), .A2(MEM_stage_inst_dmem_n20025), .ZN(MEM_stage_inst_dmem_n19994) );
INV_X1 MEM_stage_inst_dmem_U19370 ( .A(MEM_stage_inst_dmem_n20024), .ZN(MEM_stage_inst_dmem_n20025) );
NAND2_X1 MEM_stage_inst_dmem_U19369 ( .A1(MEM_stage_inst_dmem_ram_3247), .A2(MEM_stage_inst_dmem_n20024), .ZN(MEM_stage_inst_dmem_n19995) );
NAND2_X1 MEM_stage_inst_dmem_U19368 ( .A1(MEM_stage_inst_dmem_n21109), .A2(MEM_stage_inst_dmem_n20334), .ZN(MEM_stage_inst_dmem_n20024) );
NAND2_X1 MEM_stage_inst_dmem_U19367 ( .A1(MEM_stage_inst_dmem_n19993), .A2(MEM_stage_inst_dmem_n19992), .ZN(MEM_stage_inst_dmem_n9451) );
NAND2_X1 MEM_stage_inst_dmem_U19366 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n19991), .ZN(MEM_stage_inst_dmem_n19992) );
NAND2_X1 MEM_stage_inst_dmem_U19365 ( .A1(MEM_stage_inst_dmem_ram_3248), .A2(MEM_stage_inst_dmem_n19990), .ZN(MEM_stage_inst_dmem_n19993) );
NAND2_X1 MEM_stage_inst_dmem_U19364 ( .A1(MEM_stage_inst_dmem_n19989), .A2(MEM_stage_inst_dmem_n19988), .ZN(MEM_stage_inst_dmem_n9452) );
NAND2_X1 MEM_stage_inst_dmem_U19363 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n19991), .ZN(MEM_stage_inst_dmem_n19988) );
NAND2_X1 MEM_stage_inst_dmem_U19362 ( .A1(MEM_stage_inst_dmem_ram_3249), .A2(MEM_stage_inst_dmem_n19990), .ZN(MEM_stage_inst_dmem_n19989) );
NAND2_X1 MEM_stage_inst_dmem_U19361 ( .A1(MEM_stage_inst_dmem_n19987), .A2(MEM_stage_inst_dmem_n19986), .ZN(MEM_stage_inst_dmem_n9453) );
NAND2_X1 MEM_stage_inst_dmem_U19360 ( .A1(MEM_stage_inst_dmem_n20544), .A2(MEM_stage_inst_dmem_n19991), .ZN(MEM_stage_inst_dmem_n19986) );
NAND2_X1 MEM_stage_inst_dmem_U19359 ( .A1(MEM_stage_inst_dmem_ram_3250), .A2(MEM_stage_inst_dmem_n19990), .ZN(MEM_stage_inst_dmem_n19987) );
NAND2_X1 MEM_stage_inst_dmem_U19358 ( .A1(MEM_stage_inst_dmem_n19985), .A2(MEM_stage_inst_dmem_n19984), .ZN(MEM_stage_inst_dmem_n9454) );
NAND2_X1 MEM_stage_inst_dmem_U19357 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n19991), .ZN(MEM_stage_inst_dmem_n19984) );
NAND2_X1 MEM_stage_inst_dmem_U19356 ( .A1(MEM_stage_inst_dmem_ram_3251), .A2(MEM_stage_inst_dmem_n19990), .ZN(MEM_stage_inst_dmem_n19985) );
NAND2_X1 MEM_stage_inst_dmem_U19355 ( .A1(MEM_stage_inst_dmem_n19983), .A2(MEM_stage_inst_dmem_n19982), .ZN(MEM_stage_inst_dmem_n9455) );
NAND2_X1 MEM_stage_inst_dmem_U19354 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n19991), .ZN(MEM_stage_inst_dmem_n19982) );
NAND2_X1 MEM_stage_inst_dmem_U19353 ( .A1(MEM_stage_inst_dmem_ram_3252), .A2(MEM_stage_inst_dmem_n19990), .ZN(MEM_stage_inst_dmem_n19983) );
NAND2_X1 MEM_stage_inst_dmem_U19352 ( .A1(MEM_stage_inst_dmem_n19981), .A2(MEM_stage_inst_dmem_n19980), .ZN(MEM_stage_inst_dmem_n9456) );
NAND2_X1 MEM_stage_inst_dmem_U19351 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n19991), .ZN(MEM_stage_inst_dmem_n19980) );
NAND2_X1 MEM_stage_inst_dmem_U19350 ( .A1(MEM_stage_inst_dmem_ram_3253), .A2(MEM_stage_inst_dmem_n19990), .ZN(MEM_stage_inst_dmem_n19981) );
NAND2_X1 MEM_stage_inst_dmem_U19349 ( .A1(MEM_stage_inst_dmem_n19979), .A2(MEM_stage_inst_dmem_n19978), .ZN(MEM_stage_inst_dmem_n9457) );
NAND2_X1 MEM_stage_inst_dmem_U19348 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n19991), .ZN(MEM_stage_inst_dmem_n19978) );
NAND2_X1 MEM_stage_inst_dmem_U19347 ( .A1(MEM_stage_inst_dmem_ram_3254), .A2(MEM_stage_inst_dmem_n19990), .ZN(MEM_stage_inst_dmem_n19979) );
NAND2_X1 MEM_stage_inst_dmem_U19346 ( .A1(MEM_stage_inst_dmem_n19977), .A2(MEM_stage_inst_dmem_n19976), .ZN(MEM_stage_inst_dmem_n9458) );
NAND2_X1 MEM_stage_inst_dmem_U19345 ( .A1(MEM_stage_inst_dmem_n13886), .A2(MEM_stage_inst_dmem_n19991), .ZN(MEM_stage_inst_dmem_n19976) );
NAND2_X1 MEM_stage_inst_dmem_U19344 ( .A1(MEM_stage_inst_dmem_ram_3255), .A2(MEM_stage_inst_dmem_n19990), .ZN(MEM_stage_inst_dmem_n19977) );
NAND2_X1 MEM_stage_inst_dmem_U19343 ( .A1(MEM_stage_inst_dmem_n19975), .A2(MEM_stage_inst_dmem_n19974), .ZN(MEM_stage_inst_dmem_n9459) );
NAND2_X1 MEM_stage_inst_dmem_U19342 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n19991), .ZN(MEM_stage_inst_dmem_n19974) );
NAND2_X1 MEM_stage_inst_dmem_U19341 ( .A1(MEM_stage_inst_dmem_ram_3256), .A2(MEM_stage_inst_dmem_n19990), .ZN(MEM_stage_inst_dmem_n19975) );
NAND2_X1 MEM_stage_inst_dmem_U19340 ( .A1(MEM_stage_inst_dmem_n19973), .A2(MEM_stage_inst_dmem_n19972), .ZN(MEM_stage_inst_dmem_n9460) );
NAND2_X1 MEM_stage_inst_dmem_U19339 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n19991), .ZN(MEM_stage_inst_dmem_n19972) );
NAND2_X1 MEM_stage_inst_dmem_U19338 ( .A1(MEM_stage_inst_dmem_ram_3257), .A2(MEM_stage_inst_dmem_n19990), .ZN(MEM_stage_inst_dmem_n19973) );
NAND2_X1 MEM_stage_inst_dmem_U19337 ( .A1(MEM_stage_inst_dmem_n19971), .A2(MEM_stage_inst_dmem_n19970), .ZN(MEM_stage_inst_dmem_n9461) );
NAND2_X1 MEM_stage_inst_dmem_U19336 ( .A1(MEM_stage_inst_dmem_n20521), .A2(MEM_stage_inst_dmem_n19991), .ZN(MEM_stage_inst_dmem_n19970) );
NAND2_X1 MEM_stage_inst_dmem_U19335 ( .A1(MEM_stage_inst_dmem_ram_3258), .A2(MEM_stage_inst_dmem_n19990), .ZN(MEM_stage_inst_dmem_n19971) );
NAND2_X1 MEM_stage_inst_dmem_U19334 ( .A1(MEM_stage_inst_dmem_n19969), .A2(MEM_stage_inst_dmem_n19968), .ZN(MEM_stage_inst_dmem_n9462) );
NAND2_X1 MEM_stage_inst_dmem_U19333 ( .A1(MEM_stage_inst_dmem_n14705), .A2(MEM_stage_inst_dmem_n19991), .ZN(MEM_stage_inst_dmem_n19968) );
NAND2_X1 MEM_stage_inst_dmem_U19332 ( .A1(MEM_stage_inst_dmem_ram_3259), .A2(MEM_stage_inst_dmem_n19990), .ZN(MEM_stage_inst_dmem_n19969) );
NAND2_X1 MEM_stage_inst_dmem_U19331 ( .A1(MEM_stage_inst_dmem_n19967), .A2(MEM_stage_inst_dmem_n19966), .ZN(MEM_stage_inst_dmem_n9463) );
NAND2_X1 MEM_stage_inst_dmem_U19330 ( .A1(MEM_stage_inst_dmem_n14702), .A2(MEM_stage_inst_dmem_n19991), .ZN(MEM_stage_inst_dmem_n19966) );
NAND2_X1 MEM_stage_inst_dmem_U19329 ( .A1(MEM_stage_inst_dmem_ram_3260), .A2(MEM_stage_inst_dmem_n19990), .ZN(MEM_stage_inst_dmem_n19967) );
NAND2_X1 MEM_stage_inst_dmem_U19328 ( .A1(MEM_stage_inst_dmem_n19965), .A2(MEM_stage_inst_dmem_n19964), .ZN(MEM_stage_inst_dmem_n9464) );
NAND2_X1 MEM_stage_inst_dmem_U19327 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n19991), .ZN(MEM_stage_inst_dmem_n19964) );
NAND2_X1 MEM_stage_inst_dmem_U19326 ( .A1(MEM_stage_inst_dmem_ram_3261), .A2(MEM_stage_inst_dmem_n19990), .ZN(MEM_stage_inst_dmem_n19965) );
NAND2_X1 MEM_stage_inst_dmem_U19325 ( .A1(MEM_stage_inst_dmem_n19963), .A2(MEM_stage_inst_dmem_n19962), .ZN(MEM_stage_inst_dmem_n9465) );
NAND2_X1 MEM_stage_inst_dmem_U19324 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n19991), .ZN(MEM_stage_inst_dmem_n19962) );
NAND2_X1 MEM_stage_inst_dmem_U19323 ( .A1(MEM_stage_inst_dmem_ram_3262), .A2(MEM_stage_inst_dmem_n19990), .ZN(MEM_stage_inst_dmem_n19963) );
NAND2_X1 MEM_stage_inst_dmem_U19322 ( .A1(MEM_stage_inst_dmem_n19961), .A2(MEM_stage_inst_dmem_n19960), .ZN(MEM_stage_inst_dmem_n9466) );
NAND2_X1 MEM_stage_inst_dmem_U19321 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n19991), .ZN(MEM_stage_inst_dmem_n19960) );
INV_X1 MEM_stage_inst_dmem_U19320 ( .A(MEM_stage_inst_dmem_n19990), .ZN(MEM_stage_inst_dmem_n19991) );
NAND2_X1 MEM_stage_inst_dmem_U19319 ( .A1(MEM_stage_inst_dmem_ram_3263), .A2(MEM_stage_inst_dmem_n19990), .ZN(MEM_stage_inst_dmem_n19961) );
NAND2_X1 MEM_stage_inst_dmem_U19318 ( .A1(MEM_stage_inst_dmem_n21074), .A2(MEM_stage_inst_dmem_n20334), .ZN(MEM_stage_inst_dmem_n19990) );
NAND2_X1 MEM_stage_inst_dmem_U19317 ( .A1(MEM_stage_inst_dmem_n19959), .A2(MEM_stage_inst_dmem_n19958), .ZN(MEM_stage_inst_dmem_n9467) );
NAND2_X1 MEM_stage_inst_dmem_U19316 ( .A1(MEM_stage_inst_dmem_n20551), .A2(MEM_stage_inst_dmem_n19957), .ZN(MEM_stage_inst_dmem_n19958) );
NAND2_X1 MEM_stage_inst_dmem_U19315 ( .A1(MEM_stage_inst_dmem_ram_3264), .A2(MEM_stage_inst_dmem_n19956), .ZN(MEM_stage_inst_dmem_n19959) );
NAND2_X1 MEM_stage_inst_dmem_U19314 ( .A1(MEM_stage_inst_dmem_n19955), .A2(MEM_stage_inst_dmem_n19954), .ZN(MEM_stage_inst_dmem_n9468) );
NAND2_X1 MEM_stage_inst_dmem_U19313 ( .A1(MEM_stage_inst_dmem_n20547), .A2(MEM_stage_inst_dmem_n19957), .ZN(MEM_stage_inst_dmem_n19954) );
NAND2_X1 MEM_stage_inst_dmem_U19312 ( .A1(MEM_stage_inst_dmem_ram_3265), .A2(MEM_stage_inst_dmem_n19956), .ZN(MEM_stage_inst_dmem_n19955) );
NAND2_X1 MEM_stage_inst_dmem_U19311 ( .A1(MEM_stage_inst_dmem_n19953), .A2(MEM_stage_inst_dmem_n19952), .ZN(MEM_stage_inst_dmem_n9469) );
NAND2_X1 MEM_stage_inst_dmem_U19310 ( .A1(MEM_stage_inst_dmem_n20544), .A2(MEM_stage_inst_dmem_n19957), .ZN(MEM_stage_inst_dmem_n19952) );
NAND2_X1 MEM_stage_inst_dmem_U19309 ( .A1(MEM_stage_inst_dmem_ram_3266), .A2(MEM_stage_inst_dmem_n19956), .ZN(MEM_stage_inst_dmem_n19953) );
NAND2_X1 MEM_stage_inst_dmem_U19308 ( .A1(MEM_stage_inst_dmem_n19951), .A2(MEM_stage_inst_dmem_n19950), .ZN(MEM_stage_inst_dmem_n9470) );
NAND2_X1 MEM_stage_inst_dmem_U19307 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n19957), .ZN(MEM_stage_inst_dmem_n19950) );
NAND2_X1 MEM_stage_inst_dmem_U19306 ( .A1(MEM_stage_inst_dmem_ram_3267), .A2(MEM_stage_inst_dmem_n19956), .ZN(MEM_stage_inst_dmem_n19951) );
NAND2_X1 MEM_stage_inst_dmem_U19305 ( .A1(MEM_stage_inst_dmem_n19949), .A2(MEM_stage_inst_dmem_n19948), .ZN(MEM_stage_inst_dmem_n9471) );
NAND2_X1 MEM_stage_inst_dmem_U19304 ( .A1(EX_pipeline_reg_out_9), .A2(MEM_stage_inst_dmem_n19957), .ZN(MEM_stage_inst_dmem_n19948) );
NAND2_X1 MEM_stage_inst_dmem_U19303 ( .A1(MEM_stage_inst_dmem_ram_3268), .A2(MEM_stage_inst_dmem_n19956), .ZN(MEM_stage_inst_dmem_n19949) );
NAND2_X1 MEM_stage_inst_dmem_U19302 ( .A1(MEM_stage_inst_dmem_n19947), .A2(MEM_stage_inst_dmem_n19946), .ZN(MEM_stage_inst_dmem_n9472) );
NAND2_X1 MEM_stage_inst_dmem_U19301 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n19957), .ZN(MEM_stage_inst_dmem_n19946) );
NAND2_X1 MEM_stage_inst_dmem_U19300 ( .A1(MEM_stage_inst_dmem_ram_3269), .A2(MEM_stage_inst_dmem_n19956), .ZN(MEM_stage_inst_dmem_n19947) );
NAND2_X1 MEM_stage_inst_dmem_U19299 ( .A1(MEM_stage_inst_dmem_n19945), .A2(MEM_stage_inst_dmem_n19944), .ZN(MEM_stage_inst_dmem_n9473) );
NAND2_X1 MEM_stage_inst_dmem_U19298 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n19957), .ZN(MEM_stage_inst_dmem_n19944) );
NAND2_X1 MEM_stage_inst_dmem_U19297 ( .A1(MEM_stage_inst_dmem_ram_3270), .A2(MEM_stage_inst_dmem_n19956), .ZN(MEM_stage_inst_dmem_n19945) );
NAND2_X1 MEM_stage_inst_dmem_U19296 ( .A1(MEM_stage_inst_dmem_n19943), .A2(MEM_stage_inst_dmem_n19942), .ZN(MEM_stage_inst_dmem_n9474) );
NAND2_X1 MEM_stage_inst_dmem_U19295 ( .A1(MEM_stage_inst_dmem_n20530), .A2(MEM_stage_inst_dmem_n19957), .ZN(MEM_stage_inst_dmem_n19942) );
NAND2_X1 MEM_stage_inst_dmem_U19294 ( .A1(MEM_stage_inst_dmem_ram_3271), .A2(MEM_stage_inst_dmem_n19956), .ZN(MEM_stage_inst_dmem_n19943) );
NAND2_X1 MEM_stage_inst_dmem_U19293 ( .A1(MEM_stage_inst_dmem_n19941), .A2(MEM_stage_inst_dmem_n19940), .ZN(MEM_stage_inst_dmem_n9475) );
NAND2_X1 MEM_stage_inst_dmem_U19292 ( .A1(MEM_stage_inst_dmem_n20527), .A2(MEM_stage_inst_dmem_n19957), .ZN(MEM_stage_inst_dmem_n19940) );
NAND2_X1 MEM_stage_inst_dmem_U19291 ( .A1(MEM_stage_inst_dmem_ram_3272), .A2(MEM_stage_inst_dmem_n19956), .ZN(MEM_stage_inst_dmem_n19941) );
NAND2_X1 MEM_stage_inst_dmem_U19290 ( .A1(MEM_stage_inst_dmem_n19939), .A2(MEM_stage_inst_dmem_n19938), .ZN(MEM_stage_inst_dmem_n9476) );
NAND2_X1 MEM_stage_inst_dmem_U19289 ( .A1(MEM_stage_inst_dmem_n20524), .A2(MEM_stage_inst_dmem_n19957), .ZN(MEM_stage_inst_dmem_n19938) );
NAND2_X1 MEM_stage_inst_dmem_U19288 ( .A1(MEM_stage_inst_dmem_ram_3273), .A2(MEM_stage_inst_dmem_n19956), .ZN(MEM_stage_inst_dmem_n19939) );
NAND2_X1 MEM_stage_inst_dmem_U19287 ( .A1(MEM_stage_inst_dmem_n19937), .A2(MEM_stage_inst_dmem_n19936), .ZN(MEM_stage_inst_dmem_n9477) );
NAND2_X1 MEM_stage_inst_dmem_U19286 ( .A1(MEM_stage_inst_dmem_n20521), .A2(MEM_stage_inst_dmem_n19957), .ZN(MEM_stage_inst_dmem_n19936) );
NAND2_X1 MEM_stage_inst_dmem_U19285 ( .A1(MEM_stage_inst_dmem_ram_3274), .A2(MEM_stage_inst_dmem_n19956), .ZN(MEM_stage_inst_dmem_n19937) );
NAND2_X1 MEM_stage_inst_dmem_U19284 ( .A1(MEM_stage_inst_dmem_n19935), .A2(MEM_stage_inst_dmem_n19934), .ZN(MEM_stage_inst_dmem_n9478) );
NAND2_X1 MEM_stage_inst_dmem_U19283 ( .A1(MEM_stage_inst_dmem_n20518), .A2(MEM_stage_inst_dmem_n19957), .ZN(MEM_stage_inst_dmem_n19934) );
NAND2_X1 MEM_stage_inst_dmem_U19282 ( .A1(MEM_stage_inst_dmem_ram_3275), .A2(MEM_stage_inst_dmem_n19956), .ZN(MEM_stage_inst_dmem_n19935) );
NAND2_X1 MEM_stage_inst_dmem_U19281 ( .A1(MEM_stage_inst_dmem_n19933), .A2(MEM_stage_inst_dmem_n19932), .ZN(MEM_stage_inst_dmem_n9479) );
NAND2_X1 MEM_stage_inst_dmem_U19280 ( .A1(MEM_stage_inst_dmem_n20515), .A2(MEM_stage_inst_dmem_n19957), .ZN(MEM_stage_inst_dmem_n19932) );
NAND2_X1 MEM_stage_inst_dmem_U19279 ( .A1(MEM_stage_inst_dmem_ram_3276), .A2(MEM_stage_inst_dmem_n19956), .ZN(MEM_stage_inst_dmem_n19933) );
NAND2_X1 MEM_stage_inst_dmem_U19278 ( .A1(MEM_stage_inst_dmem_n19931), .A2(MEM_stage_inst_dmem_n19930), .ZN(MEM_stage_inst_dmem_n9480) );
NAND2_X1 MEM_stage_inst_dmem_U19277 ( .A1(MEM_stage_inst_dmem_n20512), .A2(MEM_stage_inst_dmem_n19957), .ZN(MEM_stage_inst_dmem_n19930) );
NAND2_X1 MEM_stage_inst_dmem_U19276 ( .A1(MEM_stage_inst_dmem_ram_3277), .A2(MEM_stage_inst_dmem_n19956), .ZN(MEM_stage_inst_dmem_n19931) );
NAND2_X1 MEM_stage_inst_dmem_U19275 ( .A1(MEM_stage_inst_dmem_n19929), .A2(MEM_stage_inst_dmem_n19928), .ZN(MEM_stage_inst_dmem_n9481) );
NAND2_X1 MEM_stage_inst_dmem_U19274 ( .A1(MEM_stage_inst_dmem_n20509), .A2(MEM_stage_inst_dmem_n19957), .ZN(MEM_stage_inst_dmem_n19928) );
NAND2_X1 MEM_stage_inst_dmem_U19273 ( .A1(MEM_stage_inst_dmem_ram_3278), .A2(MEM_stage_inst_dmem_n19956), .ZN(MEM_stage_inst_dmem_n19929) );
NAND2_X1 MEM_stage_inst_dmem_U19272 ( .A1(MEM_stage_inst_dmem_n19927), .A2(MEM_stage_inst_dmem_n19926), .ZN(MEM_stage_inst_dmem_n9482) );
NAND2_X1 MEM_stage_inst_dmem_U19271 ( .A1(MEM_stage_inst_dmem_n20506), .A2(MEM_stage_inst_dmem_n19957), .ZN(MEM_stage_inst_dmem_n19926) );
INV_X1 MEM_stage_inst_dmem_U19270 ( .A(MEM_stage_inst_dmem_n19956), .ZN(MEM_stage_inst_dmem_n19957) );
NAND2_X1 MEM_stage_inst_dmem_U19269 ( .A1(MEM_stage_inst_dmem_ram_3279), .A2(MEM_stage_inst_dmem_n19956), .ZN(MEM_stage_inst_dmem_n19927) );
NAND2_X1 MEM_stage_inst_dmem_U19268 ( .A1(MEM_stage_inst_dmem_n21039), .A2(MEM_stage_inst_dmem_n20334), .ZN(MEM_stage_inst_dmem_n19956) );
NAND2_X1 MEM_stage_inst_dmem_U19267 ( .A1(MEM_stage_inst_dmem_n19925), .A2(MEM_stage_inst_dmem_n19924), .ZN(MEM_stage_inst_dmem_n9483) );
NAND2_X1 MEM_stage_inst_dmem_U19266 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n19923), .ZN(MEM_stage_inst_dmem_n19924) );
NAND2_X1 MEM_stage_inst_dmem_U19265 ( .A1(MEM_stage_inst_dmem_ram_3280), .A2(MEM_stage_inst_dmem_n19922), .ZN(MEM_stage_inst_dmem_n19925) );
NAND2_X1 MEM_stage_inst_dmem_U19264 ( .A1(MEM_stage_inst_dmem_n19921), .A2(MEM_stage_inst_dmem_n19920), .ZN(MEM_stage_inst_dmem_n9484) );
NAND2_X1 MEM_stage_inst_dmem_U19263 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n19923), .ZN(MEM_stage_inst_dmem_n19920) );
NAND2_X1 MEM_stage_inst_dmem_U19262 ( .A1(MEM_stage_inst_dmem_ram_3281), .A2(MEM_stage_inst_dmem_n19922), .ZN(MEM_stage_inst_dmem_n19921) );
NAND2_X1 MEM_stage_inst_dmem_U19261 ( .A1(MEM_stage_inst_dmem_n19919), .A2(MEM_stage_inst_dmem_n19918), .ZN(MEM_stage_inst_dmem_n9485) );
NAND2_X1 MEM_stage_inst_dmem_U19260 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n19923), .ZN(MEM_stage_inst_dmem_n19918) );
NAND2_X1 MEM_stage_inst_dmem_U19259 ( .A1(MEM_stage_inst_dmem_ram_3282), .A2(MEM_stage_inst_dmem_n19922), .ZN(MEM_stage_inst_dmem_n19919) );
NAND2_X1 MEM_stage_inst_dmem_U19258 ( .A1(MEM_stage_inst_dmem_n19917), .A2(MEM_stage_inst_dmem_n19916), .ZN(MEM_stage_inst_dmem_n9486) );
NAND2_X1 MEM_stage_inst_dmem_U19257 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n19923), .ZN(MEM_stage_inst_dmem_n19916) );
NAND2_X1 MEM_stage_inst_dmem_U19256 ( .A1(MEM_stage_inst_dmem_ram_3283), .A2(MEM_stage_inst_dmem_n19922), .ZN(MEM_stage_inst_dmem_n19917) );
NAND2_X1 MEM_stage_inst_dmem_U19255 ( .A1(MEM_stage_inst_dmem_n19915), .A2(MEM_stage_inst_dmem_n19914), .ZN(MEM_stage_inst_dmem_n9487) );
NAND2_X1 MEM_stage_inst_dmem_U19254 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n19923), .ZN(MEM_stage_inst_dmem_n19914) );
NAND2_X1 MEM_stage_inst_dmem_U19253 ( .A1(MEM_stage_inst_dmem_ram_3284), .A2(MEM_stage_inst_dmem_n19922), .ZN(MEM_stage_inst_dmem_n19915) );
NAND2_X1 MEM_stage_inst_dmem_U19252 ( .A1(MEM_stage_inst_dmem_n19913), .A2(MEM_stage_inst_dmem_n19912), .ZN(MEM_stage_inst_dmem_n9488) );
NAND2_X1 MEM_stage_inst_dmem_U19251 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n19923), .ZN(MEM_stage_inst_dmem_n19912) );
NAND2_X1 MEM_stage_inst_dmem_U19250 ( .A1(MEM_stage_inst_dmem_ram_3285), .A2(MEM_stage_inst_dmem_n19922), .ZN(MEM_stage_inst_dmem_n19913) );
NAND2_X1 MEM_stage_inst_dmem_U19249 ( .A1(MEM_stage_inst_dmem_n19911), .A2(MEM_stage_inst_dmem_n19910), .ZN(MEM_stage_inst_dmem_n9489) );
NAND2_X1 MEM_stage_inst_dmem_U19248 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n19923), .ZN(MEM_stage_inst_dmem_n19910) );
NAND2_X1 MEM_stage_inst_dmem_U19247 ( .A1(MEM_stage_inst_dmem_ram_3286), .A2(MEM_stage_inst_dmem_n19922), .ZN(MEM_stage_inst_dmem_n19911) );
NAND2_X1 MEM_stage_inst_dmem_U19246 ( .A1(MEM_stage_inst_dmem_n19909), .A2(MEM_stage_inst_dmem_n19908), .ZN(MEM_stage_inst_dmem_n9490) );
NAND2_X1 MEM_stage_inst_dmem_U19245 ( .A1(EX_pipeline_reg_out_12), .A2(MEM_stage_inst_dmem_n19923), .ZN(MEM_stage_inst_dmem_n19908) );
NAND2_X1 MEM_stage_inst_dmem_U19244 ( .A1(MEM_stage_inst_dmem_ram_3287), .A2(MEM_stage_inst_dmem_n19922), .ZN(MEM_stage_inst_dmem_n19909) );
NAND2_X1 MEM_stage_inst_dmem_U19243 ( .A1(MEM_stage_inst_dmem_n19907), .A2(MEM_stage_inst_dmem_n19906), .ZN(MEM_stage_inst_dmem_n9491) );
NAND2_X1 MEM_stage_inst_dmem_U19242 ( .A1(MEM_stage_inst_dmem_n13883), .A2(MEM_stage_inst_dmem_n19923), .ZN(MEM_stage_inst_dmem_n19906) );
NAND2_X1 MEM_stage_inst_dmem_U19241 ( .A1(MEM_stage_inst_dmem_ram_3288), .A2(MEM_stage_inst_dmem_n19922), .ZN(MEM_stage_inst_dmem_n19907) );
NAND2_X1 MEM_stage_inst_dmem_U19240 ( .A1(MEM_stage_inst_dmem_n19905), .A2(MEM_stage_inst_dmem_n19904), .ZN(MEM_stage_inst_dmem_n9492) );
NAND2_X1 MEM_stage_inst_dmem_U19239 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n19923), .ZN(MEM_stage_inst_dmem_n19904) );
NAND2_X1 MEM_stage_inst_dmem_U19238 ( .A1(MEM_stage_inst_dmem_ram_3289), .A2(MEM_stage_inst_dmem_n19922), .ZN(MEM_stage_inst_dmem_n19905) );
NAND2_X1 MEM_stage_inst_dmem_U19237 ( .A1(MEM_stage_inst_dmem_n19903), .A2(MEM_stage_inst_dmem_n19902), .ZN(MEM_stage_inst_dmem_n9493) );
NAND2_X1 MEM_stage_inst_dmem_U19236 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n19923), .ZN(MEM_stage_inst_dmem_n19902) );
NAND2_X1 MEM_stage_inst_dmem_U19235 ( .A1(MEM_stage_inst_dmem_ram_3290), .A2(MEM_stage_inst_dmem_n19922), .ZN(MEM_stage_inst_dmem_n19903) );
NAND2_X1 MEM_stage_inst_dmem_U19234 ( .A1(MEM_stage_inst_dmem_n19901), .A2(MEM_stage_inst_dmem_n19900), .ZN(MEM_stage_inst_dmem_n9494) );
NAND2_X1 MEM_stage_inst_dmem_U19233 ( .A1(MEM_stage_inst_dmem_n13044), .A2(MEM_stage_inst_dmem_n19923), .ZN(MEM_stage_inst_dmem_n19900) );
NAND2_X1 MEM_stage_inst_dmem_U19232 ( .A1(MEM_stage_inst_dmem_ram_3291), .A2(MEM_stage_inst_dmem_n19922), .ZN(MEM_stage_inst_dmem_n19901) );
NAND2_X1 MEM_stage_inst_dmem_U19231 ( .A1(MEM_stage_inst_dmem_n19899), .A2(MEM_stage_inst_dmem_n19898), .ZN(MEM_stage_inst_dmem_n9495) );
NAND2_X1 MEM_stage_inst_dmem_U19230 ( .A1(MEM_stage_inst_dmem_n13041), .A2(MEM_stage_inst_dmem_n19923), .ZN(MEM_stage_inst_dmem_n19898) );
NAND2_X1 MEM_stage_inst_dmem_U19229 ( .A1(MEM_stage_inst_dmem_ram_3292), .A2(MEM_stage_inst_dmem_n19922), .ZN(MEM_stage_inst_dmem_n19899) );
NAND2_X1 MEM_stage_inst_dmem_U19228 ( .A1(MEM_stage_inst_dmem_n19897), .A2(MEM_stage_inst_dmem_n19896), .ZN(MEM_stage_inst_dmem_n9496) );
NAND2_X1 MEM_stage_inst_dmem_U19227 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n19923), .ZN(MEM_stage_inst_dmem_n19896) );
NAND2_X1 MEM_stage_inst_dmem_U19226 ( .A1(MEM_stage_inst_dmem_ram_3293), .A2(MEM_stage_inst_dmem_n19922), .ZN(MEM_stage_inst_dmem_n19897) );
NAND2_X1 MEM_stage_inst_dmem_U19225 ( .A1(MEM_stage_inst_dmem_n19895), .A2(MEM_stage_inst_dmem_n19894), .ZN(MEM_stage_inst_dmem_n9497) );
NAND2_X1 MEM_stage_inst_dmem_U19224 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n19923), .ZN(MEM_stage_inst_dmem_n19894) );
NAND2_X1 MEM_stage_inst_dmem_U19223 ( .A1(MEM_stage_inst_dmem_ram_3294), .A2(MEM_stage_inst_dmem_n19922), .ZN(MEM_stage_inst_dmem_n19895) );
NAND2_X1 MEM_stage_inst_dmem_U19222 ( .A1(MEM_stage_inst_dmem_n19893), .A2(MEM_stage_inst_dmem_n19892), .ZN(MEM_stage_inst_dmem_n9498) );
NAND2_X1 MEM_stage_inst_dmem_U19221 ( .A1(MEM_stage_inst_dmem_n15110), .A2(MEM_stage_inst_dmem_n19923), .ZN(MEM_stage_inst_dmem_n19892) );
INV_X1 MEM_stage_inst_dmem_U19220 ( .A(MEM_stage_inst_dmem_n19922), .ZN(MEM_stage_inst_dmem_n19923) );
NAND2_X1 MEM_stage_inst_dmem_U19219 ( .A1(MEM_stage_inst_dmem_ram_3295), .A2(MEM_stage_inst_dmem_n19922), .ZN(MEM_stage_inst_dmem_n19893) );
NAND2_X1 MEM_stage_inst_dmem_U19218 ( .A1(MEM_stage_inst_dmem_n21004), .A2(MEM_stage_inst_dmem_n20334), .ZN(MEM_stage_inst_dmem_n19922) );
NAND2_X1 MEM_stage_inst_dmem_U19217 ( .A1(MEM_stage_inst_dmem_n19891), .A2(MEM_stage_inst_dmem_n19890), .ZN(MEM_stage_inst_dmem_n9499) );
NAND2_X1 MEM_stage_inst_dmem_U19216 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n19889), .ZN(MEM_stage_inst_dmem_n19890) );
NAND2_X1 MEM_stage_inst_dmem_U19215 ( .A1(MEM_stage_inst_dmem_ram_3296), .A2(MEM_stage_inst_dmem_n19888), .ZN(MEM_stage_inst_dmem_n19891) );
NAND2_X1 MEM_stage_inst_dmem_U19214 ( .A1(MEM_stage_inst_dmem_n19887), .A2(MEM_stage_inst_dmem_n19886), .ZN(MEM_stage_inst_dmem_n9500) );
NAND2_X1 MEM_stage_inst_dmem_U19213 ( .A1(EX_pipeline_reg_out_6), .A2(MEM_stage_inst_dmem_n19889), .ZN(MEM_stage_inst_dmem_n19886) );
NAND2_X1 MEM_stage_inst_dmem_U19212 ( .A1(MEM_stage_inst_dmem_ram_3297), .A2(MEM_stage_inst_dmem_n19888), .ZN(MEM_stage_inst_dmem_n19887) );
NAND2_X1 MEM_stage_inst_dmem_U19211 ( .A1(MEM_stage_inst_dmem_n19885), .A2(MEM_stage_inst_dmem_n19884), .ZN(MEM_stage_inst_dmem_n9501) );
NAND2_X1 MEM_stage_inst_dmem_U19210 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n19889), .ZN(MEM_stage_inst_dmem_n19884) );
NAND2_X1 MEM_stage_inst_dmem_U19209 ( .A1(MEM_stage_inst_dmem_ram_3298), .A2(MEM_stage_inst_dmem_n19888), .ZN(MEM_stage_inst_dmem_n19885) );
NAND2_X1 MEM_stage_inst_dmem_U19208 ( .A1(MEM_stage_inst_dmem_n19883), .A2(MEM_stage_inst_dmem_n19882), .ZN(MEM_stage_inst_dmem_n9502) );
NAND2_X1 MEM_stage_inst_dmem_U19207 ( .A1(EX_pipeline_reg_out_8), .A2(MEM_stage_inst_dmem_n19889), .ZN(MEM_stage_inst_dmem_n19882) );
NAND2_X1 MEM_stage_inst_dmem_U19206 ( .A1(MEM_stage_inst_dmem_ram_3299), .A2(MEM_stage_inst_dmem_n19888), .ZN(MEM_stage_inst_dmem_n19883) );
NAND2_X1 MEM_stage_inst_dmem_U19205 ( .A1(MEM_stage_inst_dmem_n19881), .A2(MEM_stage_inst_dmem_n19880), .ZN(MEM_stage_inst_dmem_n9503) );
NAND2_X1 MEM_stage_inst_dmem_U19204 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n19889), .ZN(MEM_stage_inst_dmem_n19880) );
NAND2_X1 MEM_stage_inst_dmem_U19203 ( .A1(MEM_stage_inst_dmem_ram_3300), .A2(MEM_stage_inst_dmem_n19888), .ZN(MEM_stage_inst_dmem_n19881) );
NAND2_X1 MEM_stage_inst_dmem_U19202 ( .A1(MEM_stage_inst_dmem_n19879), .A2(MEM_stage_inst_dmem_n19878), .ZN(MEM_stage_inst_dmem_n9504) );
NAND2_X1 MEM_stage_inst_dmem_U19201 ( .A1(EX_pipeline_reg_out_10), .A2(MEM_stage_inst_dmem_n19889), .ZN(MEM_stage_inst_dmem_n19878) );
NAND2_X1 MEM_stage_inst_dmem_U19200 ( .A1(MEM_stage_inst_dmem_ram_3301), .A2(MEM_stage_inst_dmem_n19888), .ZN(MEM_stage_inst_dmem_n19879) );
NAND2_X1 MEM_stage_inst_dmem_U19199 ( .A1(MEM_stage_inst_dmem_n19877), .A2(MEM_stage_inst_dmem_n19876), .ZN(MEM_stage_inst_dmem_n9505) );
NAND2_X1 MEM_stage_inst_dmem_U19198 ( .A1(MEM_stage_inst_dmem_n21340), .A2(MEM_stage_inst_dmem_n19889), .ZN(MEM_stage_inst_dmem_n19876) );
NAND2_X1 MEM_stage_inst_dmem_U19197 ( .A1(MEM_stage_inst_dmem_ram_3302), .A2(MEM_stage_inst_dmem_n19888), .ZN(MEM_stage_inst_dmem_n19877) );
NAND2_X1 MEM_stage_inst_dmem_U19196 ( .A1(MEM_stage_inst_dmem_n19875), .A2(MEM_stage_inst_dmem_n19874), .ZN(MEM_stage_inst_dmem_n9506) );
NAND2_X1 MEM_stage_inst_dmem_U19195 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n19889), .ZN(MEM_stage_inst_dmem_n19874) );
NAND2_X1 MEM_stage_inst_dmem_U19194 ( .A1(MEM_stage_inst_dmem_ram_3303), .A2(MEM_stage_inst_dmem_n19888), .ZN(MEM_stage_inst_dmem_n19875) );
NAND2_X1 MEM_stage_inst_dmem_U19193 ( .A1(MEM_stage_inst_dmem_n19873), .A2(MEM_stage_inst_dmem_n19872), .ZN(MEM_stage_inst_dmem_n9507) );
NAND2_X1 MEM_stage_inst_dmem_U19192 ( .A1(MEM_stage_inst_dmem_n13051), .A2(MEM_stage_inst_dmem_n19889), .ZN(MEM_stage_inst_dmem_n19872) );
NAND2_X1 MEM_stage_inst_dmem_U19191 ( .A1(MEM_stage_inst_dmem_ram_3304), .A2(MEM_stage_inst_dmem_n19888), .ZN(MEM_stage_inst_dmem_n19873) );
NAND2_X1 MEM_stage_inst_dmem_U19190 ( .A1(MEM_stage_inst_dmem_n19871), .A2(MEM_stage_inst_dmem_n19870), .ZN(MEM_stage_inst_dmem_n9508) );
NAND2_X1 MEM_stage_inst_dmem_U19189 ( .A1(MEM_stage_inst_dmem_n16772), .A2(MEM_stage_inst_dmem_n19889), .ZN(MEM_stage_inst_dmem_n19870) );
NAND2_X1 MEM_stage_inst_dmem_U19188 ( .A1(MEM_stage_inst_dmem_ram_3305), .A2(MEM_stage_inst_dmem_n19888), .ZN(MEM_stage_inst_dmem_n19871) );
NAND2_X1 MEM_stage_inst_dmem_U19187 ( .A1(MEM_stage_inst_dmem_n19869), .A2(MEM_stage_inst_dmem_n19868), .ZN(MEM_stage_inst_dmem_n9509) );
NAND2_X1 MEM_stage_inst_dmem_U19186 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n19889), .ZN(MEM_stage_inst_dmem_n19868) );
NAND2_X1 MEM_stage_inst_dmem_U19185 ( .A1(MEM_stage_inst_dmem_ram_3306), .A2(MEM_stage_inst_dmem_n19888), .ZN(MEM_stage_inst_dmem_n19869) );
NAND2_X1 MEM_stage_inst_dmem_U19184 ( .A1(MEM_stage_inst_dmem_n19867), .A2(MEM_stage_inst_dmem_n19866), .ZN(MEM_stage_inst_dmem_n9510) );
NAND2_X1 MEM_stage_inst_dmem_U19183 ( .A1(MEM_stage_inst_dmem_n13044), .A2(MEM_stage_inst_dmem_n19889), .ZN(MEM_stage_inst_dmem_n19866) );
NAND2_X1 MEM_stage_inst_dmem_U19182 ( .A1(MEM_stage_inst_dmem_ram_3307), .A2(MEM_stage_inst_dmem_n19888), .ZN(MEM_stage_inst_dmem_n19867) );
NAND2_X1 MEM_stage_inst_dmem_U19181 ( .A1(MEM_stage_inst_dmem_n19865), .A2(MEM_stage_inst_dmem_n19864), .ZN(MEM_stage_inst_dmem_n9511) );
NAND2_X1 MEM_stage_inst_dmem_U19180 ( .A1(MEM_stage_inst_dmem_n14702), .A2(MEM_stage_inst_dmem_n19889), .ZN(MEM_stage_inst_dmem_n19864) );
NAND2_X1 MEM_stage_inst_dmem_U19179 ( .A1(MEM_stage_inst_dmem_ram_3308), .A2(MEM_stage_inst_dmem_n19888), .ZN(MEM_stage_inst_dmem_n19865) );
NAND2_X1 MEM_stage_inst_dmem_U19178 ( .A1(MEM_stage_inst_dmem_n19863), .A2(MEM_stage_inst_dmem_n19862), .ZN(MEM_stage_inst_dmem_n9512) );
NAND2_X1 MEM_stage_inst_dmem_U19177 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n19889), .ZN(MEM_stage_inst_dmem_n19862) );
NAND2_X1 MEM_stage_inst_dmem_U19176 ( .A1(MEM_stage_inst_dmem_ram_3309), .A2(MEM_stage_inst_dmem_n19888), .ZN(MEM_stage_inst_dmem_n19863) );
NAND2_X1 MEM_stage_inst_dmem_U19175 ( .A1(MEM_stage_inst_dmem_n19861), .A2(MEM_stage_inst_dmem_n19860), .ZN(MEM_stage_inst_dmem_n9513) );
NAND2_X1 MEM_stage_inst_dmem_U19174 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n19889), .ZN(MEM_stage_inst_dmem_n19860) );
NAND2_X1 MEM_stage_inst_dmem_U19173 ( .A1(MEM_stage_inst_dmem_ram_3310), .A2(MEM_stage_inst_dmem_n19888), .ZN(MEM_stage_inst_dmem_n19861) );
NAND2_X1 MEM_stage_inst_dmem_U19172 ( .A1(MEM_stage_inst_dmem_n19859), .A2(MEM_stage_inst_dmem_n19858), .ZN(MEM_stage_inst_dmem_n9514) );
NAND2_X1 MEM_stage_inst_dmem_U19171 ( .A1(MEM_stage_inst_dmem_n14693), .A2(MEM_stage_inst_dmem_n19889), .ZN(MEM_stage_inst_dmem_n19858) );
INV_X1 MEM_stage_inst_dmem_U19170 ( .A(MEM_stage_inst_dmem_n19888), .ZN(MEM_stage_inst_dmem_n19889) );
NAND2_X1 MEM_stage_inst_dmem_U19169 ( .A1(MEM_stage_inst_dmem_ram_3311), .A2(MEM_stage_inst_dmem_n19888), .ZN(MEM_stage_inst_dmem_n19859) );
NAND2_X1 MEM_stage_inst_dmem_U19168 ( .A1(MEM_stage_inst_dmem_n20969), .A2(MEM_stage_inst_dmem_n20334), .ZN(MEM_stage_inst_dmem_n19888) );
NAND2_X1 MEM_stage_inst_dmem_U19167 ( .A1(MEM_stage_inst_dmem_n19857), .A2(MEM_stage_inst_dmem_n19856), .ZN(MEM_stage_inst_dmem_n9515) );
NAND2_X1 MEM_stage_inst_dmem_U19166 ( .A1(MEM_stage_inst_dmem_n20551), .A2(MEM_stage_inst_dmem_n19855), .ZN(MEM_stage_inst_dmem_n19856) );
NAND2_X1 MEM_stage_inst_dmem_U19165 ( .A1(MEM_stage_inst_dmem_ram_3312), .A2(MEM_stage_inst_dmem_n19854), .ZN(MEM_stage_inst_dmem_n19857) );
NAND2_X1 MEM_stage_inst_dmem_U19164 ( .A1(MEM_stage_inst_dmem_n19853), .A2(MEM_stage_inst_dmem_n19852), .ZN(MEM_stage_inst_dmem_n9516) );
NAND2_X1 MEM_stage_inst_dmem_U19163 ( .A1(MEM_stage_inst_dmem_n20547), .A2(MEM_stage_inst_dmem_n19855), .ZN(MEM_stage_inst_dmem_n19852) );
NAND2_X1 MEM_stage_inst_dmem_U19162 ( .A1(MEM_stage_inst_dmem_ram_3313), .A2(MEM_stage_inst_dmem_n19854), .ZN(MEM_stage_inst_dmem_n19853) );
NAND2_X1 MEM_stage_inst_dmem_U19161 ( .A1(MEM_stage_inst_dmem_n19851), .A2(MEM_stage_inst_dmem_n19850), .ZN(MEM_stage_inst_dmem_n9517) );
NAND2_X1 MEM_stage_inst_dmem_U19160 ( .A1(MEM_stage_inst_dmem_n20544), .A2(MEM_stage_inst_dmem_n19855), .ZN(MEM_stage_inst_dmem_n19850) );
NAND2_X1 MEM_stage_inst_dmem_U19159 ( .A1(MEM_stage_inst_dmem_ram_3314), .A2(MEM_stage_inst_dmem_n19854), .ZN(MEM_stage_inst_dmem_n19851) );
NAND2_X1 MEM_stage_inst_dmem_U19158 ( .A1(MEM_stage_inst_dmem_n19849), .A2(MEM_stage_inst_dmem_n19848), .ZN(MEM_stage_inst_dmem_n9518) );
NAND2_X1 MEM_stage_inst_dmem_U19157 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n19855), .ZN(MEM_stage_inst_dmem_n19848) );
NAND2_X1 MEM_stage_inst_dmem_U19156 ( .A1(MEM_stage_inst_dmem_ram_3315), .A2(MEM_stage_inst_dmem_n19854), .ZN(MEM_stage_inst_dmem_n19849) );
NAND2_X1 MEM_stage_inst_dmem_U19155 ( .A1(MEM_stage_inst_dmem_n19847), .A2(MEM_stage_inst_dmem_n19846), .ZN(MEM_stage_inst_dmem_n9519) );
NAND2_X1 MEM_stage_inst_dmem_U19154 ( .A1(EX_pipeline_reg_out_9), .A2(MEM_stage_inst_dmem_n19855), .ZN(MEM_stage_inst_dmem_n19846) );
NAND2_X1 MEM_stage_inst_dmem_U19153 ( .A1(MEM_stage_inst_dmem_ram_3316), .A2(MEM_stage_inst_dmem_n19854), .ZN(MEM_stage_inst_dmem_n19847) );
NAND2_X1 MEM_stage_inst_dmem_U19152 ( .A1(MEM_stage_inst_dmem_n19845), .A2(MEM_stage_inst_dmem_n19844), .ZN(MEM_stage_inst_dmem_n9520) );
NAND2_X1 MEM_stage_inst_dmem_U19151 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n19855), .ZN(MEM_stage_inst_dmem_n19844) );
NAND2_X1 MEM_stage_inst_dmem_U19150 ( .A1(MEM_stage_inst_dmem_ram_3317), .A2(MEM_stage_inst_dmem_n19854), .ZN(MEM_stage_inst_dmem_n19845) );
NAND2_X1 MEM_stage_inst_dmem_U19149 ( .A1(MEM_stage_inst_dmem_n19843), .A2(MEM_stage_inst_dmem_n19842), .ZN(MEM_stage_inst_dmem_n9521) );
NAND2_X1 MEM_stage_inst_dmem_U19148 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n19855), .ZN(MEM_stage_inst_dmem_n19842) );
NAND2_X1 MEM_stage_inst_dmem_U19147 ( .A1(MEM_stage_inst_dmem_ram_3318), .A2(MEM_stage_inst_dmem_n19854), .ZN(MEM_stage_inst_dmem_n19843) );
NAND2_X1 MEM_stage_inst_dmem_U19146 ( .A1(MEM_stage_inst_dmem_n19841), .A2(MEM_stage_inst_dmem_n19840), .ZN(MEM_stage_inst_dmem_n9522) );
NAND2_X1 MEM_stage_inst_dmem_U19145 ( .A1(MEM_stage_inst_dmem_n20530), .A2(MEM_stage_inst_dmem_n19855), .ZN(MEM_stage_inst_dmem_n19840) );
NAND2_X1 MEM_stage_inst_dmem_U19144 ( .A1(MEM_stage_inst_dmem_ram_3319), .A2(MEM_stage_inst_dmem_n19854), .ZN(MEM_stage_inst_dmem_n19841) );
NAND2_X1 MEM_stage_inst_dmem_U19143 ( .A1(MEM_stage_inst_dmem_n19839), .A2(MEM_stage_inst_dmem_n19838), .ZN(MEM_stage_inst_dmem_n9523) );
NAND2_X1 MEM_stage_inst_dmem_U19142 ( .A1(MEM_stage_inst_dmem_n20527), .A2(MEM_stage_inst_dmem_n19855), .ZN(MEM_stage_inst_dmem_n19838) );
NAND2_X1 MEM_stage_inst_dmem_U19141 ( .A1(MEM_stage_inst_dmem_ram_3320), .A2(MEM_stage_inst_dmem_n19854), .ZN(MEM_stage_inst_dmem_n19839) );
NAND2_X1 MEM_stage_inst_dmem_U19140 ( .A1(MEM_stage_inst_dmem_n19837), .A2(MEM_stage_inst_dmem_n19836), .ZN(MEM_stage_inst_dmem_n9524) );
NAND2_X1 MEM_stage_inst_dmem_U19139 ( .A1(MEM_stage_inst_dmem_n20524), .A2(MEM_stage_inst_dmem_n19855), .ZN(MEM_stage_inst_dmem_n19836) );
NAND2_X1 MEM_stage_inst_dmem_U19138 ( .A1(MEM_stage_inst_dmem_ram_3321), .A2(MEM_stage_inst_dmem_n19854), .ZN(MEM_stage_inst_dmem_n19837) );
NAND2_X1 MEM_stage_inst_dmem_U19137 ( .A1(MEM_stage_inst_dmem_n19835), .A2(MEM_stage_inst_dmem_n19834), .ZN(MEM_stage_inst_dmem_n9525) );
NAND2_X1 MEM_stage_inst_dmem_U19136 ( .A1(MEM_stage_inst_dmem_n20521), .A2(MEM_stage_inst_dmem_n19855), .ZN(MEM_stage_inst_dmem_n19834) );
NAND2_X1 MEM_stage_inst_dmem_U19135 ( .A1(MEM_stage_inst_dmem_ram_3322), .A2(MEM_stage_inst_dmem_n19854), .ZN(MEM_stage_inst_dmem_n19835) );
NAND2_X1 MEM_stage_inst_dmem_U19134 ( .A1(MEM_stage_inst_dmem_n19833), .A2(MEM_stage_inst_dmem_n19832), .ZN(MEM_stage_inst_dmem_n9526) );
NAND2_X1 MEM_stage_inst_dmem_U19133 ( .A1(MEM_stage_inst_dmem_n20518), .A2(MEM_stage_inst_dmem_n19855), .ZN(MEM_stage_inst_dmem_n19832) );
NAND2_X1 MEM_stage_inst_dmem_U19132 ( .A1(MEM_stage_inst_dmem_ram_3323), .A2(MEM_stage_inst_dmem_n19854), .ZN(MEM_stage_inst_dmem_n19833) );
NAND2_X1 MEM_stage_inst_dmem_U19131 ( .A1(MEM_stage_inst_dmem_n19831), .A2(MEM_stage_inst_dmem_n19830), .ZN(MEM_stage_inst_dmem_n9527) );
NAND2_X1 MEM_stage_inst_dmem_U19130 ( .A1(MEM_stage_inst_dmem_n20515), .A2(MEM_stage_inst_dmem_n19855), .ZN(MEM_stage_inst_dmem_n19830) );
NAND2_X1 MEM_stage_inst_dmem_U19129 ( .A1(MEM_stage_inst_dmem_ram_3324), .A2(MEM_stage_inst_dmem_n19854), .ZN(MEM_stage_inst_dmem_n19831) );
NAND2_X1 MEM_stage_inst_dmem_U19128 ( .A1(MEM_stage_inst_dmem_n19829), .A2(MEM_stage_inst_dmem_n19828), .ZN(MEM_stage_inst_dmem_n9528) );
NAND2_X1 MEM_stage_inst_dmem_U19127 ( .A1(MEM_stage_inst_dmem_n20512), .A2(MEM_stage_inst_dmem_n19855), .ZN(MEM_stage_inst_dmem_n19828) );
NAND2_X1 MEM_stage_inst_dmem_U19126 ( .A1(MEM_stage_inst_dmem_ram_3325), .A2(MEM_stage_inst_dmem_n19854), .ZN(MEM_stage_inst_dmem_n19829) );
NAND2_X1 MEM_stage_inst_dmem_U19125 ( .A1(MEM_stage_inst_dmem_n19827), .A2(MEM_stage_inst_dmem_n19826), .ZN(MEM_stage_inst_dmem_n9529) );
NAND2_X1 MEM_stage_inst_dmem_U19124 ( .A1(MEM_stage_inst_dmem_n20509), .A2(MEM_stage_inst_dmem_n19855), .ZN(MEM_stage_inst_dmem_n19826) );
NAND2_X1 MEM_stage_inst_dmem_U19123 ( .A1(MEM_stage_inst_dmem_ram_3326), .A2(MEM_stage_inst_dmem_n19854), .ZN(MEM_stage_inst_dmem_n19827) );
NAND2_X1 MEM_stage_inst_dmem_U19122 ( .A1(MEM_stage_inst_dmem_n19825), .A2(MEM_stage_inst_dmem_n19824), .ZN(MEM_stage_inst_dmem_n9530) );
NAND2_X1 MEM_stage_inst_dmem_U19121 ( .A1(MEM_stage_inst_dmem_n20506), .A2(MEM_stage_inst_dmem_n19855), .ZN(MEM_stage_inst_dmem_n19824) );
NAND2_X1 MEM_stage_inst_dmem_U19120 ( .A1(MEM_stage_inst_dmem_ram_3327), .A2(MEM_stage_inst_dmem_n19854), .ZN(MEM_stage_inst_dmem_n19825) );
NAND2_X1 MEM_stage_inst_dmem_U19119 ( .A1(MEM_stage_inst_dmem_n20934), .A2(MEM_stage_inst_dmem_n20334), .ZN(MEM_stage_inst_dmem_n19854) );
NOR2_X2 MEM_stage_inst_dmem_U19118 ( .A1(MEM_stage_inst_dmem_n19823), .A2(MEM_stage_inst_dmem_n20932), .ZN(MEM_stage_inst_dmem_n20334) );
NAND2_X1 MEM_stage_inst_dmem_U19117 ( .A1(MEM_stage_inst_dmem_n19822), .A2(MEM_stage_inst_dmem_n19821), .ZN(MEM_stage_inst_dmem_n9531) );
NAND2_X1 MEM_stage_inst_dmem_U19116 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n19820), .ZN(MEM_stage_inst_dmem_n19821) );
NAND2_X1 MEM_stage_inst_dmem_U19115 ( .A1(MEM_stage_inst_dmem_ram_3328), .A2(MEM_stage_inst_dmem_n19819), .ZN(MEM_stage_inst_dmem_n19822) );
NAND2_X1 MEM_stage_inst_dmem_U19114 ( .A1(MEM_stage_inst_dmem_n19818), .A2(MEM_stage_inst_dmem_n19817), .ZN(MEM_stage_inst_dmem_n9532) );
NAND2_X1 MEM_stage_inst_dmem_U19113 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n19820), .ZN(MEM_stage_inst_dmem_n19817) );
NAND2_X1 MEM_stage_inst_dmem_U19112 ( .A1(MEM_stage_inst_dmem_ram_3329), .A2(MEM_stage_inst_dmem_n19819), .ZN(MEM_stage_inst_dmem_n19818) );
NAND2_X1 MEM_stage_inst_dmem_U19111 ( .A1(MEM_stage_inst_dmem_n19816), .A2(MEM_stage_inst_dmem_n19815), .ZN(MEM_stage_inst_dmem_n9533) );
NAND2_X1 MEM_stage_inst_dmem_U19110 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n19820), .ZN(MEM_stage_inst_dmem_n19815) );
NAND2_X1 MEM_stage_inst_dmem_U19109 ( .A1(MEM_stage_inst_dmem_ram_3330), .A2(MEM_stage_inst_dmem_n19819), .ZN(MEM_stage_inst_dmem_n19816) );
NAND2_X1 MEM_stage_inst_dmem_U19108 ( .A1(MEM_stage_inst_dmem_n19814), .A2(MEM_stage_inst_dmem_n19813), .ZN(MEM_stage_inst_dmem_n9534) );
NAND2_X1 MEM_stage_inst_dmem_U19107 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n19820), .ZN(MEM_stage_inst_dmem_n19813) );
NAND2_X1 MEM_stage_inst_dmem_U19106 ( .A1(MEM_stage_inst_dmem_ram_3331), .A2(MEM_stage_inst_dmem_n19819), .ZN(MEM_stage_inst_dmem_n19814) );
NAND2_X1 MEM_stage_inst_dmem_U19105 ( .A1(MEM_stage_inst_dmem_n19812), .A2(MEM_stage_inst_dmem_n19811), .ZN(MEM_stage_inst_dmem_n9535) );
NAND2_X1 MEM_stage_inst_dmem_U19104 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n19820), .ZN(MEM_stage_inst_dmem_n19811) );
NAND2_X1 MEM_stage_inst_dmem_U19103 ( .A1(MEM_stage_inst_dmem_ram_3332), .A2(MEM_stage_inst_dmem_n19819), .ZN(MEM_stage_inst_dmem_n19812) );
NAND2_X1 MEM_stage_inst_dmem_U19102 ( .A1(MEM_stage_inst_dmem_n19810), .A2(MEM_stage_inst_dmem_n19809), .ZN(MEM_stage_inst_dmem_n9536) );
NAND2_X1 MEM_stage_inst_dmem_U19101 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n19820), .ZN(MEM_stage_inst_dmem_n19809) );
NAND2_X1 MEM_stage_inst_dmem_U19100 ( .A1(MEM_stage_inst_dmem_ram_3333), .A2(MEM_stage_inst_dmem_n19819), .ZN(MEM_stage_inst_dmem_n19810) );
NAND2_X1 MEM_stage_inst_dmem_U19099 ( .A1(MEM_stage_inst_dmem_n19808), .A2(MEM_stage_inst_dmem_n19807), .ZN(MEM_stage_inst_dmem_n9537) );
NAND2_X1 MEM_stage_inst_dmem_U19098 ( .A1(MEM_stage_inst_dmem_n13056), .A2(MEM_stage_inst_dmem_n19820), .ZN(MEM_stage_inst_dmem_n19807) );
NAND2_X1 MEM_stage_inst_dmem_U19097 ( .A1(MEM_stage_inst_dmem_ram_3334), .A2(MEM_stage_inst_dmem_n19819), .ZN(MEM_stage_inst_dmem_n19808) );
NAND2_X1 MEM_stage_inst_dmem_U19096 ( .A1(MEM_stage_inst_dmem_n19806), .A2(MEM_stage_inst_dmem_n19805), .ZN(MEM_stage_inst_dmem_n9538) );
NAND2_X1 MEM_stage_inst_dmem_U19095 ( .A1(MEM_stage_inst_dmem_n17), .A2(MEM_stage_inst_dmem_n19820), .ZN(MEM_stage_inst_dmem_n19805) );
NAND2_X1 MEM_stage_inst_dmem_U19094 ( .A1(MEM_stage_inst_dmem_ram_3335), .A2(MEM_stage_inst_dmem_n19819), .ZN(MEM_stage_inst_dmem_n19806) );
NAND2_X1 MEM_stage_inst_dmem_U19093 ( .A1(MEM_stage_inst_dmem_n19804), .A2(MEM_stage_inst_dmem_n19803), .ZN(MEM_stage_inst_dmem_n9539) );
NAND2_X1 MEM_stage_inst_dmem_U19092 ( .A1(EX_pipeline_reg_out_13), .A2(MEM_stage_inst_dmem_n19820), .ZN(MEM_stage_inst_dmem_n19803) );
NAND2_X1 MEM_stage_inst_dmem_U19091 ( .A1(MEM_stage_inst_dmem_ram_3336), .A2(MEM_stage_inst_dmem_n19819), .ZN(MEM_stage_inst_dmem_n19804) );
NAND2_X1 MEM_stage_inst_dmem_U19090 ( .A1(MEM_stage_inst_dmem_n19802), .A2(MEM_stage_inst_dmem_n19801), .ZN(MEM_stage_inst_dmem_n9540) );
NAND2_X1 MEM_stage_inst_dmem_U19089 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n19820), .ZN(MEM_stage_inst_dmem_n19801) );
NAND2_X1 MEM_stage_inst_dmem_U19088 ( .A1(MEM_stage_inst_dmem_ram_3337), .A2(MEM_stage_inst_dmem_n19819), .ZN(MEM_stage_inst_dmem_n19802) );
NAND2_X1 MEM_stage_inst_dmem_U19087 ( .A1(MEM_stage_inst_dmem_n19800), .A2(MEM_stage_inst_dmem_n19799), .ZN(MEM_stage_inst_dmem_n9541) );
NAND2_X1 MEM_stage_inst_dmem_U19086 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n19820), .ZN(MEM_stage_inst_dmem_n19799) );
NAND2_X1 MEM_stage_inst_dmem_U19085 ( .A1(MEM_stage_inst_dmem_ram_3338), .A2(MEM_stage_inst_dmem_n19819), .ZN(MEM_stage_inst_dmem_n19800) );
NAND2_X1 MEM_stage_inst_dmem_U19084 ( .A1(MEM_stage_inst_dmem_n19798), .A2(MEM_stage_inst_dmem_n19797), .ZN(MEM_stage_inst_dmem_n9542) );
NAND2_X1 MEM_stage_inst_dmem_U19083 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n19820), .ZN(MEM_stage_inst_dmem_n19797) );
NAND2_X1 MEM_stage_inst_dmem_U19082 ( .A1(MEM_stage_inst_dmem_ram_3339), .A2(MEM_stage_inst_dmem_n19819), .ZN(MEM_stage_inst_dmem_n19798) );
NAND2_X1 MEM_stage_inst_dmem_U19081 ( .A1(MEM_stage_inst_dmem_n19796), .A2(MEM_stage_inst_dmem_n19795), .ZN(MEM_stage_inst_dmem_n9543) );
NAND2_X1 MEM_stage_inst_dmem_U19080 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n19820), .ZN(MEM_stage_inst_dmem_n19795) );
NAND2_X1 MEM_stage_inst_dmem_U19079 ( .A1(MEM_stage_inst_dmem_ram_3340), .A2(MEM_stage_inst_dmem_n19819), .ZN(MEM_stage_inst_dmem_n19796) );
NAND2_X1 MEM_stage_inst_dmem_U19078 ( .A1(MEM_stage_inst_dmem_n19794), .A2(MEM_stage_inst_dmem_n19793), .ZN(MEM_stage_inst_dmem_n9544) );
NAND2_X1 MEM_stage_inst_dmem_U19077 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n19820), .ZN(MEM_stage_inst_dmem_n19793) );
NAND2_X1 MEM_stage_inst_dmem_U19076 ( .A1(MEM_stage_inst_dmem_ram_3341), .A2(MEM_stage_inst_dmem_n19819), .ZN(MEM_stage_inst_dmem_n19794) );
NAND2_X1 MEM_stage_inst_dmem_U19075 ( .A1(MEM_stage_inst_dmem_n19792), .A2(MEM_stage_inst_dmem_n19791), .ZN(MEM_stage_inst_dmem_n9545) );
NAND2_X1 MEM_stage_inst_dmem_U19074 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n19820), .ZN(MEM_stage_inst_dmem_n19791) );
NAND2_X1 MEM_stage_inst_dmem_U19073 ( .A1(MEM_stage_inst_dmem_ram_3342), .A2(MEM_stage_inst_dmem_n19819), .ZN(MEM_stage_inst_dmem_n19792) );
NAND2_X1 MEM_stage_inst_dmem_U19072 ( .A1(MEM_stage_inst_dmem_n19790), .A2(MEM_stage_inst_dmem_n19789), .ZN(MEM_stage_inst_dmem_n9546) );
NAND2_X1 MEM_stage_inst_dmem_U19071 ( .A1(MEM_stage_inst_dmem_n14693), .A2(MEM_stage_inst_dmem_n19820), .ZN(MEM_stage_inst_dmem_n19789) );
INV_X1 MEM_stage_inst_dmem_U19070 ( .A(MEM_stage_inst_dmem_n19819), .ZN(MEM_stage_inst_dmem_n19820) );
NAND2_X1 MEM_stage_inst_dmem_U19069 ( .A1(MEM_stage_inst_dmem_ram_3343), .A2(MEM_stage_inst_dmem_n19819), .ZN(MEM_stage_inst_dmem_n19790) );
NAND2_X1 MEM_stage_inst_dmem_U19068 ( .A1(MEM_stage_inst_dmem_n21465), .A2(MEM_stage_inst_dmem_n19788), .ZN(MEM_stage_inst_dmem_n19819) );
NAND2_X1 MEM_stage_inst_dmem_U19067 ( .A1(MEM_stage_inst_dmem_n19787), .A2(MEM_stage_inst_dmem_n19786), .ZN(MEM_stage_inst_dmem_n9547) );
NAND2_X1 MEM_stage_inst_dmem_U19066 ( .A1(MEM_stage_inst_dmem_n20551), .A2(MEM_stage_inst_dmem_n19785), .ZN(MEM_stage_inst_dmem_n19786) );
NAND2_X1 MEM_stage_inst_dmem_U19065 ( .A1(MEM_stage_inst_dmem_ram_3344), .A2(MEM_stage_inst_dmem_n19784), .ZN(MEM_stage_inst_dmem_n19787) );
NAND2_X1 MEM_stage_inst_dmem_U19064 ( .A1(MEM_stage_inst_dmem_n19783), .A2(MEM_stage_inst_dmem_n19782), .ZN(MEM_stage_inst_dmem_n9548) );
NAND2_X1 MEM_stage_inst_dmem_U19063 ( .A1(MEM_stage_inst_dmem_n20547), .A2(MEM_stage_inst_dmem_n19785), .ZN(MEM_stage_inst_dmem_n19782) );
NAND2_X1 MEM_stage_inst_dmem_U19062 ( .A1(MEM_stage_inst_dmem_ram_3345), .A2(MEM_stage_inst_dmem_n19784), .ZN(MEM_stage_inst_dmem_n19783) );
NAND2_X1 MEM_stage_inst_dmem_U19061 ( .A1(MEM_stage_inst_dmem_n19781), .A2(MEM_stage_inst_dmem_n19780), .ZN(MEM_stage_inst_dmem_n9549) );
NAND2_X1 MEM_stage_inst_dmem_U19060 ( .A1(MEM_stage_inst_dmem_n20544), .A2(MEM_stage_inst_dmem_n19785), .ZN(MEM_stage_inst_dmem_n19780) );
NAND2_X1 MEM_stage_inst_dmem_U19059 ( .A1(MEM_stage_inst_dmem_ram_3346), .A2(MEM_stage_inst_dmem_n19784), .ZN(MEM_stage_inst_dmem_n19781) );
NAND2_X1 MEM_stage_inst_dmem_U19058 ( .A1(MEM_stage_inst_dmem_n19779), .A2(MEM_stage_inst_dmem_n19778), .ZN(MEM_stage_inst_dmem_n9550) );
NAND2_X1 MEM_stage_inst_dmem_U19057 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n19785), .ZN(MEM_stage_inst_dmem_n19778) );
NAND2_X1 MEM_stage_inst_dmem_U19056 ( .A1(MEM_stage_inst_dmem_ram_3347), .A2(MEM_stage_inst_dmem_n19784), .ZN(MEM_stage_inst_dmem_n19779) );
NAND2_X1 MEM_stage_inst_dmem_U19055 ( .A1(MEM_stage_inst_dmem_n19777), .A2(MEM_stage_inst_dmem_n19776), .ZN(MEM_stage_inst_dmem_n9551) );
NAND2_X1 MEM_stage_inst_dmem_U19054 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n19785), .ZN(MEM_stage_inst_dmem_n19776) );
NAND2_X1 MEM_stage_inst_dmem_U19053 ( .A1(MEM_stage_inst_dmem_ram_3348), .A2(MEM_stage_inst_dmem_n19784), .ZN(MEM_stage_inst_dmem_n19777) );
NAND2_X1 MEM_stage_inst_dmem_U19052 ( .A1(MEM_stage_inst_dmem_n19775), .A2(MEM_stage_inst_dmem_n19774), .ZN(MEM_stage_inst_dmem_n9552) );
NAND2_X1 MEM_stage_inst_dmem_U19051 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n19785), .ZN(MEM_stage_inst_dmem_n19774) );
NAND2_X1 MEM_stage_inst_dmem_U19050 ( .A1(MEM_stage_inst_dmem_ram_3349), .A2(MEM_stage_inst_dmem_n19784), .ZN(MEM_stage_inst_dmem_n19775) );
NAND2_X1 MEM_stage_inst_dmem_U19049 ( .A1(MEM_stage_inst_dmem_n19773), .A2(MEM_stage_inst_dmem_n19772), .ZN(MEM_stage_inst_dmem_n9553) );
NAND2_X1 MEM_stage_inst_dmem_U19048 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n19785), .ZN(MEM_stage_inst_dmem_n19772) );
NAND2_X1 MEM_stage_inst_dmem_U19047 ( .A1(MEM_stage_inst_dmem_ram_3350), .A2(MEM_stage_inst_dmem_n19784), .ZN(MEM_stage_inst_dmem_n19773) );
NAND2_X1 MEM_stage_inst_dmem_U19046 ( .A1(MEM_stage_inst_dmem_n19771), .A2(MEM_stage_inst_dmem_n19770), .ZN(MEM_stage_inst_dmem_n9554) );
NAND2_X1 MEM_stage_inst_dmem_U19045 ( .A1(MEM_stage_inst_dmem_n20530), .A2(MEM_stage_inst_dmem_n19785), .ZN(MEM_stage_inst_dmem_n19770) );
NAND2_X1 MEM_stage_inst_dmem_U19044 ( .A1(MEM_stage_inst_dmem_ram_3351), .A2(MEM_stage_inst_dmem_n19784), .ZN(MEM_stage_inst_dmem_n19771) );
NAND2_X1 MEM_stage_inst_dmem_U19043 ( .A1(MEM_stage_inst_dmem_n19769), .A2(MEM_stage_inst_dmem_n19768), .ZN(MEM_stage_inst_dmem_n9555) );
NAND2_X1 MEM_stage_inst_dmem_U19042 ( .A1(MEM_stage_inst_dmem_n20527), .A2(MEM_stage_inst_dmem_n19785), .ZN(MEM_stage_inst_dmem_n19768) );
NAND2_X1 MEM_stage_inst_dmem_U19041 ( .A1(MEM_stage_inst_dmem_ram_3352), .A2(MEM_stage_inst_dmem_n19784), .ZN(MEM_stage_inst_dmem_n19769) );
NAND2_X1 MEM_stage_inst_dmem_U19040 ( .A1(MEM_stage_inst_dmem_n19767), .A2(MEM_stage_inst_dmem_n19766), .ZN(MEM_stage_inst_dmem_n9556) );
NAND2_X1 MEM_stage_inst_dmem_U19039 ( .A1(MEM_stage_inst_dmem_n20524), .A2(MEM_stage_inst_dmem_n19785), .ZN(MEM_stage_inst_dmem_n19766) );
NAND2_X1 MEM_stage_inst_dmem_U19038 ( .A1(MEM_stage_inst_dmem_ram_3353), .A2(MEM_stage_inst_dmem_n19784), .ZN(MEM_stage_inst_dmem_n19767) );
NAND2_X1 MEM_stage_inst_dmem_U19037 ( .A1(MEM_stage_inst_dmem_n19765), .A2(MEM_stage_inst_dmem_n19764), .ZN(MEM_stage_inst_dmem_n9557) );
NAND2_X1 MEM_stage_inst_dmem_U19036 ( .A1(MEM_stage_inst_dmem_n20521), .A2(MEM_stage_inst_dmem_n19785), .ZN(MEM_stage_inst_dmem_n19764) );
NAND2_X1 MEM_stage_inst_dmem_U19035 ( .A1(MEM_stage_inst_dmem_ram_3354), .A2(MEM_stage_inst_dmem_n19784), .ZN(MEM_stage_inst_dmem_n19765) );
NAND2_X1 MEM_stage_inst_dmem_U19034 ( .A1(MEM_stage_inst_dmem_n19763), .A2(MEM_stage_inst_dmem_n19762), .ZN(MEM_stage_inst_dmem_n9558) );
NAND2_X1 MEM_stage_inst_dmem_U19033 ( .A1(MEM_stage_inst_dmem_n20518), .A2(MEM_stage_inst_dmem_n19785), .ZN(MEM_stage_inst_dmem_n19762) );
NAND2_X1 MEM_stage_inst_dmem_U19032 ( .A1(MEM_stage_inst_dmem_ram_3355), .A2(MEM_stage_inst_dmem_n19784), .ZN(MEM_stage_inst_dmem_n19763) );
NAND2_X1 MEM_stage_inst_dmem_U19031 ( .A1(MEM_stage_inst_dmem_n19761), .A2(MEM_stage_inst_dmem_n19760), .ZN(MEM_stage_inst_dmem_n9559) );
NAND2_X1 MEM_stage_inst_dmem_U19030 ( .A1(MEM_stage_inst_dmem_n20515), .A2(MEM_stage_inst_dmem_n19785), .ZN(MEM_stage_inst_dmem_n19760) );
NAND2_X1 MEM_stage_inst_dmem_U19029 ( .A1(MEM_stage_inst_dmem_ram_3356), .A2(MEM_stage_inst_dmem_n19784), .ZN(MEM_stage_inst_dmem_n19761) );
NAND2_X1 MEM_stage_inst_dmem_U19028 ( .A1(MEM_stage_inst_dmem_n19759), .A2(MEM_stage_inst_dmem_n19758), .ZN(MEM_stage_inst_dmem_n9560) );
NAND2_X1 MEM_stage_inst_dmem_U19027 ( .A1(MEM_stage_inst_dmem_n20512), .A2(MEM_stage_inst_dmem_n19785), .ZN(MEM_stage_inst_dmem_n19758) );
NAND2_X1 MEM_stage_inst_dmem_U19026 ( .A1(MEM_stage_inst_dmem_ram_3357), .A2(MEM_stage_inst_dmem_n19784), .ZN(MEM_stage_inst_dmem_n19759) );
NAND2_X1 MEM_stage_inst_dmem_U19025 ( .A1(MEM_stage_inst_dmem_n19757), .A2(MEM_stage_inst_dmem_n19756), .ZN(MEM_stage_inst_dmem_n9561) );
NAND2_X1 MEM_stage_inst_dmem_U19024 ( .A1(MEM_stage_inst_dmem_n20509), .A2(MEM_stage_inst_dmem_n19785), .ZN(MEM_stage_inst_dmem_n19756) );
NAND2_X1 MEM_stage_inst_dmem_U19023 ( .A1(MEM_stage_inst_dmem_ram_3358), .A2(MEM_stage_inst_dmem_n19784), .ZN(MEM_stage_inst_dmem_n19757) );
NAND2_X1 MEM_stage_inst_dmem_U19022 ( .A1(MEM_stage_inst_dmem_n19755), .A2(MEM_stage_inst_dmem_n19754), .ZN(MEM_stage_inst_dmem_n9562) );
NAND2_X1 MEM_stage_inst_dmem_U19021 ( .A1(MEM_stage_inst_dmem_n20506), .A2(MEM_stage_inst_dmem_n19785), .ZN(MEM_stage_inst_dmem_n19754) );
INV_X1 MEM_stage_inst_dmem_U19020 ( .A(MEM_stage_inst_dmem_n19784), .ZN(MEM_stage_inst_dmem_n19785) );
NAND2_X1 MEM_stage_inst_dmem_U19019 ( .A1(MEM_stage_inst_dmem_ram_3359), .A2(MEM_stage_inst_dmem_n19784), .ZN(MEM_stage_inst_dmem_n19755) );
NAND2_X1 MEM_stage_inst_dmem_U19018 ( .A1(MEM_stage_inst_dmem_n21429), .A2(MEM_stage_inst_dmem_n19788), .ZN(MEM_stage_inst_dmem_n19784) );
NAND2_X1 MEM_stage_inst_dmem_U19017 ( .A1(MEM_stage_inst_dmem_n19753), .A2(MEM_stage_inst_dmem_n19752), .ZN(MEM_stage_inst_dmem_n9563) );
NAND2_X1 MEM_stage_inst_dmem_U19016 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n19751), .ZN(MEM_stage_inst_dmem_n19752) );
NAND2_X1 MEM_stage_inst_dmem_U19015 ( .A1(MEM_stage_inst_dmem_ram_3360), .A2(MEM_stage_inst_dmem_n19750), .ZN(MEM_stage_inst_dmem_n19753) );
NAND2_X1 MEM_stage_inst_dmem_U19014 ( .A1(MEM_stage_inst_dmem_n19749), .A2(MEM_stage_inst_dmem_n19748), .ZN(MEM_stage_inst_dmem_n9564) );
NAND2_X1 MEM_stage_inst_dmem_U19013 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n19751), .ZN(MEM_stage_inst_dmem_n19748) );
NAND2_X1 MEM_stage_inst_dmem_U19012 ( .A1(MEM_stage_inst_dmem_ram_3361), .A2(MEM_stage_inst_dmem_n19750), .ZN(MEM_stage_inst_dmem_n19749) );
NAND2_X1 MEM_stage_inst_dmem_U19011 ( .A1(MEM_stage_inst_dmem_n19747), .A2(MEM_stage_inst_dmem_n19746), .ZN(MEM_stage_inst_dmem_n9565) );
NAND2_X1 MEM_stage_inst_dmem_U19010 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n19751), .ZN(MEM_stage_inst_dmem_n19746) );
NAND2_X1 MEM_stage_inst_dmem_U19009 ( .A1(MEM_stage_inst_dmem_ram_3362), .A2(MEM_stage_inst_dmem_n19750), .ZN(MEM_stage_inst_dmem_n19747) );
NAND2_X1 MEM_stage_inst_dmem_U19008 ( .A1(MEM_stage_inst_dmem_n19745), .A2(MEM_stage_inst_dmem_n19744), .ZN(MEM_stage_inst_dmem_n9566) );
NAND2_X1 MEM_stage_inst_dmem_U19007 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n19751), .ZN(MEM_stage_inst_dmem_n19744) );
NAND2_X1 MEM_stage_inst_dmem_U19006 ( .A1(MEM_stage_inst_dmem_ram_3363), .A2(MEM_stage_inst_dmem_n19750), .ZN(MEM_stage_inst_dmem_n19745) );
NAND2_X1 MEM_stage_inst_dmem_U19005 ( .A1(MEM_stage_inst_dmem_n19743), .A2(MEM_stage_inst_dmem_n19742), .ZN(MEM_stage_inst_dmem_n9567) );
NAND2_X1 MEM_stage_inst_dmem_U19004 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n19751), .ZN(MEM_stage_inst_dmem_n19742) );
NAND2_X1 MEM_stage_inst_dmem_U19003 ( .A1(MEM_stage_inst_dmem_ram_3364), .A2(MEM_stage_inst_dmem_n19750), .ZN(MEM_stage_inst_dmem_n19743) );
NAND2_X1 MEM_stage_inst_dmem_U19002 ( .A1(MEM_stage_inst_dmem_n19741), .A2(MEM_stage_inst_dmem_n19740), .ZN(MEM_stage_inst_dmem_n9568) );
NAND2_X1 MEM_stage_inst_dmem_U19001 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n19751), .ZN(MEM_stage_inst_dmem_n19740) );
NAND2_X1 MEM_stage_inst_dmem_U19000 ( .A1(MEM_stage_inst_dmem_ram_3365), .A2(MEM_stage_inst_dmem_n19750), .ZN(MEM_stage_inst_dmem_n19741) );
NAND2_X1 MEM_stage_inst_dmem_U18999 ( .A1(MEM_stage_inst_dmem_n19739), .A2(MEM_stage_inst_dmem_n19738), .ZN(MEM_stage_inst_dmem_n9569) );
NAND2_X1 MEM_stage_inst_dmem_U18998 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n19751), .ZN(MEM_stage_inst_dmem_n19738) );
NAND2_X1 MEM_stage_inst_dmem_U18997 ( .A1(MEM_stage_inst_dmem_ram_3366), .A2(MEM_stage_inst_dmem_n19750), .ZN(MEM_stage_inst_dmem_n19739) );
NAND2_X1 MEM_stage_inst_dmem_U18996 ( .A1(MEM_stage_inst_dmem_n19737), .A2(MEM_stage_inst_dmem_n19736), .ZN(MEM_stage_inst_dmem_n9570) );
NAND2_X1 MEM_stage_inst_dmem_U18995 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n19751), .ZN(MEM_stage_inst_dmem_n19736) );
NAND2_X1 MEM_stage_inst_dmem_U18994 ( .A1(MEM_stage_inst_dmem_ram_3367), .A2(MEM_stage_inst_dmem_n19750), .ZN(MEM_stage_inst_dmem_n19737) );
NAND2_X1 MEM_stage_inst_dmem_U18993 ( .A1(MEM_stage_inst_dmem_n19735), .A2(MEM_stage_inst_dmem_n19734), .ZN(MEM_stage_inst_dmem_n9571) );
NAND2_X1 MEM_stage_inst_dmem_U18992 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n19751), .ZN(MEM_stage_inst_dmem_n19734) );
NAND2_X1 MEM_stage_inst_dmem_U18991 ( .A1(MEM_stage_inst_dmem_ram_3368), .A2(MEM_stage_inst_dmem_n19750), .ZN(MEM_stage_inst_dmem_n19735) );
NAND2_X1 MEM_stage_inst_dmem_U18990 ( .A1(MEM_stage_inst_dmem_n19733), .A2(MEM_stage_inst_dmem_n19732), .ZN(MEM_stage_inst_dmem_n9572) );
NAND2_X1 MEM_stage_inst_dmem_U18989 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n19751), .ZN(MEM_stage_inst_dmem_n19732) );
NAND2_X1 MEM_stage_inst_dmem_U18988 ( .A1(MEM_stage_inst_dmem_ram_3369), .A2(MEM_stage_inst_dmem_n19750), .ZN(MEM_stage_inst_dmem_n19733) );
NAND2_X1 MEM_stage_inst_dmem_U18987 ( .A1(MEM_stage_inst_dmem_n19731), .A2(MEM_stage_inst_dmem_n19730), .ZN(MEM_stage_inst_dmem_n9573) );
NAND2_X1 MEM_stage_inst_dmem_U18986 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n19751), .ZN(MEM_stage_inst_dmem_n19730) );
NAND2_X1 MEM_stage_inst_dmem_U18985 ( .A1(MEM_stage_inst_dmem_ram_3370), .A2(MEM_stage_inst_dmem_n19750), .ZN(MEM_stage_inst_dmem_n19731) );
NAND2_X1 MEM_stage_inst_dmem_U18984 ( .A1(MEM_stage_inst_dmem_n19729), .A2(MEM_stage_inst_dmem_n19728), .ZN(MEM_stage_inst_dmem_n9574) );
NAND2_X1 MEM_stage_inst_dmem_U18983 ( .A1(MEM_stage_inst_dmem_n18004), .A2(MEM_stage_inst_dmem_n19751), .ZN(MEM_stage_inst_dmem_n19728) );
NAND2_X1 MEM_stage_inst_dmem_U18982 ( .A1(MEM_stage_inst_dmem_ram_3371), .A2(MEM_stage_inst_dmem_n19750), .ZN(MEM_stage_inst_dmem_n19729) );
NAND2_X1 MEM_stage_inst_dmem_U18981 ( .A1(MEM_stage_inst_dmem_n19727), .A2(MEM_stage_inst_dmem_n19726), .ZN(MEM_stage_inst_dmem_n9575) );
NAND2_X1 MEM_stage_inst_dmem_U18980 ( .A1(MEM_stage_inst_dmem_n21474), .A2(MEM_stage_inst_dmem_n19751), .ZN(MEM_stage_inst_dmem_n19726) );
NAND2_X1 MEM_stage_inst_dmem_U18979 ( .A1(MEM_stage_inst_dmem_ram_3372), .A2(MEM_stage_inst_dmem_n19750), .ZN(MEM_stage_inst_dmem_n19727) );
NAND2_X1 MEM_stage_inst_dmem_U18978 ( .A1(MEM_stage_inst_dmem_n19725), .A2(MEM_stage_inst_dmem_n19724), .ZN(MEM_stage_inst_dmem_n9576) );
NAND2_X1 MEM_stage_inst_dmem_U18977 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n19751), .ZN(MEM_stage_inst_dmem_n19724) );
NAND2_X1 MEM_stage_inst_dmem_U18976 ( .A1(MEM_stage_inst_dmem_ram_3373), .A2(MEM_stage_inst_dmem_n19750), .ZN(MEM_stage_inst_dmem_n19725) );
NAND2_X1 MEM_stage_inst_dmem_U18975 ( .A1(MEM_stage_inst_dmem_n19723), .A2(MEM_stage_inst_dmem_n19722), .ZN(MEM_stage_inst_dmem_n9577) );
NAND2_X1 MEM_stage_inst_dmem_U18974 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n19751), .ZN(MEM_stage_inst_dmem_n19722) );
NAND2_X1 MEM_stage_inst_dmem_U18973 ( .A1(MEM_stage_inst_dmem_ram_3374), .A2(MEM_stage_inst_dmem_n19750), .ZN(MEM_stage_inst_dmem_n19723) );
NAND2_X1 MEM_stage_inst_dmem_U18972 ( .A1(MEM_stage_inst_dmem_n19721), .A2(MEM_stage_inst_dmem_n19720), .ZN(MEM_stage_inst_dmem_n9578) );
NAND2_X1 MEM_stage_inst_dmem_U18971 ( .A1(MEM_stage_inst_dmem_n16343), .A2(MEM_stage_inst_dmem_n19751), .ZN(MEM_stage_inst_dmem_n19720) );
INV_X1 MEM_stage_inst_dmem_U18970 ( .A(MEM_stage_inst_dmem_n19750), .ZN(MEM_stage_inst_dmem_n19751) );
NAND2_X1 MEM_stage_inst_dmem_U18969 ( .A1(MEM_stage_inst_dmem_ram_3375), .A2(MEM_stage_inst_dmem_n19750), .ZN(MEM_stage_inst_dmem_n19721) );
NAND2_X1 MEM_stage_inst_dmem_U18968 ( .A1(MEM_stage_inst_dmem_n21394), .A2(MEM_stage_inst_dmem_n19788), .ZN(MEM_stage_inst_dmem_n19750) );
NAND2_X1 MEM_stage_inst_dmem_U18967 ( .A1(MEM_stage_inst_dmem_n19719), .A2(MEM_stage_inst_dmem_n19718), .ZN(MEM_stage_inst_dmem_n9579) );
NAND2_X1 MEM_stage_inst_dmem_U18966 ( .A1(MEM_stage_inst_dmem_n20551), .A2(MEM_stage_inst_dmem_n19717), .ZN(MEM_stage_inst_dmem_n19718) );
NAND2_X1 MEM_stage_inst_dmem_U18965 ( .A1(MEM_stage_inst_dmem_ram_3376), .A2(MEM_stage_inst_dmem_n19716), .ZN(MEM_stage_inst_dmem_n19719) );
NAND2_X1 MEM_stage_inst_dmem_U18964 ( .A1(MEM_stage_inst_dmem_n19715), .A2(MEM_stage_inst_dmem_n19714), .ZN(MEM_stage_inst_dmem_n9580) );
NAND2_X1 MEM_stage_inst_dmem_U18963 ( .A1(MEM_stage_inst_dmem_n20547), .A2(MEM_stage_inst_dmem_n19717), .ZN(MEM_stage_inst_dmem_n19714) );
NAND2_X1 MEM_stage_inst_dmem_U18962 ( .A1(MEM_stage_inst_dmem_ram_3377), .A2(MEM_stage_inst_dmem_n19716), .ZN(MEM_stage_inst_dmem_n19715) );
NAND2_X1 MEM_stage_inst_dmem_U18961 ( .A1(MEM_stage_inst_dmem_n19713), .A2(MEM_stage_inst_dmem_n19712), .ZN(MEM_stage_inst_dmem_n9581) );
NAND2_X1 MEM_stage_inst_dmem_U18960 ( .A1(MEM_stage_inst_dmem_n20544), .A2(MEM_stage_inst_dmem_n19717), .ZN(MEM_stage_inst_dmem_n19712) );
NAND2_X1 MEM_stage_inst_dmem_U18959 ( .A1(MEM_stage_inst_dmem_ram_3378), .A2(MEM_stage_inst_dmem_n19716), .ZN(MEM_stage_inst_dmem_n19713) );
NAND2_X1 MEM_stage_inst_dmem_U18958 ( .A1(MEM_stage_inst_dmem_n19711), .A2(MEM_stage_inst_dmem_n19710), .ZN(MEM_stage_inst_dmem_n9582) );
NAND2_X1 MEM_stage_inst_dmem_U18957 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n19717), .ZN(MEM_stage_inst_dmem_n19710) );
NAND2_X1 MEM_stage_inst_dmem_U18956 ( .A1(MEM_stage_inst_dmem_ram_3379), .A2(MEM_stage_inst_dmem_n19716), .ZN(MEM_stage_inst_dmem_n19711) );
NAND2_X1 MEM_stage_inst_dmem_U18955 ( .A1(MEM_stage_inst_dmem_n19709), .A2(MEM_stage_inst_dmem_n19708), .ZN(MEM_stage_inst_dmem_n9583) );
NAND2_X1 MEM_stage_inst_dmem_U18954 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n19717), .ZN(MEM_stage_inst_dmem_n19708) );
NAND2_X1 MEM_stage_inst_dmem_U18953 ( .A1(MEM_stage_inst_dmem_ram_3380), .A2(MEM_stage_inst_dmem_n19716), .ZN(MEM_stage_inst_dmem_n19709) );
NAND2_X1 MEM_stage_inst_dmem_U18952 ( .A1(MEM_stage_inst_dmem_n19707), .A2(MEM_stage_inst_dmem_n19706), .ZN(MEM_stage_inst_dmem_n9584) );
NAND2_X1 MEM_stage_inst_dmem_U18951 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n19717), .ZN(MEM_stage_inst_dmem_n19706) );
NAND2_X1 MEM_stage_inst_dmem_U18950 ( .A1(MEM_stage_inst_dmem_ram_3381), .A2(MEM_stage_inst_dmem_n19716), .ZN(MEM_stage_inst_dmem_n19707) );
NAND2_X1 MEM_stage_inst_dmem_U18949 ( .A1(MEM_stage_inst_dmem_n19705), .A2(MEM_stage_inst_dmem_n19704), .ZN(MEM_stage_inst_dmem_n9585) );
NAND2_X1 MEM_stage_inst_dmem_U18948 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n19717), .ZN(MEM_stage_inst_dmem_n19704) );
NAND2_X1 MEM_stage_inst_dmem_U18947 ( .A1(MEM_stage_inst_dmem_ram_3382), .A2(MEM_stage_inst_dmem_n19716), .ZN(MEM_stage_inst_dmem_n19705) );
NAND2_X1 MEM_stage_inst_dmem_U18946 ( .A1(MEM_stage_inst_dmem_n19703), .A2(MEM_stage_inst_dmem_n19702), .ZN(MEM_stage_inst_dmem_n9586) );
NAND2_X1 MEM_stage_inst_dmem_U18945 ( .A1(MEM_stage_inst_dmem_n20530), .A2(MEM_stage_inst_dmem_n19717), .ZN(MEM_stage_inst_dmem_n19702) );
NAND2_X1 MEM_stage_inst_dmem_U18944 ( .A1(MEM_stage_inst_dmem_ram_3383), .A2(MEM_stage_inst_dmem_n19716), .ZN(MEM_stage_inst_dmem_n19703) );
NAND2_X1 MEM_stage_inst_dmem_U18943 ( .A1(MEM_stage_inst_dmem_n19701), .A2(MEM_stage_inst_dmem_n19700), .ZN(MEM_stage_inst_dmem_n9587) );
NAND2_X1 MEM_stage_inst_dmem_U18942 ( .A1(MEM_stage_inst_dmem_n20527), .A2(MEM_stage_inst_dmem_n19717), .ZN(MEM_stage_inst_dmem_n19700) );
NAND2_X1 MEM_stage_inst_dmem_U18941 ( .A1(MEM_stage_inst_dmem_ram_3384), .A2(MEM_stage_inst_dmem_n19716), .ZN(MEM_stage_inst_dmem_n19701) );
NAND2_X1 MEM_stage_inst_dmem_U18940 ( .A1(MEM_stage_inst_dmem_n19699), .A2(MEM_stage_inst_dmem_n19698), .ZN(MEM_stage_inst_dmem_n9588) );
NAND2_X1 MEM_stage_inst_dmem_U18939 ( .A1(MEM_stage_inst_dmem_n20524), .A2(MEM_stage_inst_dmem_n19717), .ZN(MEM_stage_inst_dmem_n19698) );
NAND2_X1 MEM_stage_inst_dmem_U18938 ( .A1(MEM_stage_inst_dmem_ram_3385), .A2(MEM_stage_inst_dmem_n19716), .ZN(MEM_stage_inst_dmem_n19699) );
NAND2_X1 MEM_stage_inst_dmem_U18937 ( .A1(MEM_stage_inst_dmem_n19697), .A2(MEM_stage_inst_dmem_n19696), .ZN(MEM_stage_inst_dmem_n9589) );
NAND2_X1 MEM_stage_inst_dmem_U18936 ( .A1(MEM_stage_inst_dmem_n20521), .A2(MEM_stage_inst_dmem_n19717), .ZN(MEM_stage_inst_dmem_n19696) );
NAND2_X1 MEM_stage_inst_dmem_U18935 ( .A1(MEM_stage_inst_dmem_ram_3386), .A2(MEM_stage_inst_dmem_n19716), .ZN(MEM_stage_inst_dmem_n19697) );
NAND2_X1 MEM_stage_inst_dmem_U18934 ( .A1(MEM_stage_inst_dmem_n19695), .A2(MEM_stage_inst_dmem_n19694), .ZN(MEM_stage_inst_dmem_n9590) );
NAND2_X1 MEM_stage_inst_dmem_U18933 ( .A1(MEM_stage_inst_dmem_n20518), .A2(MEM_stage_inst_dmem_n19717), .ZN(MEM_stage_inst_dmem_n19694) );
NAND2_X1 MEM_stage_inst_dmem_U18932 ( .A1(MEM_stage_inst_dmem_ram_3387), .A2(MEM_stage_inst_dmem_n19716), .ZN(MEM_stage_inst_dmem_n19695) );
NAND2_X1 MEM_stage_inst_dmem_U18931 ( .A1(MEM_stage_inst_dmem_n19693), .A2(MEM_stage_inst_dmem_n19692), .ZN(MEM_stage_inst_dmem_n9591) );
NAND2_X1 MEM_stage_inst_dmem_U18930 ( .A1(MEM_stage_inst_dmem_n20515), .A2(MEM_stage_inst_dmem_n19717), .ZN(MEM_stage_inst_dmem_n19692) );
NAND2_X1 MEM_stage_inst_dmem_U18929 ( .A1(MEM_stage_inst_dmem_ram_3388), .A2(MEM_stage_inst_dmem_n19716), .ZN(MEM_stage_inst_dmem_n19693) );
NAND2_X1 MEM_stage_inst_dmem_U18928 ( .A1(MEM_stage_inst_dmem_n19691), .A2(MEM_stage_inst_dmem_n19690), .ZN(MEM_stage_inst_dmem_n9592) );
NAND2_X1 MEM_stage_inst_dmem_U18927 ( .A1(MEM_stage_inst_dmem_n20512), .A2(MEM_stage_inst_dmem_n19717), .ZN(MEM_stage_inst_dmem_n19690) );
NAND2_X1 MEM_stage_inst_dmem_U18926 ( .A1(MEM_stage_inst_dmem_ram_3389), .A2(MEM_stage_inst_dmem_n19716), .ZN(MEM_stage_inst_dmem_n19691) );
NAND2_X1 MEM_stage_inst_dmem_U18925 ( .A1(MEM_stage_inst_dmem_n19689), .A2(MEM_stage_inst_dmem_n19688), .ZN(MEM_stage_inst_dmem_n9593) );
NAND2_X1 MEM_stage_inst_dmem_U18924 ( .A1(MEM_stage_inst_dmem_n20509), .A2(MEM_stage_inst_dmem_n19717), .ZN(MEM_stage_inst_dmem_n19688) );
NAND2_X1 MEM_stage_inst_dmem_U18923 ( .A1(MEM_stage_inst_dmem_ram_3390), .A2(MEM_stage_inst_dmem_n19716), .ZN(MEM_stage_inst_dmem_n19689) );
NAND2_X1 MEM_stage_inst_dmem_U18922 ( .A1(MEM_stage_inst_dmem_n19687), .A2(MEM_stage_inst_dmem_n19686), .ZN(MEM_stage_inst_dmem_n9594) );
NAND2_X1 MEM_stage_inst_dmem_U18921 ( .A1(MEM_stage_inst_dmem_n20506), .A2(MEM_stage_inst_dmem_n19717), .ZN(MEM_stage_inst_dmem_n19686) );
INV_X1 MEM_stage_inst_dmem_U18920 ( .A(MEM_stage_inst_dmem_n19716), .ZN(MEM_stage_inst_dmem_n19717) );
NAND2_X1 MEM_stage_inst_dmem_U18919 ( .A1(MEM_stage_inst_dmem_ram_3391), .A2(MEM_stage_inst_dmem_n19716), .ZN(MEM_stage_inst_dmem_n19687) );
NAND2_X1 MEM_stage_inst_dmem_U18918 ( .A1(MEM_stage_inst_dmem_n21359), .A2(MEM_stage_inst_dmem_n19788), .ZN(MEM_stage_inst_dmem_n19716) );
NAND2_X1 MEM_stage_inst_dmem_U18917 ( .A1(MEM_stage_inst_dmem_n19685), .A2(MEM_stage_inst_dmem_n19684), .ZN(MEM_stage_inst_dmem_n9595) );
NAND2_X1 MEM_stage_inst_dmem_U18916 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n19683), .ZN(MEM_stage_inst_dmem_n19684) );
NAND2_X1 MEM_stage_inst_dmem_U18915 ( .A1(MEM_stage_inst_dmem_ram_3392), .A2(MEM_stage_inst_dmem_n19682), .ZN(MEM_stage_inst_dmem_n19685) );
NAND2_X1 MEM_stage_inst_dmem_U18914 ( .A1(MEM_stage_inst_dmem_n19681), .A2(MEM_stage_inst_dmem_n19680), .ZN(MEM_stage_inst_dmem_n9596) );
NAND2_X1 MEM_stage_inst_dmem_U18913 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n19683), .ZN(MEM_stage_inst_dmem_n19680) );
NAND2_X1 MEM_stage_inst_dmem_U18912 ( .A1(MEM_stage_inst_dmem_ram_3393), .A2(MEM_stage_inst_dmem_n19682), .ZN(MEM_stage_inst_dmem_n19681) );
NAND2_X1 MEM_stage_inst_dmem_U18911 ( .A1(MEM_stage_inst_dmem_n19679), .A2(MEM_stage_inst_dmem_n19678), .ZN(MEM_stage_inst_dmem_n9597) );
NAND2_X1 MEM_stage_inst_dmem_U18910 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n19683), .ZN(MEM_stage_inst_dmem_n19678) );
NAND2_X1 MEM_stage_inst_dmem_U18909 ( .A1(MEM_stage_inst_dmem_ram_3394), .A2(MEM_stage_inst_dmem_n19682), .ZN(MEM_stage_inst_dmem_n19679) );
NAND2_X1 MEM_stage_inst_dmem_U18908 ( .A1(MEM_stage_inst_dmem_n19677), .A2(MEM_stage_inst_dmem_n19676), .ZN(MEM_stage_inst_dmem_n9598) );
NAND2_X1 MEM_stage_inst_dmem_U18907 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n19683), .ZN(MEM_stage_inst_dmem_n19676) );
NAND2_X1 MEM_stage_inst_dmem_U18906 ( .A1(MEM_stage_inst_dmem_ram_3395), .A2(MEM_stage_inst_dmem_n19682), .ZN(MEM_stage_inst_dmem_n19677) );
NAND2_X1 MEM_stage_inst_dmem_U18905 ( .A1(MEM_stage_inst_dmem_n19675), .A2(MEM_stage_inst_dmem_n19674), .ZN(MEM_stage_inst_dmem_n9599) );
NAND2_X1 MEM_stage_inst_dmem_U18904 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n19683), .ZN(MEM_stage_inst_dmem_n19674) );
NAND2_X1 MEM_stage_inst_dmem_U18903 ( .A1(MEM_stage_inst_dmem_ram_3396), .A2(MEM_stage_inst_dmem_n19682), .ZN(MEM_stage_inst_dmem_n19675) );
NAND2_X1 MEM_stage_inst_dmem_U18902 ( .A1(MEM_stage_inst_dmem_n19673), .A2(MEM_stage_inst_dmem_n19672), .ZN(MEM_stage_inst_dmem_n9600) );
NAND2_X1 MEM_stage_inst_dmem_U18901 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n19683), .ZN(MEM_stage_inst_dmem_n19672) );
NAND2_X1 MEM_stage_inst_dmem_U18900 ( .A1(MEM_stage_inst_dmem_ram_3397), .A2(MEM_stage_inst_dmem_n19682), .ZN(MEM_stage_inst_dmem_n19673) );
NAND2_X1 MEM_stage_inst_dmem_U18899 ( .A1(MEM_stage_inst_dmem_n19671), .A2(MEM_stage_inst_dmem_n19670), .ZN(MEM_stage_inst_dmem_n9601) );
NAND2_X1 MEM_stage_inst_dmem_U18898 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n19683), .ZN(MEM_stage_inst_dmem_n19670) );
NAND2_X1 MEM_stage_inst_dmem_U18897 ( .A1(MEM_stage_inst_dmem_ram_3398), .A2(MEM_stage_inst_dmem_n19682), .ZN(MEM_stage_inst_dmem_n19671) );
NAND2_X1 MEM_stage_inst_dmem_U18896 ( .A1(MEM_stage_inst_dmem_n19669), .A2(MEM_stage_inst_dmem_n19668), .ZN(MEM_stage_inst_dmem_n9602) );
NAND2_X1 MEM_stage_inst_dmem_U18895 ( .A1(MEM_stage_inst_dmem_n20530), .A2(MEM_stage_inst_dmem_n19683), .ZN(MEM_stage_inst_dmem_n19668) );
NAND2_X1 MEM_stage_inst_dmem_U18894 ( .A1(MEM_stage_inst_dmem_ram_3399), .A2(MEM_stage_inst_dmem_n19682), .ZN(MEM_stage_inst_dmem_n19669) );
NAND2_X1 MEM_stage_inst_dmem_U18893 ( .A1(MEM_stage_inst_dmem_n19667), .A2(MEM_stage_inst_dmem_n19666), .ZN(MEM_stage_inst_dmem_n9603) );
NAND2_X1 MEM_stage_inst_dmem_U18892 ( .A1(EX_pipeline_reg_out_13), .A2(MEM_stage_inst_dmem_n19683), .ZN(MEM_stage_inst_dmem_n19666) );
NAND2_X1 MEM_stage_inst_dmem_U18891 ( .A1(MEM_stage_inst_dmem_ram_3400), .A2(MEM_stage_inst_dmem_n19682), .ZN(MEM_stage_inst_dmem_n19667) );
NAND2_X1 MEM_stage_inst_dmem_U18890 ( .A1(MEM_stage_inst_dmem_n19665), .A2(MEM_stage_inst_dmem_n19664), .ZN(MEM_stage_inst_dmem_n9604) );
NAND2_X1 MEM_stage_inst_dmem_U18889 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n19683), .ZN(MEM_stage_inst_dmem_n19664) );
NAND2_X1 MEM_stage_inst_dmem_U18888 ( .A1(MEM_stage_inst_dmem_ram_3401), .A2(MEM_stage_inst_dmem_n19682), .ZN(MEM_stage_inst_dmem_n19665) );
NAND2_X1 MEM_stage_inst_dmem_U18887 ( .A1(MEM_stage_inst_dmem_n19663), .A2(MEM_stage_inst_dmem_n19662), .ZN(MEM_stage_inst_dmem_n9605) );
NAND2_X1 MEM_stage_inst_dmem_U18886 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n19683), .ZN(MEM_stage_inst_dmem_n19662) );
NAND2_X1 MEM_stage_inst_dmem_U18885 ( .A1(MEM_stage_inst_dmem_ram_3402), .A2(MEM_stage_inst_dmem_n19682), .ZN(MEM_stage_inst_dmem_n19663) );
NAND2_X1 MEM_stage_inst_dmem_U18884 ( .A1(MEM_stage_inst_dmem_n19661), .A2(MEM_stage_inst_dmem_n19660), .ZN(MEM_stage_inst_dmem_n9606) );
NAND2_X1 MEM_stage_inst_dmem_U18883 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n19683), .ZN(MEM_stage_inst_dmem_n19660) );
NAND2_X1 MEM_stage_inst_dmem_U18882 ( .A1(MEM_stage_inst_dmem_ram_3403), .A2(MEM_stage_inst_dmem_n19682), .ZN(MEM_stage_inst_dmem_n19661) );
NAND2_X1 MEM_stage_inst_dmem_U18881 ( .A1(MEM_stage_inst_dmem_n19659), .A2(MEM_stage_inst_dmem_n19658), .ZN(MEM_stage_inst_dmem_n9607) );
NAND2_X1 MEM_stage_inst_dmem_U18880 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n19683), .ZN(MEM_stage_inst_dmem_n19658) );
NAND2_X1 MEM_stage_inst_dmem_U18879 ( .A1(MEM_stage_inst_dmem_ram_3404), .A2(MEM_stage_inst_dmem_n19682), .ZN(MEM_stage_inst_dmem_n19659) );
NAND2_X1 MEM_stage_inst_dmem_U18878 ( .A1(MEM_stage_inst_dmem_n19657), .A2(MEM_stage_inst_dmem_n19656), .ZN(MEM_stage_inst_dmem_n9608) );
NAND2_X1 MEM_stage_inst_dmem_U18877 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n19683), .ZN(MEM_stage_inst_dmem_n19656) );
NAND2_X1 MEM_stage_inst_dmem_U18876 ( .A1(MEM_stage_inst_dmem_ram_3405), .A2(MEM_stage_inst_dmem_n19682), .ZN(MEM_stage_inst_dmem_n19657) );
NAND2_X1 MEM_stage_inst_dmem_U18875 ( .A1(MEM_stage_inst_dmem_n19655), .A2(MEM_stage_inst_dmem_n19654), .ZN(MEM_stage_inst_dmem_n9609) );
NAND2_X1 MEM_stage_inst_dmem_U18874 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n19683), .ZN(MEM_stage_inst_dmem_n19654) );
NAND2_X1 MEM_stage_inst_dmem_U18873 ( .A1(MEM_stage_inst_dmem_ram_3406), .A2(MEM_stage_inst_dmem_n19682), .ZN(MEM_stage_inst_dmem_n19655) );
NAND2_X1 MEM_stage_inst_dmem_U18872 ( .A1(MEM_stage_inst_dmem_n19653), .A2(MEM_stage_inst_dmem_n19652), .ZN(MEM_stage_inst_dmem_n9610) );
NAND2_X1 MEM_stage_inst_dmem_U18871 ( .A1(MEM_stage_inst_dmem_n16343), .A2(MEM_stage_inst_dmem_n19683), .ZN(MEM_stage_inst_dmem_n19652) );
INV_X1 MEM_stage_inst_dmem_U18870 ( .A(MEM_stage_inst_dmem_n19682), .ZN(MEM_stage_inst_dmem_n19683) );
NAND2_X1 MEM_stage_inst_dmem_U18869 ( .A1(MEM_stage_inst_dmem_ram_3407), .A2(MEM_stage_inst_dmem_n19682), .ZN(MEM_stage_inst_dmem_n19653) );
NAND2_X1 MEM_stage_inst_dmem_U18868 ( .A1(MEM_stage_inst_dmem_n21319), .A2(MEM_stage_inst_dmem_n19788), .ZN(MEM_stage_inst_dmem_n19682) );
NAND2_X1 MEM_stage_inst_dmem_U18867 ( .A1(MEM_stage_inst_dmem_n19651), .A2(MEM_stage_inst_dmem_n19650), .ZN(MEM_stage_inst_dmem_n9611) );
NAND2_X1 MEM_stage_inst_dmem_U18866 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n19649), .ZN(MEM_stage_inst_dmem_n19650) );
NAND2_X1 MEM_stage_inst_dmem_U18865 ( .A1(MEM_stage_inst_dmem_ram_3408), .A2(MEM_stage_inst_dmem_n19648), .ZN(MEM_stage_inst_dmem_n19651) );
NAND2_X1 MEM_stage_inst_dmem_U18864 ( .A1(MEM_stage_inst_dmem_n19647), .A2(MEM_stage_inst_dmem_n19646), .ZN(MEM_stage_inst_dmem_n9612) );
NAND2_X1 MEM_stage_inst_dmem_U18863 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n19649), .ZN(MEM_stage_inst_dmem_n19646) );
NAND2_X1 MEM_stage_inst_dmem_U18862 ( .A1(MEM_stage_inst_dmem_ram_3409), .A2(MEM_stage_inst_dmem_n19648), .ZN(MEM_stage_inst_dmem_n19647) );
NAND2_X1 MEM_stage_inst_dmem_U18861 ( .A1(MEM_stage_inst_dmem_n19645), .A2(MEM_stage_inst_dmem_n19644), .ZN(MEM_stage_inst_dmem_n9613) );
NAND2_X1 MEM_stage_inst_dmem_U18860 ( .A1(MEM_stage_inst_dmem_n18027), .A2(MEM_stage_inst_dmem_n19649), .ZN(MEM_stage_inst_dmem_n19644) );
NAND2_X1 MEM_stage_inst_dmem_U18859 ( .A1(MEM_stage_inst_dmem_ram_3410), .A2(MEM_stage_inst_dmem_n19648), .ZN(MEM_stage_inst_dmem_n19645) );
NAND2_X1 MEM_stage_inst_dmem_U18858 ( .A1(MEM_stage_inst_dmem_n19643), .A2(MEM_stage_inst_dmem_n19642), .ZN(MEM_stage_inst_dmem_n9614) );
NAND2_X1 MEM_stage_inst_dmem_U18857 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n19649), .ZN(MEM_stage_inst_dmem_n19642) );
NAND2_X1 MEM_stage_inst_dmem_U18856 ( .A1(MEM_stage_inst_dmem_ram_3411), .A2(MEM_stage_inst_dmem_n19648), .ZN(MEM_stage_inst_dmem_n19643) );
NAND2_X1 MEM_stage_inst_dmem_U18855 ( .A1(MEM_stage_inst_dmem_n19641), .A2(MEM_stage_inst_dmem_n19640), .ZN(MEM_stage_inst_dmem_n9615) );
NAND2_X1 MEM_stage_inst_dmem_U18854 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n19649), .ZN(MEM_stage_inst_dmem_n19640) );
NAND2_X1 MEM_stage_inst_dmem_U18853 ( .A1(MEM_stage_inst_dmem_ram_3412), .A2(MEM_stage_inst_dmem_n19648), .ZN(MEM_stage_inst_dmem_n19641) );
NAND2_X1 MEM_stage_inst_dmem_U18852 ( .A1(MEM_stage_inst_dmem_n19639), .A2(MEM_stage_inst_dmem_n19638), .ZN(MEM_stage_inst_dmem_n9616) );
NAND2_X1 MEM_stage_inst_dmem_U18851 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n19649), .ZN(MEM_stage_inst_dmem_n19638) );
NAND2_X1 MEM_stage_inst_dmem_U18850 ( .A1(MEM_stage_inst_dmem_ram_3413), .A2(MEM_stage_inst_dmem_n19648), .ZN(MEM_stage_inst_dmem_n19639) );
NAND2_X1 MEM_stage_inst_dmem_U18849 ( .A1(MEM_stage_inst_dmem_n19637), .A2(MEM_stage_inst_dmem_n19636), .ZN(MEM_stage_inst_dmem_n9617) );
NAND2_X1 MEM_stage_inst_dmem_U18848 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n19649), .ZN(MEM_stage_inst_dmem_n19636) );
NAND2_X1 MEM_stage_inst_dmem_U18847 ( .A1(MEM_stage_inst_dmem_ram_3414), .A2(MEM_stage_inst_dmem_n19648), .ZN(MEM_stage_inst_dmem_n19637) );
NAND2_X1 MEM_stage_inst_dmem_U18846 ( .A1(MEM_stage_inst_dmem_n19635), .A2(MEM_stage_inst_dmem_n19634), .ZN(MEM_stage_inst_dmem_n9618) );
NAND2_X1 MEM_stage_inst_dmem_U18845 ( .A1(MEM_stage_inst_dmem_n17), .A2(MEM_stage_inst_dmem_n19649), .ZN(MEM_stage_inst_dmem_n19634) );
NAND2_X1 MEM_stage_inst_dmem_U18844 ( .A1(MEM_stage_inst_dmem_ram_3415), .A2(MEM_stage_inst_dmem_n19648), .ZN(MEM_stage_inst_dmem_n19635) );
NAND2_X1 MEM_stage_inst_dmem_U18843 ( .A1(MEM_stage_inst_dmem_n19633), .A2(MEM_stage_inst_dmem_n19632), .ZN(MEM_stage_inst_dmem_n9619) );
NAND2_X1 MEM_stage_inst_dmem_U18842 ( .A1(MEM_stage_inst_dmem_n18013), .A2(MEM_stage_inst_dmem_n19649), .ZN(MEM_stage_inst_dmem_n19632) );
NAND2_X1 MEM_stage_inst_dmem_U18841 ( .A1(MEM_stage_inst_dmem_ram_3416), .A2(MEM_stage_inst_dmem_n19648), .ZN(MEM_stage_inst_dmem_n19633) );
NAND2_X1 MEM_stage_inst_dmem_U18840 ( .A1(MEM_stage_inst_dmem_n19631), .A2(MEM_stage_inst_dmem_n19630), .ZN(MEM_stage_inst_dmem_n9620) );
NAND2_X1 MEM_stage_inst_dmem_U18839 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n19649), .ZN(MEM_stage_inst_dmem_n19630) );
NAND2_X1 MEM_stage_inst_dmem_U18838 ( .A1(MEM_stage_inst_dmem_ram_3417), .A2(MEM_stage_inst_dmem_n19648), .ZN(MEM_stage_inst_dmem_n19631) );
NAND2_X1 MEM_stage_inst_dmem_U18837 ( .A1(MEM_stage_inst_dmem_n19629), .A2(MEM_stage_inst_dmem_n19628), .ZN(MEM_stage_inst_dmem_n9621) );
NAND2_X1 MEM_stage_inst_dmem_U18836 ( .A1(MEM_stage_inst_dmem_n18007), .A2(MEM_stage_inst_dmem_n19649), .ZN(MEM_stage_inst_dmem_n19628) );
NAND2_X1 MEM_stage_inst_dmem_U18835 ( .A1(MEM_stage_inst_dmem_ram_3418), .A2(MEM_stage_inst_dmem_n19648), .ZN(MEM_stage_inst_dmem_n19629) );
NAND2_X1 MEM_stage_inst_dmem_U18834 ( .A1(MEM_stage_inst_dmem_n19627), .A2(MEM_stage_inst_dmem_n19626), .ZN(MEM_stage_inst_dmem_n9622) );
NAND2_X1 MEM_stage_inst_dmem_U18833 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n19649), .ZN(MEM_stage_inst_dmem_n19626) );
NAND2_X1 MEM_stage_inst_dmem_U18832 ( .A1(MEM_stage_inst_dmem_ram_3419), .A2(MEM_stage_inst_dmem_n19648), .ZN(MEM_stage_inst_dmem_n19627) );
NAND2_X1 MEM_stage_inst_dmem_U18831 ( .A1(MEM_stage_inst_dmem_n19625), .A2(MEM_stage_inst_dmem_n19624), .ZN(MEM_stage_inst_dmem_n9623) );
NAND2_X1 MEM_stage_inst_dmem_U18830 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n19649), .ZN(MEM_stage_inst_dmem_n19624) );
NAND2_X1 MEM_stage_inst_dmem_U18829 ( .A1(MEM_stage_inst_dmem_ram_3420), .A2(MEM_stage_inst_dmem_n19648), .ZN(MEM_stage_inst_dmem_n19625) );
NAND2_X1 MEM_stage_inst_dmem_U18828 ( .A1(MEM_stage_inst_dmem_n19623), .A2(MEM_stage_inst_dmem_n19622), .ZN(MEM_stage_inst_dmem_n9624) );
NAND2_X1 MEM_stage_inst_dmem_U18827 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n19649), .ZN(MEM_stage_inst_dmem_n19622) );
NAND2_X1 MEM_stage_inst_dmem_U18826 ( .A1(MEM_stage_inst_dmem_ram_3421), .A2(MEM_stage_inst_dmem_n19648), .ZN(MEM_stage_inst_dmem_n19623) );
NAND2_X1 MEM_stage_inst_dmem_U18825 ( .A1(MEM_stage_inst_dmem_n19621), .A2(MEM_stage_inst_dmem_n19620), .ZN(MEM_stage_inst_dmem_n9625) );
NAND2_X1 MEM_stage_inst_dmem_U18824 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n19649), .ZN(MEM_stage_inst_dmem_n19620) );
NAND2_X1 MEM_stage_inst_dmem_U18823 ( .A1(MEM_stage_inst_dmem_ram_3422), .A2(MEM_stage_inst_dmem_n19648), .ZN(MEM_stage_inst_dmem_n19621) );
NAND2_X1 MEM_stage_inst_dmem_U18822 ( .A1(MEM_stage_inst_dmem_n19619), .A2(MEM_stage_inst_dmem_n19618), .ZN(MEM_stage_inst_dmem_n9626) );
NAND2_X1 MEM_stage_inst_dmem_U18821 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n19649), .ZN(MEM_stage_inst_dmem_n19618) );
INV_X1 MEM_stage_inst_dmem_U18820 ( .A(MEM_stage_inst_dmem_n19648), .ZN(MEM_stage_inst_dmem_n19649) );
NAND2_X1 MEM_stage_inst_dmem_U18819 ( .A1(MEM_stage_inst_dmem_ram_3423), .A2(MEM_stage_inst_dmem_n19648), .ZN(MEM_stage_inst_dmem_n19619) );
NAND2_X1 MEM_stage_inst_dmem_U18818 ( .A1(MEM_stage_inst_dmem_n21284), .A2(MEM_stage_inst_dmem_n19788), .ZN(MEM_stage_inst_dmem_n19648) );
NAND2_X1 MEM_stage_inst_dmem_U18817 ( .A1(MEM_stage_inst_dmem_n19617), .A2(MEM_stage_inst_dmem_n19616), .ZN(MEM_stage_inst_dmem_n9627) );
NAND2_X1 MEM_stage_inst_dmem_U18816 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n19615), .ZN(MEM_stage_inst_dmem_n19616) );
NAND2_X1 MEM_stage_inst_dmem_U18815 ( .A1(MEM_stage_inst_dmem_ram_3424), .A2(MEM_stage_inst_dmem_n19614), .ZN(MEM_stage_inst_dmem_n19617) );
NAND2_X1 MEM_stage_inst_dmem_U18814 ( .A1(MEM_stage_inst_dmem_n19613), .A2(MEM_stage_inst_dmem_n19612), .ZN(MEM_stage_inst_dmem_n9628) );
NAND2_X1 MEM_stage_inst_dmem_U18813 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n19615), .ZN(MEM_stage_inst_dmem_n19612) );
NAND2_X1 MEM_stage_inst_dmem_U18812 ( .A1(MEM_stage_inst_dmem_ram_3425), .A2(MEM_stage_inst_dmem_n19614), .ZN(MEM_stage_inst_dmem_n19613) );
NAND2_X1 MEM_stage_inst_dmem_U18811 ( .A1(MEM_stage_inst_dmem_n19611), .A2(MEM_stage_inst_dmem_n19610), .ZN(MEM_stage_inst_dmem_n9629) );
NAND2_X1 MEM_stage_inst_dmem_U18810 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n19615), .ZN(MEM_stage_inst_dmem_n19610) );
NAND2_X1 MEM_stage_inst_dmem_U18809 ( .A1(MEM_stage_inst_dmem_ram_3426), .A2(MEM_stage_inst_dmem_n19614), .ZN(MEM_stage_inst_dmem_n19611) );
NAND2_X1 MEM_stage_inst_dmem_U18808 ( .A1(MEM_stage_inst_dmem_n19609), .A2(MEM_stage_inst_dmem_n19608), .ZN(MEM_stage_inst_dmem_n9630) );
NAND2_X1 MEM_stage_inst_dmem_U18807 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n19615), .ZN(MEM_stage_inst_dmem_n19608) );
NAND2_X1 MEM_stage_inst_dmem_U18806 ( .A1(MEM_stage_inst_dmem_ram_3427), .A2(MEM_stage_inst_dmem_n19614), .ZN(MEM_stage_inst_dmem_n19609) );
NAND2_X1 MEM_stage_inst_dmem_U18805 ( .A1(MEM_stage_inst_dmem_n19607), .A2(MEM_stage_inst_dmem_n19606), .ZN(MEM_stage_inst_dmem_n9631) );
NAND2_X1 MEM_stage_inst_dmem_U18804 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n19615), .ZN(MEM_stage_inst_dmem_n19606) );
NAND2_X1 MEM_stage_inst_dmem_U18803 ( .A1(MEM_stage_inst_dmem_ram_3428), .A2(MEM_stage_inst_dmem_n19614), .ZN(MEM_stage_inst_dmem_n19607) );
NAND2_X1 MEM_stage_inst_dmem_U18802 ( .A1(MEM_stage_inst_dmem_n19605), .A2(MEM_stage_inst_dmem_n19604), .ZN(MEM_stage_inst_dmem_n9632) );
NAND2_X1 MEM_stage_inst_dmem_U18801 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n19615), .ZN(MEM_stage_inst_dmem_n19604) );
NAND2_X1 MEM_stage_inst_dmem_U18800 ( .A1(MEM_stage_inst_dmem_ram_3429), .A2(MEM_stage_inst_dmem_n19614), .ZN(MEM_stage_inst_dmem_n19605) );
NAND2_X1 MEM_stage_inst_dmem_U18799 ( .A1(MEM_stage_inst_dmem_n19603), .A2(MEM_stage_inst_dmem_n19602), .ZN(MEM_stage_inst_dmem_n9633) );
NAND2_X1 MEM_stage_inst_dmem_U18798 ( .A1(MEM_stage_inst_dmem_n14717), .A2(MEM_stage_inst_dmem_n19615), .ZN(MEM_stage_inst_dmem_n19602) );
NAND2_X1 MEM_stage_inst_dmem_U18797 ( .A1(MEM_stage_inst_dmem_ram_3430), .A2(MEM_stage_inst_dmem_n19614), .ZN(MEM_stage_inst_dmem_n19603) );
NAND2_X1 MEM_stage_inst_dmem_U18796 ( .A1(MEM_stage_inst_dmem_n19601), .A2(MEM_stage_inst_dmem_n19600), .ZN(MEM_stage_inst_dmem_n9634) );
NAND2_X1 MEM_stage_inst_dmem_U18795 ( .A1(MEM_stage_inst_dmem_n18875), .A2(MEM_stage_inst_dmem_n19615), .ZN(MEM_stage_inst_dmem_n19600) );
NAND2_X1 MEM_stage_inst_dmem_U18794 ( .A1(MEM_stage_inst_dmem_ram_3431), .A2(MEM_stage_inst_dmem_n19614), .ZN(MEM_stage_inst_dmem_n19601) );
NAND2_X1 MEM_stage_inst_dmem_U18793 ( .A1(MEM_stage_inst_dmem_n19599), .A2(MEM_stage_inst_dmem_n19598), .ZN(MEM_stage_inst_dmem_n9635) );
NAND2_X1 MEM_stage_inst_dmem_U18792 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n19615), .ZN(MEM_stage_inst_dmem_n19598) );
NAND2_X1 MEM_stage_inst_dmem_U18791 ( .A1(MEM_stage_inst_dmem_ram_3432), .A2(MEM_stage_inst_dmem_n19614), .ZN(MEM_stage_inst_dmem_n19599) );
NAND2_X1 MEM_stage_inst_dmem_U18790 ( .A1(MEM_stage_inst_dmem_n19597), .A2(MEM_stage_inst_dmem_n19596), .ZN(MEM_stage_inst_dmem_n9636) );
NAND2_X1 MEM_stage_inst_dmem_U18789 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n19615), .ZN(MEM_stage_inst_dmem_n19596) );
NAND2_X1 MEM_stage_inst_dmem_U18788 ( .A1(MEM_stage_inst_dmem_ram_3433), .A2(MEM_stage_inst_dmem_n19614), .ZN(MEM_stage_inst_dmem_n19597) );
NAND2_X1 MEM_stage_inst_dmem_U18787 ( .A1(MEM_stage_inst_dmem_n19595), .A2(MEM_stage_inst_dmem_n19594), .ZN(MEM_stage_inst_dmem_n9637) );
NAND2_X1 MEM_stage_inst_dmem_U18786 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n19615), .ZN(MEM_stage_inst_dmem_n19594) );
NAND2_X1 MEM_stage_inst_dmem_U18785 ( .A1(MEM_stage_inst_dmem_ram_3434), .A2(MEM_stage_inst_dmem_n19614), .ZN(MEM_stage_inst_dmem_n19595) );
NAND2_X1 MEM_stage_inst_dmem_U18784 ( .A1(MEM_stage_inst_dmem_n19593), .A2(MEM_stage_inst_dmem_n19592), .ZN(MEM_stage_inst_dmem_n9638) );
NAND2_X1 MEM_stage_inst_dmem_U18783 ( .A1(MEM_stage_inst_dmem_n18004), .A2(MEM_stage_inst_dmem_n19615), .ZN(MEM_stage_inst_dmem_n19592) );
NAND2_X1 MEM_stage_inst_dmem_U18782 ( .A1(MEM_stage_inst_dmem_ram_3435), .A2(MEM_stage_inst_dmem_n19614), .ZN(MEM_stage_inst_dmem_n19593) );
NAND2_X1 MEM_stage_inst_dmem_U18781 ( .A1(MEM_stage_inst_dmem_n19591), .A2(MEM_stage_inst_dmem_n19590), .ZN(MEM_stage_inst_dmem_n9639) );
NAND2_X1 MEM_stage_inst_dmem_U18780 ( .A1(MEM_stage_inst_dmem_n18001), .A2(MEM_stage_inst_dmem_n19615), .ZN(MEM_stage_inst_dmem_n19590) );
NAND2_X1 MEM_stage_inst_dmem_U18779 ( .A1(MEM_stage_inst_dmem_ram_3436), .A2(MEM_stage_inst_dmem_n19614), .ZN(MEM_stage_inst_dmem_n19591) );
NAND2_X1 MEM_stage_inst_dmem_U18778 ( .A1(MEM_stage_inst_dmem_n19589), .A2(MEM_stage_inst_dmem_n19588), .ZN(MEM_stage_inst_dmem_n9640) );
NAND2_X1 MEM_stage_inst_dmem_U18777 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n19615), .ZN(MEM_stage_inst_dmem_n19588) );
NAND2_X1 MEM_stage_inst_dmem_U18776 ( .A1(MEM_stage_inst_dmem_ram_3437), .A2(MEM_stage_inst_dmem_n19614), .ZN(MEM_stage_inst_dmem_n19589) );
NAND2_X1 MEM_stage_inst_dmem_U18775 ( .A1(MEM_stage_inst_dmem_n19587), .A2(MEM_stage_inst_dmem_n19586), .ZN(MEM_stage_inst_dmem_n9641) );
NAND2_X1 MEM_stage_inst_dmem_U18774 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n19615), .ZN(MEM_stage_inst_dmem_n19586) );
NAND2_X1 MEM_stage_inst_dmem_U18773 ( .A1(MEM_stage_inst_dmem_ram_3438), .A2(MEM_stage_inst_dmem_n19614), .ZN(MEM_stage_inst_dmem_n19587) );
NAND2_X1 MEM_stage_inst_dmem_U18772 ( .A1(MEM_stage_inst_dmem_n19585), .A2(MEM_stage_inst_dmem_n19584), .ZN(MEM_stage_inst_dmem_n9642) );
NAND2_X1 MEM_stage_inst_dmem_U18771 ( .A1(MEM_stage_inst_dmem_n15110), .A2(MEM_stage_inst_dmem_n19615), .ZN(MEM_stage_inst_dmem_n19584) );
INV_X1 MEM_stage_inst_dmem_U18770 ( .A(MEM_stage_inst_dmem_n19614), .ZN(MEM_stage_inst_dmem_n19615) );
NAND2_X1 MEM_stage_inst_dmem_U18769 ( .A1(MEM_stage_inst_dmem_ram_3439), .A2(MEM_stage_inst_dmem_n19614), .ZN(MEM_stage_inst_dmem_n19585) );
NAND2_X1 MEM_stage_inst_dmem_U18768 ( .A1(MEM_stage_inst_dmem_n21249), .A2(MEM_stage_inst_dmem_n19788), .ZN(MEM_stage_inst_dmem_n19614) );
NAND2_X1 MEM_stage_inst_dmem_U18767 ( .A1(MEM_stage_inst_dmem_n19583), .A2(MEM_stage_inst_dmem_n19582), .ZN(MEM_stage_inst_dmem_n9643) );
NAND2_X1 MEM_stage_inst_dmem_U18766 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n19581), .ZN(MEM_stage_inst_dmem_n19582) );
NAND2_X1 MEM_stage_inst_dmem_U18765 ( .A1(MEM_stage_inst_dmem_ram_3440), .A2(MEM_stage_inst_dmem_n19580), .ZN(MEM_stage_inst_dmem_n19583) );
NAND2_X1 MEM_stage_inst_dmem_U18764 ( .A1(MEM_stage_inst_dmem_n19579), .A2(MEM_stage_inst_dmem_n19578), .ZN(MEM_stage_inst_dmem_n9644) );
NAND2_X1 MEM_stage_inst_dmem_U18763 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n19581), .ZN(MEM_stage_inst_dmem_n19578) );
NAND2_X1 MEM_stage_inst_dmem_U18762 ( .A1(MEM_stage_inst_dmem_ram_3441), .A2(MEM_stage_inst_dmem_n19580), .ZN(MEM_stage_inst_dmem_n19579) );
NAND2_X1 MEM_stage_inst_dmem_U18761 ( .A1(MEM_stage_inst_dmem_n19577), .A2(MEM_stage_inst_dmem_n19576), .ZN(MEM_stage_inst_dmem_n9645) );
NAND2_X1 MEM_stage_inst_dmem_U18760 ( .A1(EX_pipeline_reg_out_7), .A2(MEM_stage_inst_dmem_n19581), .ZN(MEM_stage_inst_dmem_n19576) );
NAND2_X1 MEM_stage_inst_dmem_U18759 ( .A1(MEM_stage_inst_dmem_ram_3442), .A2(MEM_stage_inst_dmem_n19580), .ZN(MEM_stage_inst_dmem_n19577) );
NAND2_X1 MEM_stage_inst_dmem_U18758 ( .A1(MEM_stage_inst_dmem_n19575), .A2(MEM_stage_inst_dmem_n19574), .ZN(MEM_stage_inst_dmem_n9646) );
NAND2_X1 MEM_stage_inst_dmem_U18757 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n19581), .ZN(MEM_stage_inst_dmem_n19574) );
NAND2_X1 MEM_stage_inst_dmem_U18756 ( .A1(MEM_stage_inst_dmem_ram_3443), .A2(MEM_stage_inst_dmem_n19580), .ZN(MEM_stage_inst_dmem_n19575) );
NAND2_X1 MEM_stage_inst_dmem_U18755 ( .A1(MEM_stage_inst_dmem_n19573), .A2(MEM_stage_inst_dmem_n19572), .ZN(MEM_stage_inst_dmem_n9647) );
NAND2_X1 MEM_stage_inst_dmem_U18754 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n19581), .ZN(MEM_stage_inst_dmem_n19572) );
NAND2_X1 MEM_stage_inst_dmem_U18753 ( .A1(MEM_stage_inst_dmem_ram_3444), .A2(MEM_stage_inst_dmem_n19580), .ZN(MEM_stage_inst_dmem_n19573) );
NAND2_X1 MEM_stage_inst_dmem_U18752 ( .A1(MEM_stage_inst_dmem_n19571), .A2(MEM_stage_inst_dmem_n19570), .ZN(MEM_stage_inst_dmem_n9648) );
NAND2_X1 MEM_stage_inst_dmem_U18751 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n19581), .ZN(MEM_stage_inst_dmem_n19570) );
NAND2_X1 MEM_stage_inst_dmem_U18750 ( .A1(MEM_stage_inst_dmem_ram_3445), .A2(MEM_stage_inst_dmem_n19580), .ZN(MEM_stage_inst_dmem_n19571) );
NAND2_X1 MEM_stage_inst_dmem_U18749 ( .A1(MEM_stage_inst_dmem_n19569), .A2(MEM_stage_inst_dmem_n19568), .ZN(MEM_stage_inst_dmem_n9649) );
NAND2_X1 MEM_stage_inst_dmem_U18748 ( .A1(MEM_stage_inst_dmem_n14717), .A2(MEM_stage_inst_dmem_n19581), .ZN(MEM_stage_inst_dmem_n19568) );
NAND2_X1 MEM_stage_inst_dmem_U18747 ( .A1(MEM_stage_inst_dmem_ram_3446), .A2(MEM_stage_inst_dmem_n19580), .ZN(MEM_stage_inst_dmem_n19569) );
NAND2_X1 MEM_stage_inst_dmem_U18746 ( .A1(MEM_stage_inst_dmem_n19567), .A2(MEM_stage_inst_dmem_n19566), .ZN(MEM_stage_inst_dmem_n9650) );
NAND2_X1 MEM_stage_inst_dmem_U18745 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n19581), .ZN(MEM_stage_inst_dmem_n19566) );
NAND2_X1 MEM_stage_inst_dmem_U18744 ( .A1(MEM_stage_inst_dmem_ram_3447), .A2(MEM_stage_inst_dmem_n19580), .ZN(MEM_stage_inst_dmem_n19567) );
NAND2_X1 MEM_stage_inst_dmem_U18743 ( .A1(MEM_stage_inst_dmem_n19565), .A2(MEM_stage_inst_dmem_n19564), .ZN(MEM_stage_inst_dmem_n9651) );
NAND2_X1 MEM_stage_inst_dmem_U18742 ( .A1(MEM_stage_inst_dmem_n13051), .A2(MEM_stage_inst_dmem_n19581), .ZN(MEM_stage_inst_dmem_n19564) );
NAND2_X1 MEM_stage_inst_dmem_U18741 ( .A1(MEM_stage_inst_dmem_ram_3448), .A2(MEM_stage_inst_dmem_n19580), .ZN(MEM_stage_inst_dmem_n19565) );
NAND2_X1 MEM_stage_inst_dmem_U18740 ( .A1(MEM_stage_inst_dmem_n19563), .A2(MEM_stage_inst_dmem_n19562), .ZN(MEM_stage_inst_dmem_n9652) );
NAND2_X1 MEM_stage_inst_dmem_U18739 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n19581), .ZN(MEM_stage_inst_dmem_n19562) );
NAND2_X1 MEM_stage_inst_dmem_U18738 ( .A1(MEM_stage_inst_dmem_ram_3449), .A2(MEM_stage_inst_dmem_n19580), .ZN(MEM_stage_inst_dmem_n19563) );
NAND2_X1 MEM_stage_inst_dmem_U18737 ( .A1(MEM_stage_inst_dmem_n19561), .A2(MEM_stage_inst_dmem_n19560), .ZN(MEM_stage_inst_dmem_n9653) );
NAND2_X1 MEM_stage_inst_dmem_U18736 ( .A1(EX_pipeline_reg_out_15), .A2(MEM_stage_inst_dmem_n19581), .ZN(MEM_stage_inst_dmem_n19560) );
NAND2_X1 MEM_stage_inst_dmem_U18735 ( .A1(MEM_stage_inst_dmem_ram_3450), .A2(MEM_stage_inst_dmem_n19580), .ZN(MEM_stage_inst_dmem_n19561) );
NAND2_X1 MEM_stage_inst_dmem_U18734 ( .A1(MEM_stage_inst_dmem_n19559), .A2(MEM_stage_inst_dmem_n19558), .ZN(MEM_stage_inst_dmem_n9654) );
NAND2_X1 MEM_stage_inst_dmem_U18733 ( .A1(MEM_stage_inst_dmem_n20904), .A2(MEM_stage_inst_dmem_n19581), .ZN(MEM_stage_inst_dmem_n19558) );
NAND2_X1 MEM_stage_inst_dmem_U18732 ( .A1(MEM_stage_inst_dmem_ram_3451), .A2(MEM_stage_inst_dmem_n19580), .ZN(MEM_stage_inst_dmem_n19559) );
NAND2_X1 MEM_stage_inst_dmem_U18731 ( .A1(MEM_stage_inst_dmem_n19557), .A2(MEM_stage_inst_dmem_n19556), .ZN(MEM_stage_inst_dmem_n9655) );
NAND2_X1 MEM_stage_inst_dmem_U18730 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n19581), .ZN(MEM_stage_inst_dmem_n19556) );
NAND2_X1 MEM_stage_inst_dmem_U18729 ( .A1(MEM_stage_inst_dmem_ram_3452), .A2(MEM_stage_inst_dmem_n19580), .ZN(MEM_stage_inst_dmem_n19557) );
NAND2_X1 MEM_stage_inst_dmem_U18728 ( .A1(MEM_stage_inst_dmem_n19555), .A2(MEM_stage_inst_dmem_n19554), .ZN(MEM_stage_inst_dmem_n9656) );
NAND2_X1 MEM_stage_inst_dmem_U18727 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n19581), .ZN(MEM_stage_inst_dmem_n19554) );
NAND2_X1 MEM_stage_inst_dmem_U18726 ( .A1(MEM_stage_inst_dmem_ram_3453), .A2(MEM_stage_inst_dmem_n19580), .ZN(MEM_stage_inst_dmem_n19555) );
NAND2_X1 MEM_stage_inst_dmem_U18725 ( .A1(MEM_stage_inst_dmem_n19553), .A2(MEM_stage_inst_dmem_n19552), .ZN(MEM_stage_inst_dmem_n9657) );
NAND2_X1 MEM_stage_inst_dmem_U18724 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n19581), .ZN(MEM_stage_inst_dmem_n19552) );
NAND2_X1 MEM_stage_inst_dmem_U18723 ( .A1(MEM_stage_inst_dmem_ram_3454), .A2(MEM_stage_inst_dmem_n19580), .ZN(MEM_stage_inst_dmem_n19553) );
NAND2_X1 MEM_stage_inst_dmem_U18722 ( .A1(MEM_stage_inst_dmem_n19551), .A2(MEM_stage_inst_dmem_n19550), .ZN(MEM_stage_inst_dmem_n9658) );
NAND2_X1 MEM_stage_inst_dmem_U18721 ( .A1(EX_pipeline_reg_out_20), .A2(MEM_stage_inst_dmem_n19581), .ZN(MEM_stage_inst_dmem_n19550) );
NAND2_X1 MEM_stage_inst_dmem_U18720 ( .A1(MEM_stage_inst_dmem_ram_3455), .A2(MEM_stage_inst_dmem_n19580), .ZN(MEM_stage_inst_dmem_n19551) );
NAND2_X1 MEM_stage_inst_dmem_U18719 ( .A1(MEM_stage_inst_dmem_n21214), .A2(MEM_stage_inst_dmem_n19788), .ZN(MEM_stage_inst_dmem_n19580) );
NAND2_X1 MEM_stage_inst_dmem_U18718 ( .A1(MEM_stage_inst_dmem_n19549), .A2(MEM_stage_inst_dmem_n19548), .ZN(MEM_stage_inst_dmem_n9659) );
NAND2_X1 MEM_stage_inst_dmem_U18717 ( .A1(MEM_stage_inst_dmem_n20551), .A2(MEM_stage_inst_dmem_n19547), .ZN(MEM_stage_inst_dmem_n19548) );
NAND2_X1 MEM_stage_inst_dmem_U18716 ( .A1(MEM_stage_inst_dmem_ram_3456), .A2(MEM_stage_inst_dmem_n19546), .ZN(MEM_stage_inst_dmem_n19549) );
NAND2_X1 MEM_stage_inst_dmem_U18715 ( .A1(MEM_stage_inst_dmem_n19545), .A2(MEM_stage_inst_dmem_n19544), .ZN(MEM_stage_inst_dmem_n9660) );
NAND2_X1 MEM_stage_inst_dmem_U18714 ( .A1(MEM_stage_inst_dmem_n20547), .A2(MEM_stage_inst_dmem_n19547), .ZN(MEM_stage_inst_dmem_n19544) );
NAND2_X1 MEM_stage_inst_dmem_U18713 ( .A1(MEM_stage_inst_dmem_ram_3457), .A2(MEM_stage_inst_dmem_n19546), .ZN(MEM_stage_inst_dmem_n19545) );
NAND2_X1 MEM_stage_inst_dmem_U18712 ( .A1(MEM_stage_inst_dmem_n19543), .A2(MEM_stage_inst_dmem_n19542), .ZN(MEM_stage_inst_dmem_n9661) );
NAND2_X1 MEM_stage_inst_dmem_U18711 ( .A1(MEM_stage_inst_dmem_n20544), .A2(MEM_stage_inst_dmem_n19547), .ZN(MEM_stage_inst_dmem_n19542) );
NAND2_X1 MEM_stage_inst_dmem_U18710 ( .A1(MEM_stage_inst_dmem_ram_3458), .A2(MEM_stage_inst_dmem_n19546), .ZN(MEM_stage_inst_dmem_n19543) );
NAND2_X1 MEM_stage_inst_dmem_U18709 ( .A1(MEM_stage_inst_dmem_n19541), .A2(MEM_stage_inst_dmem_n19540), .ZN(MEM_stage_inst_dmem_n9662) );
NAND2_X1 MEM_stage_inst_dmem_U18708 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n19547), .ZN(MEM_stage_inst_dmem_n19540) );
NAND2_X1 MEM_stage_inst_dmem_U18707 ( .A1(MEM_stage_inst_dmem_ram_3459), .A2(MEM_stage_inst_dmem_n19546), .ZN(MEM_stage_inst_dmem_n19541) );
NAND2_X1 MEM_stage_inst_dmem_U18706 ( .A1(MEM_stage_inst_dmem_n19539), .A2(MEM_stage_inst_dmem_n19538), .ZN(MEM_stage_inst_dmem_n9663) );
NAND2_X1 MEM_stage_inst_dmem_U18705 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n19547), .ZN(MEM_stage_inst_dmem_n19538) );
NAND2_X1 MEM_stage_inst_dmem_U18704 ( .A1(MEM_stage_inst_dmem_ram_3460), .A2(MEM_stage_inst_dmem_n19546), .ZN(MEM_stage_inst_dmem_n19539) );
NAND2_X1 MEM_stage_inst_dmem_U18703 ( .A1(MEM_stage_inst_dmem_n19537), .A2(MEM_stage_inst_dmem_n19536), .ZN(MEM_stage_inst_dmem_n9664) );
NAND2_X1 MEM_stage_inst_dmem_U18702 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n19547), .ZN(MEM_stage_inst_dmem_n19536) );
NAND2_X1 MEM_stage_inst_dmem_U18701 ( .A1(MEM_stage_inst_dmem_ram_3461), .A2(MEM_stage_inst_dmem_n19546), .ZN(MEM_stage_inst_dmem_n19537) );
NAND2_X1 MEM_stage_inst_dmem_U18700 ( .A1(MEM_stage_inst_dmem_n19535), .A2(MEM_stage_inst_dmem_n19534), .ZN(MEM_stage_inst_dmem_n9665) );
NAND2_X1 MEM_stage_inst_dmem_U18699 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n19547), .ZN(MEM_stage_inst_dmem_n19534) );
NAND2_X1 MEM_stage_inst_dmem_U18698 ( .A1(MEM_stage_inst_dmem_ram_3462), .A2(MEM_stage_inst_dmem_n19546), .ZN(MEM_stage_inst_dmem_n19535) );
NAND2_X1 MEM_stage_inst_dmem_U18697 ( .A1(MEM_stage_inst_dmem_n19533), .A2(MEM_stage_inst_dmem_n19532), .ZN(MEM_stage_inst_dmem_n9666) );
NAND2_X1 MEM_stage_inst_dmem_U18696 ( .A1(MEM_stage_inst_dmem_n20530), .A2(MEM_stage_inst_dmem_n19547), .ZN(MEM_stage_inst_dmem_n19532) );
NAND2_X1 MEM_stage_inst_dmem_U18695 ( .A1(MEM_stage_inst_dmem_ram_3463), .A2(MEM_stage_inst_dmem_n19546), .ZN(MEM_stage_inst_dmem_n19533) );
NAND2_X1 MEM_stage_inst_dmem_U18694 ( .A1(MEM_stage_inst_dmem_n19531), .A2(MEM_stage_inst_dmem_n19530), .ZN(MEM_stage_inst_dmem_n9667) );
NAND2_X1 MEM_stage_inst_dmem_U18693 ( .A1(MEM_stage_inst_dmem_n20527), .A2(MEM_stage_inst_dmem_n19547), .ZN(MEM_stage_inst_dmem_n19530) );
NAND2_X1 MEM_stage_inst_dmem_U18692 ( .A1(MEM_stage_inst_dmem_ram_3464), .A2(MEM_stage_inst_dmem_n19546), .ZN(MEM_stage_inst_dmem_n19531) );
NAND2_X1 MEM_stage_inst_dmem_U18691 ( .A1(MEM_stage_inst_dmem_n19529), .A2(MEM_stage_inst_dmem_n19528), .ZN(MEM_stage_inst_dmem_n9668) );
NAND2_X1 MEM_stage_inst_dmem_U18690 ( .A1(MEM_stage_inst_dmem_n20524), .A2(MEM_stage_inst_dmem_n19547), .ZN(MEM_stage_inst_dmem_n19528) );
NAND2_X1 MEM_stage_inst_dmem_U18689 ( .A1(MEM_stage_inst_dmem_ram_3465), .A2(MEM_stage_inst_dmem_n19546), .ZN(MEM_stage_inst_dmem_n19529) );
NAND2_X1 MEM_stage_inst_dmem_U18688 ( .A1(MEM_stage_inst_dmem_n19527), .A2(MEM_stage_inst_dmem_n19526), .ZN(MEM_stage_inst_dmem_n9669) );
NAND2_X1 MEM_stage_inst_dmem_U18687 ( .A1(MEM_stage_inst_dmem_n20521), .A2(MEM_stage_inst_dmem_n19547), .ZN(MEM_stage_inst_dmem_n19526) );
NAND2_X1 MEM_stage_inst_dmem_U18686 ( .A1(MEM_stage_inst_dmem_ram_3466), .A2(MEM_stage_inst_dmem_n19546), .ZN(MEM_stage_inst_dmem_n19527) );
NAND2_X1 MEM_stage_inst_dmem_U18685 ( .A1(MEM_stage_inst_dmem_n19525), .A2(MEM_stage_inst_dmem_n19524), .ZN(MEM_stage_inst_dmem_n9670) );
NAND2_X1 MEM_stage_inst_dmem_U18684 ( .A1(MEM_stage_inst_dmem_n20518), .A2(MEM_stage_inst_dmem_n19547), .ZN(MEM_stage_inst_dmem_n19524) );
NAND2_X1 MEM_stage_inst_dmem_U18683 ( .A1(MEM_stage_inst_dmem_ram_3467), .A2(MEM_stage_inst_dmem_n19546), .ZN(MEM_stage_inst_dmem_n19525) );
NAND2_X1 MEM_stage_inst_dmem_U18682 ( .A1(MEM_stage_inst_dmem_n19523), .A2(MEM_stage_inst_dmem_n19522), .ZN(MEM_stage_inst_dmem_n9671) );
NAND2_X1 MEM_stage_inst_dmem_U18681 ( .A1(MEM_stage_inst_dmem_n20515), .A2(MEM_stage_inst_dmem_n19547), .ZN(MEM_stage_inst_dmem_n19522) );
NAND2_X1 MEM_stage_inst_dmem_U18680 ( .A1(MEM_stage_inst_dmem_ram_3468), .A2(MEM_stage_inst_dmem_n19546), .ZN(MEM_stage_inst_dmem_n19523) );
NAND2_X1 MEM_stage_inst_dmem_U18679 ( .A1(MEM_stage_inst_dmem_n19521), .A2(MEM_stage_inst_dmem_n19520), .ZN(MEM_stage_inst_dmem_n9672) );
NAND2_X1 MEM_stage_inst_dmem_U18678 ( .A1(MEM_stage_inst_dmem_n20512), .A2(MEM_stage_inst_dmem_n19547), .ZN(MEM_stage_inst_dmem_n19520) );
NAND2_X1 MEM_stage_inst_dmem_U18677 ( .A1(MEM_stage_inst_dmem_ram_3469), .A2(MEM_stage_inst_dmem_n19546), .ZN(MEM_stage_inst_dmem_n19521) );
NAND2_X1 MEM_stage_inst_dmem_U18676 ( .A1(MEM_stage_inst_dmem_n19519), .A2(MEM_stage_inst_dmem_n19518), .ZN(MEM_stage_inst_dmem_n9673) );
NAND2_X1 MEM_stage_inst_dmem_U18675 ( .A1(MEM_stage_inst_dmem_n20509), .A2(MEM_stage_inst_dmem_n19547), .ZN(MEM_stage_inst_dmem_n19518) );
NAND2_X1 MEM_stage_inst_dmem_U18674 ( .A1(MEM_stage_inst_dmem_ram_3470), .A2(MEM_stage_inst_dmem_n19546), .ZN(MEM_stage_inst_dmem_n19519) );
NAND2_X1 MEM_stage_inst_dmem_U18673 ( .A1(MEM_stage_inst_dmem_n19517), .A2(MEM_stage_inst_dmem_n19516), .ZN(MEM_stage_inst_dmem_n9674) );
NAND2_X1 MEM_stage_inst_dmem_U18672 ( .A1(MEM_stage_inst_dmem_n20506), .A2(MEM_stage_inst_dmem_n19547), .ZN(MEM_stage_inst_dmem_n19516) );
INV_X1 MEM_stage_inst_dmem_U18671 ( .A(MEM_stage_inst_dmem_n19546), .ZN(MEM_stage_inst_dmem_n19547) );
NAND2_X1 MEM_stage_inst_dmem_U18670 ( .A1(MEM_stage_inst_dmem_ram_3471), .A2(MEM_stage_inst_dmem_n19546), .ZN(MEM_stage_inst_dmem_n19517) );
NAND2_X1 MEM_stage_inst_dmem_U18669 ( .A1(MEM_stage_inst_dmem_n21179), .A2(MEM_stage_inst_dmem_n19788), .ZN(MEM_stage_inst_dmem_n19546) );
NAND2_X1 MEM_stage_inst_dmem_U18668 ( .A1(MEM_stage_inst_dmem_n19515), .A2(MEM_stage_inst_dmem_n19514), .ZN(MEM_stage_inst_dmem_n9675) );
NAND2_X1 MEM_stage_inst_dmem_U18667 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n19513), .ZN(MEM_stage_inst_dmem_n19514) );
NAND2_X1 MEM_stage_inst_dmem_U18666 ( .A1(MEM_stage_inst_dmem_ram_3472), .A2(MEM_stage_inst_dmem_n19512), .ZN(MEM_stage_inst_dmem_n19515) );
NAND2_X1 MEM_stage_inst_dmem_U18665 ( .A1(MEM_stage_inst_dmem_n19511), .A2(MEM_stage_inst_dmem_n19510), .ZN(MEM_stage_inst_dmem_n9676) );
NAND2_X1 MEM_stage_inst_dmem_U18664 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n19513), .ZN(MEM_stage_inst_dmem_n19510) );
NAND2_X1 MEM_stage_inst_dmem_U18663 ( .A1(MEM_stage_inst_dmem_ram_3473), .A2(MEM_stage_inst_dmem_n19512), .ZN(MEM_stage_inst_dmem_n19511) );
NAND2_X1 MEM_stage_inst_dmem_U18662 ( .A1(MEM_stage_inst_dmem_n19509), .A2(MEM_stage_inst_dmem_n19508), .ZN(MEM_stage_inst_dmem_n9677) );
NAND2_X1 MEM_stage_inst_dmem_U18661 ( .A1(MEM_stage_inst_dmem_n18027), .A2(MEM_stage_inst_dmem_n19513), .ZN(MEM_stage_inst_dmem_n19508) );
NAND2_X1 MEM_stage_inst_dmem_U18660 ( .A1(MEM_stage_inst_dmem_ram_3474), .A2(MEM_stage_inst_dmem_n19512), .ZN(MEM_stage_inst_dmem_n19509) );
NAND2_X1 MEM_stage_inst_dmem_U18659 ( .A1(MEM_stage_inst_dmem_n19507), .A2(MEM_stage_inst_dmem_n19506), .ZN(MEM_stage_inst_dmem_n9678) );
NAND2_X1 MEM_stage_inst_dmem_U18658 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n19513), .ZN(MEM_stage_inst_dmem_n19506) );
NAND2_X1 MEM_stage_inst_dmem_U18657 ( .A1(MEM_stage_inst_dmem_ram_3475), .A2(MEM_stage_inst_dmem_n19512), .ZN(MEM_stage_inst_dmem_n19507) );
NAND2_X1 MEM_stage_inst_dmem_U18656 ( .A1(MEM_stage_inst_dmem_n19505), .A2(MEM_stage_inst_dmem_n19504), .ZN(MEM_stage_inst_dmem_n9679) );
NAND2_X1 MEM_stage_inst_dmem_U18655 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n19513), .ZN(MEM_stage_inst_dmem_n19504) );
NAND2_X1 MEM_stage_inst_dmem_U18654 ( .A1(MEM_stage_inst_dmem_ram_3476), .A2(MEM_stage_inst_dmem_n19512), .ZN(MEM_stage_inst_dmem_n19505) );
NAND2_X1 MEM_stage_inst_dmem_U18653 ( .A1(MEM_stage_inst_dmem_n19503), .A2(MEM_stage_inst_dmem_n19502), .ZN(MEM_stage_inst_dmem_n9680) );
NAND2_X1 MEM_stage_inst_dmem_U18652 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n19513), .ZN(MEM_stage_inst_dmem_n19502) );
NAND2_X1 MEM_stage_inst_dmem_U18651 ( .A1(MEM_stage_inst_dmem_ram_3477), .A2(MEM_stage_inst_dmem_n19512), .ZN(MEM_stage_inst_dmem_n19503) );
NAND2_X1 MEM_stage_inst_dmem_U18650 ( .A1(MEM_stage_inst_dmem_n19501), .A2(MEM_stage_inst_dmem_n19500), .ZN(MEM_stage_inst_dmem_n9681) );
NAND2_X1 MEM_stage_inst_dmem_U18649 ( .A1(EX_pipeline_reg_out_11), .A2(MEM_stage_inst_dmem_n19513), .ZN(MEM_stage_inst_dmem_n19500) );
NAND2_X1 MEM_stage_inst_dmem_U18648 ( .A1(MEM_stage_inst_dmem_ram_3478), .A2(MEM_stage_inst_dmem_n19512), .ZN(MEM_stage_inst_dmem_n19501) );
NAND2_X1 MEM_stage_inst_dmem_U18647 ( .A1(MEM_stage_inst_dmem_n19499), .A2(MEM_stage_inst_dmem_n19498), .ZN(MEM_stage_inst_dmem_n9682) );
NAND2_X1 MEM_stage_inst_dmem_U18646 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n19513), .ZN(MEM_stage_inst_dmem_n19498) );
NAND2_X1 MEM_stage_inst_dmem_U18645 ( .A1(MEM_stage_inst_dmem_ram_3479), .A2(MEM_stage_inst_dmem_n19512), .ZN(MEM_stage_inst_dmem_n19499) );
NAND2_X1 MEM_stage_inst_dmem_U18644 ( .A1(MEM_stage_inst_dmem_n19497), .A2(MEM_stage_inst_dmem_n19496), .ZN(MEM_stage_inst_dmem_n9683) );
NAND2_X1 MEM_stage_inst_dmem_U18643 ( .A1(MEM_stage_inst_dmem_n21335), .A2(MEM_stage_inst_dmem_n19513), .ZN(MEM_stage_inst_dmem_n19496) );
NAND2_X1 MEM_stage_inst_dmem_U18642 ( .A1(MEM_stage_inst_dmem_ram_3480), .A2(MEM_stage_inst_dmem_n19512), .ZN(MEM_stage_inst_dmem_n19497) );
NAND2_X1 MEM_stage_inst_dmem_U18641 ( .A1(MEM_stage_inst_dmem_n19495), .A2(MEM_stage_inst_dmem_n19494), .ZN(MEM_stage_inst_dmem_n9684) );
NAND2_X1 MEM_stage_inst_dmem_U18640 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n19513), .ZN(MEM_stage_inst_dmem_n19494) );
NAND2_X1 MEM_stage_inst_dmem_U18639 ( .A1(MEM_stage_inst_dmem_ram_3481), .A2(MEM_stage_inst_dmem_n19512), .ZN(MEM_stage_inst_dmem_n19495) );
NAND2_X1 MEM_stage_inst_dmem_U18638 ( .A1(MEM_stage_inst_dmem_n19493), .A2(MEM_stage_inst_dmem_n19492), .ZN(MEM_stage_inst_dmem_n9685) );
NAND2_X1 MEM_stage_inst_dmem_U18637 ( .A1(MEM_stage_inst_dmem_n18007), .A2(MEM_stage_inst_dmem_n19513), .ZN(MEM_stage_inst_dmem_n19492) );
NAND2_X1 MEM_stage_inst_dmem_U18636 ( .A1(MEM_stage_inst_dmem_ram_3482), .A2(MEM_stage_inst_dmem_n19512), .ZN(MEM_stage_inst_dmem_n19493) );
NAND2_X1 MEM_stage_inst_dmem_U18635 ( .A1(MEM_stage_inst_dmem_n19491), .A2(MEM_stage_inst_dmem_n19490), .ZN(MEM_stage_inst_dmem_n9686) );
NAND2_X1 MEM_stage_inst_dmem_U18634 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n19513), .ZN(MEM_stage_inst_dmem_n19490) );
NAND2_X1 MEM_stage_inst_dmem_U18633 ( .A1(MEM_stage_inst_dmem_ram_3483), .A2(MEM_stage_inst_dmem_n19512), .ZN(MEM_stage_inst_dmem_n19491) );
NAND2_X1 MEM_stage_inst_dmem_U18632 ( .A1(MEM_stage_inst_dmem_n19489), .A2(MEM_stage_inst_dmem_n19488), .ZN(MEM_stage_inst_dmem_n9687) );
NAND2_X1 MEM_stage_inst_dmem_U18631 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n19513), .ZN(MEM_stage_inst_dmem_n19488) );
NAND2_X1 MEM_stage_inst_dmem_U18630 ( .A1(MEM_stage_inst_dmem_ram_3484), .A2(MEM_stage_inst_dmem_n19512), .ZN(MEM_stage_inst_dmem_n19489) );
NAND2_X1 MEM_stage_inst_dmem_U18629 ( .A1(MEM_stage_inst_dmem_n19487), .A2(MEM_stage_inst_dmem_n19486), .ZN(MEM_stage_inst_dmem_n9688) );
NAND2_X1 MEM_stage_inst_dmem_U18628 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n19513), .ZN(MEM_stage_inst_dmem_n19486) );
NAND2_X1 MEM_stage_inst_dmem_U18627 ( .A1(MEM_stage_inst_dmem_ram_3485), .A2(MEM_stage_inst_dmem_n19512), .ZN(MEM_stage_inst_dmem_n19487) );
NAND2_X1 MEM_stage_inst_dmem_U18626 ( .A1(MEM_stage_inst_dmem_n19485), .A2(MEM_stage_inst_dmem_n19484), .ZN(MEM_stage_inst_dmem_n9689) );
NAND2_X1 MEM_stage_inst_dmem_U18625 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n19513), .ZN(MEM_stage_inst_dmem_n19484) );
NAND2_X1 MEM_stage_inst_dmem_U18624 ( .A1(MEM_stage_inst_dmem_ram_3486), .A2(MEM_stage_inst_dmem_n19512), .ZN(MEM_stage_inst_dmem_n19485) );
NAND2_X1 MEM_stage_inst_dmem_U18623 ( .A1(MEM_stage_inst_dmem_n19483), .A2(MEM_stage_inst_dmem_n19482), .ZN(MEM_stage_inst_dmem_n9690) );
NAND2_X1 MEM_stage_inst_dmem_U18622 ( .A1(MEM_stage_inst_dmem_n14693), .A2(MEM_stage_inst_dmem_n19513), .ZN(MEM_stage_inst_dmem_n19482) );
INV_X1 MEM_stage_inst_dmem_U18621 ( .A(MEM_stage_inst_dmem_n19512), .ZN(MEM_stage_inst_dmem_n19513) );
NAND2_X1 MEM_stage_inst_dmem_U18620 ( .A1(MEM_stage_inst_dmem_ram_3487), .A2(MEM_stage_inst_dmem_n19512), .ZN(MEM_stage_inst_dmem_n19483) );
NAND2_X1 MEM_stage_inst_dmem_U18619 ( .A1(MEM_stage_inst_dmem_n21144), .A2(MEM_stage_inst_dmem_n19788), .ZN(MEM_stage_inst_dmem_n19512) );
NAND2_X1 MEM_stage_inst_dmem_U18618 ( .A1(MEM_stage_inst_dmem_n19481), .A2(MEM_stage_inst_dmem_n19480), .ZN(MEM_stage_inst_dmem_n9691) );
NAND2_X1 MEM_stage_inst_dmem_U18617 ( .A1(MEM_stage_inst_dmem_n20551), .A2(MEM_stage_inst_dmem_n19479), .ZN(MEM_stage_inst_dmem_n19480) );
NAND2_X1 MEM_stage_inst_dmem_U18616 ( .A1(MEM_stage_inst_dmem_ram_3488), .A2(MEM_stage_inst_dmem_n19478), .ZN(MEM_stage_inst_dmem_n19481) );
NAND2_X1 MEM_stage_inst_dmem_U18615 ( .A1(MEM_stage_inst_dmem_n19477), .A2(MEM_stage_inst_dmem_n19476), .ZN(MEM_stage_inst_dmem_n9692) );
NAND2_X1 MEM_stage_inst_dmem_U18614 ( .A1(MEM_stage_inst_dmem_n20547), .A2(MEM_stage_inst_dmem_n19479), .ZN(MEM_stage_inst_dmem_n19476) );
NAND2_X1 MEM_stage_inst_dmem_U18613 ( .A1(MEM_stage_inst_dmem_ram_3489), .A2(MEM_stage_inst_dmem_n19478), .ZN(MEM_stage_inst_dmem_n19477) );
NAND2_X1 MEM_stage_inst_dmem_U18612 ( .A1(MEM_stage_inst_dmem_n19475), .A2(MEM_stage_inst_dmem_n19474), .ZN(MEM_stage_inst_dmem_n9693) );
NAND2_X1 MEM_stage_inst_dmem_U18611 ( .A1(MEM_stage_inst_dmem_n20544), .A2(MEM_stage_inst_dmem_n19479), .ZN(MEM_stage_inst_dmem_n19474) );
NAND2_X1 MEM_stage_inst_dmem_U18610 ( .A1(MEM_stage_inst_dmem_ram_3490), .A2(MEM_stage_inst_dmem_n19478), .ZN(MEM_stage_inst_dmem_n19475) );
NAND2_X1 MEM_stage_inst_dmem_U18609 ( .A1(MEM_stage_inst_dmem_n19473), .A2(MEM_stage_inst_dmem_n19472), .ZN(MEM_stage_inst_dmem_n9694) );
NAND2_X1 MEM_stage_inst_dmem_U18608 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n19479), .ZN(MEM_stage_inst_dmem_n19472) );
NAND2_X1 MEM_stage_inst_dmem_U18607 ( .A1(MEM_stage_inst_dmem_ram_3491), .A2(MEM_stage_inst_dmem_n19478), .ZN(MEM_stage_inst_dmem_n19473) );
NAND2_X1 MEM_stage_inst_dmem_U18606 ( .A1(MEM_stage_inst_dmem_n19471), .A2(MEM_stage_inst_dmem_n19470), .ZN(MEM_stage_inst_dmem_n9695) );
NAND2_X1 MEM_stage_inst_dmem_U18605 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n19479), .ZN(MEM_stage_inst_dmem_n19470) );
NAND2_X1 MEM_stage_inst_dmem_U18604 ( .A1(MEM_stage_inst_dmem_ram_3492), .A2(MEM_stage_inst_dmem_n19478), .ZN(MEM_stage_inst_dmem_n19471) );
NAND2_X1 MEM_stage_inst_dmem_U18603 ( .A1(MEM_stage_inst_dmem_n19469), .A2(MEM_stage_inst_dmem_n19468), .ZN(MEM_stage_inst_dmem_n9696) );
NAND2_X1 MEM_stage_inst_dmem_U18602 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n19479), .ZN(MEM_stage_inst_dmem_n19468) );
NAND2_X1 MEM_stage_inst_dmem_U18601 ( .A1(MEM_stage_inst_dmem_ram_3493), .A2(MEM_stage_inst_dmem_n19478), .ZN(MEM_stage_inst_dmem_n19469) );
NAND2_X1 MEM_stage_inst_dmem_U18600 ( .A1(MEM_stage_inst_dmem_n19467), .A2(MEM_stage_inst_dmem_n19466), .ZN(MEM_stage_inst_dmem_n9697) );
NAND2_X1 MEM_stage_inst_dmem_U18599 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n19479), .ZN(MEM_stage_inst_dmem_n19466) );
NAND2_X1 MEM_stage_inst_dmem_U18598 ( .A1(MEM_stage_inst_dmem_ram_3494), .A2(MEM_stage_inst_dmem_n19478), .ZN(MEM_stage_inst_dmem_n19467) );
NAND2_X1 MEM_stage_inst_dmem_U18597 ( .A1(MEM_stage_inst_dmem_n19465), .A2(MEM_stage_inst_dmem_n19464), .ZN(MEM_stage_inst_dmem_n9698) );
NAND2_X1 MEM_stage_inst_dmem_U18596 ( .A1(MEM_stage_inst_dmem_n20530), .A2(MEM_stage_inst_dmem_n19479), .ZN(MEM_stage_inst_dmem_n19464) );
NAND2_X1 MEM_stage_inst_dmem_U18595 ( .A1(MEM_stage_inst_dmem_ram_3495), .A2(MEM_stage_inst_dmem_n19478), .ZN(MEM_stage_inst_dmem_n19465) );
NAND2_X1 MEM_stage_inst_dmem_U18594 ( .A1(MEM_stage_inst_dmem_n19463), .A2(MEM_stage_inst_dmem_n19462), .ZN(MEM_stage_inst_dmem_n9699) );
NAND2_X1 MEM_stage_inst_dmem_U18593 ( .A1(MEM_stage_inst_dmem_n20527), .A2(MEM_stage_inst_dmem_n19479), .ZN(MEM_stage_inst_dmem_n19462) );
NAND2_X1 MEM_stage_inst_dmem_U18592 ( .A1(MEM_stage_inst_dmem_ram_3496), .A2(MEM_stage_inst_dmem_n19478), .ZN(MEM_stage_inst_dmem_n19463) );
NAND2_X1 MEM_stage_inst_dmem_U18591 ( .A1(MEM_stage_inst_dmem_n19461), .A2(MEM_stage_inst_dmem_n19460), .ZN(MEM_stage_inst_dmem_n9700) );
NAND2_X1 MEM_stage_inst_dmem_U18590 ( .A1(MEM_stage_inst_dmem_n20524), .A2(MEM_stage_inst_dmem_n19479), .ZN(MEM_stage_inst_dmem_n19460) );
NAND2_X1 MEM_stage_inst_dmem_U18589 ( .A1(MEM_stage_inst_dmem_ram_3497), .A2(MEM_stage_inst_dmem_n19478), .ZN(MEM_stage_inst_dmem_n19461) );
NAND2_X1 MEM_stage_inst_dmem_U18588 ( .A1(MEM_stage_inst_dmem_n19459), .A2(MEM_stage_inst_dmem_n19458), .ZN(MEM_stage_inst_dmem_n9701) );
NAND2_X1 MEM_stage_inst_dmem_U18587 ( .A1(MEM_stage_inst_dmem_n20521), .A2(MEM_stage_inst_dmem_n19479), .ZN(MEM_stage_inst_dmem_n19458) );
NAND2_X1 MEM_stage_inst_dmem_U18586 ( .A1(MEM_stage_inst_dmem_ram_3498), .A2(MEM_stage_inst_dmem_n19478), .ZN(MEM_stage_inst_dmem_n19459) );
NAND2_X1 MEM_stage_inst_dmem_U18585 ( .A1(MEM_stage_inst_dmem_n19457), .A2(MEM_stage_inst_dmem_n19456), .ZN(MEM_stage_inst_dmem_n9702) );
NAND2_X1 MEM_stage_inst_dmem_U18584 ( .A1(MEM_stage_inst_dmem_n20518), .A2(MEM_stage_inst_dmem_n19479), .ZN(MEM_stage_inst_dmem_n19456) );
NAND2_X1 MEM_stage_inst_dmem_U18583 ( .A1(MEM_stage_inst_dmem_ram_3499), .A2(MEM_stage_inst_dmem_n19478), .ZN(MEM_stage_inst_dmem_n19457) );
NAND2_X1 MEM_stage_inst_dmem_U18582 ( .A1(MEM_stage_inst_dmem_n19455), .A2(MEM_stage_inst_dmem_n19454), .ZN(MEM_stage_inst_dmem_n9703) );
NAND2_X1 MEM_stage_inst_dmem_U18581 ( .A1(MEM_stage_inst_dmem_n20515), .A2(MEM_stage_inst_dmem_n19479), .ZN(MEM_stage_inst_dmem_n19454) );
NAND2_X1 MEM_stage_inst_dmem_U18580 ( .A1(MEM_stage_inst_dmem_ram_3500), .A2(MEM_stage_inst_dmem_n19478), .ZN(MEM_stage_inst_dmem_n19455) );
NAND2_X1 MEM_stage_inst_dmem_U18579 ( .A1(MEM_stage_inst_dmem_n19453), .A2(MEM_stage_inst_dmem_n19452), .ZN(MEM_stage_inst_dmem_n9704) );
NAND2_X1 MEM_stage_inst_dmem_U18578 ( .A1(MEM_stage_inst_dmem_n20512), .A2(MEM_stage_inst_dmem_n19479), .ZN(MEM_stage_inst_dmem_n19452) );
NAND2_X1 MEM_stage_inst_dmem_U18577 ( .A1(MEM_stage_inst_dmem_ram_3501), .A2(MEM_stage_inst_dmem_n19478), .ZN(MEM_stage_inst_dmem_n19453) );
NAND2_X1 MEM_stage_inst_dmem_U18576 ( .A1(MEM_stage_inst_dmem_n19451), .A2(MEM_stage_inst_dmem_n19450), .ZN(MEM_stage_inst_dmem_n9705) );
NAND2_X1 MEM_stage_inst_dmem_U18575 ( .A1(MEM_stage_inst_dmem_n20509), .A2(MEM_stage_inst_dmem_n19479), .ZN(MEM_stage_inst_dmem_n19450) );
NAND2_X1 MEM_stage_inst_dmem_U18574 ( .A1(MEM_stage_inst_dmem_ram_3502), .A2(MEM_stage_inst_dmem_n19478), .ZN(MEM_stage_inst_dmem_n19451) );
NAND2_X1 MEM_stage_inst_dmem_U18573 ( .A1(MEM_stage_inst_dmem_n19449), .A2(MEM_stage_inst_dmem_n19448), .ZN(MEM_stage_inst_dmem_n9706) );
NAND2_X1 MEM_stage_inst_dmem_U18572 ( .A1(MEM_stage_inst_dmem_n20506), .A2(MEM_stage_inst_dmem_n19479), .ZN(MEM_stage_inst_dmem_n19448) );
INV_X1 MEM_stage_inst_dmem_U18571 ( .A(MEM_stage_inst_dmem_n19478), .ZN(MEM_stage_inst_dmem_n19479) );
NAND2_X1 MEM_stage_inst_dmem_U18570 ( .A1(MEM_stage_inst_dmem_ram_3503), .A2(MEM_stage_inst_dmem_n19478), .ZN(MEM_stage_inst_dmem_n19449) );
NAND2_X1 MEM_stage_inst_dmem_U18569 ( .A1(MEM_stage_inst_dmem_n21109), .A2(MEM_stage_inst_dmem_n19788), .ZN(MEM_stage_inst_dmem_n19478) );
NAND2_X1 MEM_stage_inst_dmem_U18568 ( .A1(MEM_stage_inst_dmem_n19447), .A2(MEM_stage_inst_dmem_n19446), .ZN(MEM_stage_inst_dmem_n9707) );
NAND2_X1 MEM_stage_inst_dmem_U18567 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n19445), .ZN(MEM_stage_inst_dmem_n19446) );
NAND2_X1 MEM_stage_inst_dmem_U18566 ( .A1(MEM_stage_inst_dmem_ram_3504), .A2(MEM_stage_inst_dmem_n19444), .ZN(MEM_stage_inst_dmem_n19447) );
NAND2_X1 MEM_stage_inst_dmem_U18565 ( .A1(MEM_stage_inst_dmem_n19443), .A2(MEM_stage_inst_dmem_n19442), .ZN(MEM_stage_inst_dmem_n9708) );
NAND2_X1 MEM_stage_inst_dmem_U18564 ( .A1(MEM_stage_inst_dmem_n109), .A2(MEM_stage_inst_dmem_n19445), .ZN(MEM_stage_inst_dmem_n19442) );
NAND2_X1 MEM_stage_inst_dmem_U18563 ( .A1(MEM_stage_inst_dmem_ram_3505), .A2(MEM_stage_inst_dmem_n19444), .ZN(MEM_stage_inst_dmem_n19443) );
NAND2_X1 MEM_stage_inst_dmem_U18562 ( .A1(MEM_stage_inst_dmem_n19441), .A2(MEM_stage_inst_dmem_n19440), .ZN(MEM_stage_inst_dmem_n9709) );
NAND2_X1 MEM_stage_inst_dmem_U18561 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n19445), .ZN(MEM_stage_inst_dmem_n19440) );
NAND2_X1 MEM_stage_inst_dmem_U18560 ( .A1(MEM_stage_inst_dmem_ram_3506), .A2(MEM_stage_inst_dmem_n19444), .ZN(MEM_stage_inst_dmem_n19441) );
NAND2_X1 MEM_stage_inst_dmem_U18559 ( .A1(MEM_stage_inst_dmem_n19439), .A2(MEM_stage_inst_dmem_n19438), .ZN(MEM_stage_inst_dmem_n9710) );
NAND2_X1 MEM_stage_inst_dmem_U18558 ( .A1(MEM_stage_inst_dmem_n13064), .A2(MEM_stage_inst_dmem_n19445), .ZN(MEM_stage_inst_dmem_n19438) );
NAND2_X1 MEM_stage_inst_dmem_U18557 ( .A1(MEM_stage_inst_dmem_ram_3507), .A2(MEM_stage_inst_dmem_n19444), .ZN(MEM_stage_inst_dmem_n19439) );
NAND2_X1 MEM_stage_inst_dmem_U18556 ( .A1(MEM_stage_inst_dmem_n19437), .A2(MEM_stage_inst_dmem_n19436), .ZN(MEM_stage_inst_dmem_n9711) );
NAND2_X1 MEM_stage_inst_dmem_U18555 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n19445), .ZN(MEM_stage_inst_dmem_n19436) );
NAND2_X1 MEM_stage_inst_dmem_U18554 ( .A1(MEM_stage_inst_dmem_ram_3508), .A2(MEM_stage_inst_dmem_n19444), .ZN(MEM_stage_inst_dmem_n19437) );
NAND2_X1 MEM_stage_inst_dmem_U18553 ( .A1(MEM_stage_inst_dmem_n19435), .A2(MEM_stage_inst_dmem_n19434), .ZN(MEM_stage_inst_dmem_n9712) );
NAND2_X1 MEM_stage_inst_dmem_U18552 ( .A1(MEM_stage_inst_dmem_n13059), .A2(MEM_stage_inst_dmem_n19445), .ZN(MEM_stage_inst_dmem_n19434) );
NAND2_X1 MEM_stage_inst_dmem_U18551 ( .A1(MEM_stage_inst_dmem_ram_3509), .A2(MEM_stage_inst_dmem_n19444), .ZN(MEM_stage_inst_dmem_n19435) );
NAND2_X1 MEM_stage_inst_dmem_U18550 ( .A1(MEM_stage_inst_dmem_n19433), .A2(MEM_stage_inst_dmem_n19432), .ZN(MEM_stage_inst_dmem_n9713) );
NAND2_X1 MEM_stage_inst_dmem_U18549 ( .A1(MEM_stage_inst_dmem_n13056), .A2(MEM_stage_inst_dmem_n19445), .ZN(MEM_stage_inst_dmem_n19432) );
NAND2_X1 MEM_stage_inst_dmem_U18548 ( .A1(MEM_stage_inst_dmem_ram_3510), .A2(MEM_stage_inst_dmem_n19444), .ZN(MEM_stage_inst_dmem_n19433) );
NAND2_X1 MEM_stage_inst_dmem_U18547 ( .A1(MEM_stage_inst_dmem_n19431), .A2(MEM_stage_inst_dmem_n19430), .ZN(MEM_stage_inst_dmem_n9714) );
NAND2_X1 MEM_stage_inst_dmem_U18546 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n19445), .ZN(MEM_stage_inst_dmem_n19430) );
NAND2_X1 MEM_stage_inst_dmem_U18545 ( .A1(MEM_stage_inst_dmem_ram_3511), .A2(MEM_stage_inst_dmem_n19444), .ZN(MEM_stage_inst_dmem_n19431) );
NAND2_X1 MEM_stage_inst_dmem_U18544 ( .A1(MEM_stage_inst_dmem_n19429), .A2(MEM_stage_inst_dmem_n19428), .ZN(MEM_stage_inst_dmem_n9715) );
NAND2_X1 MEM_stage_inst_dmem_U18543 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n19445), .ZN(MEM_stage_inst_dmem_n19428) );
NAND2_X1 MEM_stage_inst_dmem_U18542 ( .A1(MEM_stage_inst_dmem_ram_3512), .A2(MEM_stage_inst_dmem_n19444), .ZN(MEM_stage_inst_dmem_n19429) );
NAND2_X1 MEM_stage_inst_dmem_U18541 ( .A1(MEM_stage_inst_dmem_n19427), .A2(MEM_stage_inst_dmem_n19426), .ZN(MEM_stage_inst_dmem_n9716) );
NAND2_X1 MEM_stage_inst_dmem_U18540 ( .A1(MEM_stage_inst_dmem_n16772), .A2(MEM_stage_inst_dmem_n19445), .ZN(MEM_stage_inst_dmem_n19426) );
NAND2_X1 MEM_stage_inst_dmem_U18539 ( .A1(MEM_stage_inst_dmem_ram_3513), .A2(MEM_stage_inst_dmem_n19444), .ZN(MEM_stage_inst_dmem_n19427) );
NAND2_X1 MEM_stage_inst_dmem_U18538 ( .A1(MEM_stage_inst_dmem_n19425), .A2(MEM_stage_inst_dmem_n19424), .ZN(MEM_stage_inst_dmem_n9717) );
NAND2_X1 MEM_stage_inst_dmem_U18537 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n19445), .ZN(MEM_stage_inst_dmem_n19424) );
NAND2_X1 MEM_stage_inst_dmem_U18536 ( .A1(MEM_stage_inst_dmem_ram_3514), .A2(MEM_stage_inst_dmem_n19444), .ZN(MEM_stage_inst_dmem_n19425) );
NAND2_X1 MEM_stage_inst_dmem_U18535 ( .A1(MEM_stage_inst_dmem_n19423), .A2(MEM_stage_inst_dmem_n19422), .ZN(MEM_stage_inst_dmem_n9718) );
NAND2_X1 MEM_stage_inst_dmem_U18534 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n19445), .ZN(MEM_stage_inst_dmem_n19422) );
NAND2_X1 MEM_stage_inst_dmem_U18533 ( .A1(MEM_stage_inst_dmem_ram_3515), .A2(MEM_stage_inst_dmem_n19444), .ZN(MEM_stage_inst_dmem_n19423) );
NAND2_X1 MEM_stage_inst_dmem_U18532 ( .A1(MEM_stage_inst_dmem_n19421), .A2(MEM_stage_inst_dmem_n19420), .ZN(MEM_stage_inst_dmem_n9719) );
NAND2_X1 MEM_stage_inst_dmem_U18531 ( .A1(MEM_stage_inst_dmem_n14702), .A2(MEM_stage_inst_dmem_n19445), .ZN(MEM_stage_inst_dmem_n19420) );
NAND2_X1 MEM_stage_inst_dmem_U18530 ( .A1(MEM_stage_inst_dmem_ram_3516), .A2(MEM_stage_inst_dmem_n19444), .ZN(MEM_stage_inst_dmem_n19421) );
NAND2_X1 MEM_stage_inst_dmem_U18529 ( .A1(MEM_stage_inst_dmem_n19419), .A2(MEM_stage_inst_dmem_n19418), .ZN(MEM_stage_inst_dmem_n9720) );
NAND2_X1 MEM_stage_inst_dmem_U18528 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n19445), .ZN(MEM_stage_inst_dmem_n19418) );
NAND2_X1 MEM_stage_inst_dmem_U18527 ( .A1(MEM_stage_inst_dmem_ram_3517), .A2(MEM_stage_inst_dmem_n19444), .ZN(MEM_stage_inst_dmem_n19419) );
NAND2_X1 MEM_stage_inst_dmem_U18526 ( .A1(MEM_stage_inst_dmem_n19417), .A2(MEM_stage_inst_dmem_n19416), .ZN(MEM_stage_inst_dmem_n9721) );
NAND2_X1 MEM_stage_inst_dmem_U18525 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n19445), .ZN(MEM_stage_inst_dmem_n19416) );
NAND2_X1 MEM_stage_inst_dmem_U18524 ( .A1(MEM_stage_inst_dmem_ram_3518), .A2(MEM_stage_inst_dmem_n19444), .ZN(MEM_stage_inst_dmem_n19417) );
NAND2_X1 MEM_stage_inst_dmem_U18523 ( .A1(MEM_stage_inst_dmem_n19415), .A2(MEM_stage_inst_dmem_n19414), .ZN(MEM_stage_inst_dmem_n9722) );
NAND2_X1 MEM_stage_inst_dmem_U18522 ( .A1(MEM_stage_inst_dmem_n20506), .A2(MEM_stage_inst_dmem_n19445), .ZN(MEM_stage_inst_dmem_n19414) );
INV_X1 MEM_stage_inst_dmem_U18521 ( .A(MEM_stage_inst_dmem_n19444), .ZN(MEM_stage_inst_dmem_n19445) );
NAND2_X1 MEM_stage_inst_dmem_U18520 ( .A1(MEM_stage_inst_dmem_ram_3519), .A2(MEM_stage_inst_dmem_n19444), .ZN(MEM_stage_inst_dmem_n19415) );
NAND2_X1 MEM_stage_inst_dmem_U18519 ( .A1(MEM_stage_inst_dmem_n21074), .A2(MEM_stage_inst_dmem_n19788), .ZN(MEM_stage_inst_dmem_n19444) );
NAND2_X1 MEM_stage_inst_dmem_U18518 ( .A1(MEM_stage_inst_dmem_n19413), .A2(MEM_stage_inst_dmem_n19412), .ZN(MEM_stage_inst_dmem_n9723) );
NAND2_X1 MEM_stage_inst_dmem_U18517 ( .A1(MEM_stage_inst_dmem_n20551), .A2(MEM_stage_inst_dmem_n19411), .ZN(MEM_stage_inst_dmem_n19412) );
NAND2_X1 MEM_stage_inst_dmem_U18516 ( .A1(MEM_stage_inst_dmem_ram_3520), .A2(MEM_stage_inst_dmem_n19410), .ZN(MEM_stage_inst_dmem_n19413) );
NAND2_X1 MEM_stage_inst_dmem_U18515 ( .A1(MEM_stage_inst_dmem_n19409), .A2(MEM_stage_inst_dmem_n19408), .ZN(MEM_stage_inst_dmem_n9724) );
NAND2_X1 MEM_stage_inst_dmem_U18514 ( .A1(MEM_stage_inst_dmem_n20547), .A2(MEM_stage_inst_dmem_n19411), .ZN(MEM_stage_inst_dmem_n19408) );
NAND2_X1 MEM_stage_inst_dmem_U18513 ( .A1(MEM_stage_inst_dmem_ram_3521), .A2(MEM_stage_inst_dmem_n19410), .ZN(MEM_stage_inst_dmem_n19409) );
NAND2_X1 MEM_stage_inst_dmem_U18512 ( .A1(MEM_stage_inst_dmem_n19407), .A2(MEM_stage_inst_dmem_n19406), .ZN(MEM_stage_inst_dmem_n9725) );
NAND2_X1 MEM_stage_inst_dmem_U18511 ( .A1(MEM_stage_inst_dmem_n20544), .A2(MEM_stage_inst_dmem_n19411), .ZN(MEM_stage_inst_dmem_n19406) );
NAND2_X1 MEM_stage_inst_dmem_U18510 ( .A1(MEM_stage_inst_dmem_ram_3522), .A2(MEM_stage_inst_dmem_n19410), .ZN(MEM_stage_inst_dmem_n19407) );
NAND2_X1 MEM_stage_inst_dmem_U18509 ( .A1(MEM_stage_inst_dmem_n19405), .A2(MEM_stage_inst_dmem_n19404), .ZN(MEM_stage_inst_dmem_n9726) );
NAND2_X1 MEM_stage_inst_dmem_U18508 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n19411), .ZN(MEM_stage_inst_dmem_n19404) );
NAND2_X1 MEM_stage_inst_dmem_U18507 ( .A1(MEM_stage_inst_dmem_ram_3523), .A2(MEM_stage_inst_dmem_n19410), .ZN(MEM_stage_inst_dmem_n19405) );
NAND2_X1 MEM_stage_inst_dmem_U18506 ( .A1(MEM_stage_inst_dmem_n19403), .A2(MEM_stage_inst_dmem_n19402), .ZN(MEM_stage_inst_dmem_n9727) );
NAND2_X1 MEM_stage_inst_dmem_U18505 ( .A1(EX_pipeline_reg_out_9), .A2(MEM_stage_inst_dmem_n19411), .ZN(MEM_stage_inst_dmem_n19402) );
NAND2_X1 MEM_stage_inst_dmem_U18504 ( .A1(MEM_stage_inst_dmem_ram_3524), .A2(MEM_stage_inst_dmem_n19410), .ZN(MEM_stage_inst_dmem_n19403) );
NAND2_X1 MEM_stage_inst_dmem_U18503 ( .A1(MEM_stage_inst_dmem_n19401), .A2(MEM_stage_inst_dmem_n19400), .ZN(MEM_stage_inst_dmem_n9728) );
NAND2_X1 MEM_stage_inst_dmem_U18502 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n19411), .ZN(MEM_stage_inst_dmem_n19400) );
NAND2_X1 MEM_stage_inst_dmem_U18501 ( .A1(MEM_stage_inst_dmem_ram_3525), .A2(MEM_stage_inst_dmem_n19410), .ZN(MEM_stage_inst_dmem_n19401) );
NAND2_X1 MEM_stage_inst_dmem_U18500 ( .A1(MEM_stage_inst_dmem_n19399), .A2(MEM_stage_inst_dmem_n19398), .ZN(MEM_stage_inst_dmem_n9729) );
NAND2_X1 MEM_stage_inst_dmem_U18499 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n19411), .ZN(MEM_stage_inst_dmem_n19398) );
NAND2_X1 MEM_stage_inst_dmem_U18498 ( .A1(MEM_stage_inst_dmem_ram_3526), .A2(MEM_stage_inst_dmem_n19410), .ZN(MEM_stage_inst_dmem_n19399) );
NAND2_X1 MEM_stage_inst_dmem_U18497 ( .A1(MEM_stage_inst_dmem_n19397), .A2(MEM_stage_inst_dmem_n19396), .ZN(MEM_stage_inst_dmem_n9730) );
NAND2_X1 MEM_stage_inst_dmem_U18496 ( .A1(MEM_stage_inst_dmem_n20530), .A2(MEM_stage_inst_dmem_n19411), .ZN(MEM_stage_inst_dmem_n19396) );
NAND2_X1 MEM_stage_inst_dmem_U18495 ( .A1(MEM_stage_inst_dmem_ram_3527), .A2(MEM_stage_inst_dmem_n19410), .ZN(MEM_stage_inst_dmem_n19397) );
NAND2_X1 MEM_stage_inst_dmem_U18494 ( .A1(MEM_stage_inst_dmem_n19395), .A2(MEM_stage_inst_dmem_n19394), .ZN(MEM_stage_inst_dmem_n9731) );
NAND2_X1 MEM_stage_inst_dmem_U18493 ( .A1(MEM_stage_inst_dmem_n20527), .A2(MEM_stage_inst_dmem_n19411), .ZN(MEM_stage_inst_dmem_n19394) );
NAND2_X1 MEM_stage_inst_dmem_U18492 ( .A1(MEM_stage_inst_dmem_ram_3528), .A2(MEM_stage_inst_dmem_n19410), .ZN(MEM_stage_inst_dmem_n19395) );
NAND2_X1 MEM_stage_inst_dmem_U18491 ( .A1(MEM_stage_inst_dmem_n19393), .A2(MEM_stage_inst_dmem_n19392), .ZN(MEM_stage_inst_dmem_n9732) );
NAND2_X1 MEM_stage_inst_dmem_U18490 ( .A1(MEM_stage_inst_dmem_n20524), .A2(MEM_stage_inst_dmem_n19411), .ZN(MEM_stage_inst_dmem_n19392) );
NAND2_X1 MEM_stage_inst_dmem_U18489 ( .A1(MEM_stage_inst_dmem_ram_3529), .A2(MEM_stage_inst_dmem_n19410), .ZN(MEM_stage_inst_dmem_n19393) );
NAND2_X1 MEM_stage_inst_dmem_U18488 ( .A1(MEM_stage_inst_dmem_n19391), .A2(MEM_stage_inst_dmem_n19390), .ZN(MEM_stage_inst_dmem_n9733) );
NAND2_X1 MEM_stage_inst_dmem_U18487 ( .A1(MEM_stage_inst_dmem_n20521), .A2(MEM_stage_inst_dmem_n19411), .ZN(MEM_stage_inst_dmem_n19390) );
NAND2_X1 MEM_stage_inst_dmem_U18486 ( .A1(MEM_stage_inst_dmem_ram_3530), .A2(MEM_stage_inst_dmem_n19410), .ZN(MEM_stage_inst_dmem_n19391) );
NAND2_X1 MEM_stage_inst_dmem_U18485 ( .A1(MEM_stage_inst_dmem_n19389), .A2(MEM_stage_inst_dmem_n19388), .ZN(MEM_stage_inst_dmem_n9734) );
NAND2_X1 MEM_stage_inst_dmem_U18484 ( .A1(MEM_stage_inst_dmem_n20518), .A2(MEM_stage_inst_dmem_n19411), .ZN(MEM_stage_inst_dmem_n19388) );
NAND2_X1 MEM_stage_inst_dmem_U18483 ( .A1(MEM_stage_inst_dmem_ram_3531), .A2(MEM_stage_inst_dmem_n19410), .ZN(MEM_stage_inst_dmem_n19389) );
NAND2_X1 MEM_stage_inst_dmem_U18482 ( .A1(MEM_stage_inst_dmem_n19387), .A2(MEM_stage_inst_dmem_n19386), .ZN(MEM_stage_inst_dmem_n9735) );
NAND2_X1 MEM_stage_inst_dmem_U18481 ( .A1(MEM_stage_inst_dmem_n20515), .A2(MEM_stage_inst_dmem_n19411), .ZN(MEM_stage_inst_dmem_n19386) );
NAND2_X1 MEM_stage_inst_dmem_U18480 ( .A1(MEM_stage_inst_dmem_ram_3532), .A2(MEM_stage_inst_dmem_n19410), .ZN(MEM_stage_inst_dmem_n19387) );
NAND2_X1 MEM_stage_inst_dmem_U18479 ( .A1(MEM_stage_inst_dmem_n19385), .A2(MEM_stage_inst_dmem_n19384), .ZN(MEM_stage_inst_dmem_n9736) );
NAND2_X1 MEM_stage_inst_dmem_U18478 ( .A1(MEM_stage_inst_dmem_n20512), .A2(MEM_stage_inst_dmem_n19411), .ZN(MEM_stage_inst_dmem_n19384) );
NAND2_X1 MEM_stage_inst_dmem_U18477 ( .A1(MEM_stage_inst_dmem_ram_3533), .A2(MEM_stage_inst_dmem_n19410), .ZN(MEM_stage_inst_dmem_n19385) );
NAND2_X1 MEM_stage_inst_dmem_U18476 ( .A1(MEM_stage_inst_dmem_n19383), .A2(MEM_stage_inst_dmem_n19382), .ZN(MEM_stage_inst_dmem_n9737) );
NAND2_X1 MEM_stage_inst_dmem_U18475 ( .A1(MEM_stage_inst_dmem_n20509), .A2(MEM_stage_inst_dmem_n19411), .ZN(MEM_stage_inst_dmem_n19382) );
NAND2_X1 MEM_stage_inst_dmem_U18474 ( .A1(MEM_stage_inst_dmem_ram_3534), .A2(MEM_stage_inst_dmem_n19410), .ZN(MEM_stage_inst_dmem_n19383) );
NAND2_X1 MEM_stage_inst_dmem_U18473 ( .A1(MEM_stage_inst_dmem_n19381), .A2(MEM_stage_inst_dmem_n19380), .ZN(MEM_stage_inst_dmem_n9738) );
NAND2_X1 MEM_stage_inst_dmem_U18472 ( .A1(MEM_stage_inst_dmem_n20506), .A2(MEM_stage_inst_dmem_n19411), .ZN(MEM_stage_inst_dmem_n19380) );
INV_X1 MEM_stage_inst_dmem_U18471 ( .A(MEM_stage_inst_dmem_n19410), .ZN(MEM_stage_inst_dmem_n19411) );
NAND2_X1 MEM_stage_inst_dmem_U18470 ( .A1(MEM_stage_inst_dmem_ram_3535), .A2(MEM_stage_inst_dmem_n19410), .ZN(MEM_stage_inst_dmem_n19381) );
NAND2_X1 MEM_stage_inst_dmem_U18469 ( .A1(MEM_stage_inst_dmem_n21039), .A2(MEM_stage_inst_dmem_n19788), .ZN(MEM_stage_inst_dmem_n19410) );
NAND2_X1 MEM_stage_inst_dmem_U18468 ( .A1(MEM_stage_inst_dmem_n19379), .A2(MEM_stage_inst_dmem_n19378), .ZN(MEM_stage_inst_dmem_n9739) );
NAND2_X1 MEM_stage_inst_dmem_U18467 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n19377), .ZN(MEM_stage_inst_dmem_n19378) );
NAND2_X1 MEM_stage_inst_dmem_U18466 ( .A1(MEM_stage_inst_dmem_ram_3536), .A2(MEM_stage_inst_dmem_n19376), .ZN(MEM_stage_inst_dmem_n19379) );
NAND2_X1 MEM_stage_inst_dmem_U18465 ( .A1(MEM_stage_inst_dmem_n19375), .A2(MEM_stage_inst_dmem_n19374), .ZN(MEM_stage_inst_dmem_n9740) );
NAND2_X1 MEM_stage_inst_dmem_U18464 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n19377), .ZN(MEM_stage_inst_dmem_n19374) );
NAND2_X1 MEM_stage_inst_dmem_U18463 ( .A1(MEM_stage_inst_dmem_ram_3537), .A2(MEM_stage_inst_dmem_n19376), .ZN(MEM_stage_inst_dmem_n19375) );
NAND2_X1 MEM_stage_inst_dmem_U18462 ( .A1(MEM_stage_inst_dmem_n19373), .A2(MEM_stage_inst_dmem_n19372), .ZN(MEM_stage_inst_dmem_n9741) );
NAND2_X1 MEM_stage_inst_dmem_U18461 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n19377), .ZN(MEM_stage_inst_dmem_n19372) );
NAND2_X1 MEM_stage_inst_dmem_U18460 ( .A1(MEM_stage_inst_dmem_ram_3538), .A2(MEM_stage_inst_dmem_n19376), .ZN(MEM_stage_inst_dmem_n19373) );
NAND2_X1 MEM_stage_inst_dmem_U18459 ( .A1(MEM_stage_inst_dmem_n19371), .A2(MEM_stage_inst_dmem_n19370), .ZN(MEM_stage_inst_dmem_n9742) );
NAND2_X1 MEM_stage_inst_dmem_U18458 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n19377), .ZN(MEM_stage_inst_dmem_n19370) );
NAND2_X1 MEM_stage_inst_dmem_U18457 ( .A1(MEM_stage_inst_dmem_ram_3539), .A2(MEM_stage_inst_dmem_n19376), .ZN(MEM_stage_inst_dmem_n19371) );
NAND2_X1 MEM_stage_inst_dmem_U18456 ( .A1(MEM_stage_inst_dmem_n19369), .A2(MEM_stage_inst_dmem_n19368), .ZN(MEM_stage_inst_dmem_n9743) );
NAND2_X1 MEM_stage_inst_dmem_U18455 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n19377), .ZN(MEM_stage_inst_dmem_n19368) );
NAND2_X1 MEM_stage_inst_dmem_U18454 ( .A1(MEM_stage_inst_dmem_ram_3540), .A2(MEM_stage_inst_dmem_n19376), .ZN(MEM_stage_inst_dmem_n19369) );
NAND2_X1 MEM_stage_inst_dmem_U18453 ( .A1(MEM_stage_inst_dmem_n19367), .A2(MEM_stage_inst_dmem_n19366), .ZN(MEM_stage_inst_dmem_n9744) );
NAND2_X1 MEM_stage_inst_dmem_U18452 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n19377), .ZN(MEM_stage_inst_dmem_n19366) );
NAND2_X1 MEM_stage_inst_dmem_U18451 ( .A1(MEM_stage_inst_dmem_ram_3541), .A2(MEM_stage_inst_dmem_n19376), .ZN(MEM_stage_inst_dmem_n19367) );
NAND2_X1 MEM_stage_inst_dmem_U18450 ( .A1(MEM_stage_inst_dmem_n19365), .A2(MEM_stage_inst_dmem_n19364), .ZN(MEM_stage_inst_dmem_n9745) );
NAND2_X1 MEM_stage_inst_dmem_U18449 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n19377), .ZN(MEM_stage_inst_dmem_n19364) );
NAND2_X1 MEM_stage_inst_dmem_U18448 ( .A1(MEM_stage_inst_dmem_ram_3542), .A2(MEM_stage_inst_dmem_n19376), .ZN(MEM_stage_inst_dmem_n19365) );
NAND2_X1 MEM_stage_inst_dmem_U18447 ( .A1(MEM_stage_inst_dmem_n19363), .A2(MEM_stage_inst_dmem_n19362), .ZN(MEM_stage_inst_dmem_n9746) );
NAND2_X1 MEM_stage_inst_dmem_U18446 ( .A1(MEM_stage_inst_dmem_n16361), .A2(MEM_stage_inst_dmem_n19377), .ZN(MEM_stage_inst_dmem_n19362) );
NAND2_X1 MEM_stage_inst_dmem_U18445 ( .A1(MEM_stage_inst_dmem_ram_3543), .A2(MEM_stage_inst_dmem_n19376), .ZN(MEM_stage_inst_dmem_n19363) );
NAND2_X1 MEM_stage_inst_dmem_U18444 ( .A1(MEM_stage_inst_dmem_n19361), .A2(MEM_stage_inst_dmem_n19360), .ZN(MEM_stage_inst_dmem_n9747) );
NAND2_X1 MEM_stage_inst_dmem_U18443 ( .A1(MEM_stage_inst_dmem_n111), .A2(MEM_stage_inst_dmem_n19377), .ZN(MEM_stage_inst_dmem_n19360) );
NAND2_X1 MEM_stage_inst_dmem_U18442 ( .A1(MEM_stage_inst_dmem_ram_3544), .A2(MEM_stage_inst_dmem_n19376), .ZN(MEM_stage_inst_dmem_n19361) );
NAND2_X1 MEM_stage_inst_dmem_U18441 ( .A1(MEM_stage_inst_dmem_n19359), .A2(MEM_stage_inst_dmem_n19358), .ZN(MEM_stage_inst_dmem_n9748) );
NAND2_X1 MEM_stage_inst_dmem_U18440 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n19377), .ZN(MEM_stage_inst_dmem_n19358) );
NAND2_X1 MEM_stage_inst_dmem_U18439 ( .A1(MEM_stage_inst_dmem_ram_3545), .A2(MEM_stage_inst_dmem_n19376), .ZN(MEM_stage_inst_dmem_n19359) );
NAND2_X1 MEM_stage_inst_dmem_U18438 ( .A1(MEM_stage_inst_dmem_n19357), .A2(MEM_stage_inst_dmem_n19356), .ZN(MEM_stage_inst_dmem_n9749) );
NAND2_X1 MEM_stage_inst_dmem_U18437 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n19377), .ZN(MEM_stage_inst_dmem_n19356) );
NAND2_X1 MEM_stage_inst_dmem_U18436 ( .A1(MEM_stage_inst_dmem_ram_3546), .A2(MEM_stage_inst_dmem_n19376), .ZN(MEM_stage_inst_dmem_n19357) );
NAND2_X1 MEM_stage_inst_dmem_U18435 ( .A1(MEM_stage_inst_dmem_n19355), .A2(MEM_stage_inst_dmem_n19354), .ZN(MEM_stage_inst_dmem_n9750) );
NAND2_X1 MEM_stage_inst_dmem_U18434 ( .A1(MEM_stage_inst_dmem_n18864), .A2(MEM_stage_inst_dmem_n19377), .ZN(MEM_stage_inst_dmem_n19354) );
NAND2_X1 MEM_stage_inst_dmem_U18433 ( .A1(MEM_stage_inst_dmem_ram_3547), .A2(MEM_stage_inst_dmem_n19376), .ZN(MEM_stage_inst_dmem_n19355) );
NAND2_X1 MEM_stage_inst_dmem_U18432 ( .A1(MEM_stage_inst_dmem_n19353), .A2(MEM_stage_inst_dmem_n19352), .ZN(MEM_stage_inst_dmem_n9751) );
NAND2_X1 MEM_stage_inst_dmem_U18431 ( .A1(MEM_stage_inst_dmem_n18861), .A2(MEM_stage_inst_dmem_n19377), .ZN(MEM_stage_inst_dmem_n19352) );
NAND2_X1 MEM_stage_inst_dmem_U18430 ( .A1(MEM_stage_inst_dmem_ram_3548), .A2(MEM_stage_inst_dmem_n19376), .ZN(MEM_stage_inst_dmem_n19353) );
NAND2_X1 MEM_stage_inst_dmem_U18429 ( .A1(MEM_stage_inst_dmem_n19351), .A2(MEM_stage_inst_dmem_n19350), .ZN(MEM_stage_inst_dmem_n9752) );
NAND2_X1 MEM_stage_inst_dmem_U18428 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n19377), .ZN(MEM_stage_inst_dmem_n19350) );
NAND2_X1 MEM_stage_inst_dmem_U18427 ( .A1(MEM_stage_inst_dmem_ram_3549), .A2(MEM_stage_inst_dmem_n19376), .ZN(MEM_stage_inst_dmem_n19351) );
NAND2_X1 MEM_stage_inst_dmem_U18426 ( .A1(MEM_stage_inst_dmem_n19349), .A2(MEM_stage_inst_dmem_n19348), .ZN(MEM_stage_inst_dmem_n9753) );
NAND2_X1 MEM_stage_inst_dmem_U18425 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n19377), .ZN(MEM_stage_inst_dmem_n19348) );
NAND2_X1 MEM_stage_inst_dmem_U18424 ( .A1(MEM_stage_inst_dmem_ram_3550), .A2(MEM_stage_inst_dmem_n19376), .ZN(MEM_stage_inst_dmem_n19349) );
NAND2_X1 MEM_stage_inst_dmem_U18423 ( .A1(MEM_stage_inst_dmem_n19347), .A2(MEM_stage_inst_dmem_n19346), .ZN(MEM_stage_inst_dmem_n9754) );
NAND2_X1 MEM_stage_inst_dmem_U18422 ( .A1(MEM_stage_inst_dmem_n16343), .A2(MEM_stage_inst_dmem_n19377), .ZN(MEM_stage_inst_dmem_n19346) );
INV_X1 MEM_stage_inst_dmem_U18421 ( .A(MEM_stage_inst_dmem_n19376), .ZN(MEM_stage_inst_dmem_n19377) );
NAND2_X1 MEM_stage_inst_dmem_U18420 ( .A1(MEM_stage_inst_dmem_ram_3551), .A2(MEM_stage_inst_dmem_n19376), .ZN(MEM_stage_inst_dmem_n19347) );
NAND2_X1 MEM_stage_inst_dmem_U18419 ( .A1(MEM_stage_inst_dmem_n21004), .A2(MEM_stage_inst_dmem_n19788), .ZN(MEM_stage_inst_dmem_n19376) );
NAND2_X1 MEM_stage_inst_dmem_U18418 ( .A1(MEM_stage_inst_dmem_n19345), .A2(MEM_stage_inst_dmem_n19344), .ZN(MEM_stage_inst_dmem_n9755) );
NAND2_X1 MEM_stage_inst_dmem_U18417 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n19343), .ZN(MEM_stage_inst_dmem_n19344) );
NAND2_X1 MEM_stage_inst_dmem_U18416 ( .A1(MEM_stage_inst_dmem_ram_3552), .A2(MEM_stage_inst_dmem_n19342), .ZN(MEM_stage_inst_dmem_n19345) );
NAND2_X1 MEM_stage_inst_dmem_U18415 ( .A1(MEM_stage_inst_dmem_n19341), .A2(MEM_stage_inst_dmem_n19340), .ZN(MEM_stage_inst_dmem_n9756) );
NAND2_X1 MEM_stage_inst_dmem_U18414 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n19343), .ZN(MEM_stage_inst_dmem_n19340) );
NAND2_X1 MEM_stage_inst_dmem_U18413 ( .A1(MEM_stage_inst_dmem_ram_3553), .A2(MEM_stage_inst_dmem_n19342), .ZN(MEM_stage_inst_dmem_n19341) );
NAND2_X1 MEM_stage_inst_dmem_U18412 ( .A1(MEM_stage_inst_dmem_n19339), .A2(MEM_stage_inst_dmem_n19338), .ZN(MEM_stage_inst_dmem_n9757) );
NAND2_X1 MEM_stage_inst_dmem_U18411 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n19343), .ZN(MEM_stage_inst_dmem_n19338) );
NAND2_X1 MEM_stage_inst_dmem_U18410 ( .A1(MEM_stage_inst_dmem_ram_3554), .A2(MEM_stage_inst_dmem_n19342), .ZN(MEM_stage_inst_dmem_n19339) );
NAND2_X1 MEM_stage_inst_dmem_U18409 ( .A1(MEM_stage_inst_dmem_n19337), .A2(MEM_stage_inst_dmem_n19336), .ZN(MEM_stage_inst_dmem_n9758) );
NAND2_X1 MEM_stage_inst_dmem_U18408 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n19343), .ZN(MEM_stage_inst_dmem_n19336) );
NAND2_X1 MEM_stage_inst_dmem_U18407 ( .A1(MEM_stage_inst_dmem_ram_3555), .A2(MEM_stage_inst_dmem_n19342), .ZN(MEM_stage_inst_dmem_n19337) );
NAND2_X1 MEM_stage_inst_dmem_U18406 ( .A1(MEM_stage_inst_dmem_n19335), .A2(MEM_stage_inst_dmem_n19334), .ZN(MEM_stage_inst_dmem_n9759) );
NAND2_X1 MEM_stage_inst_dmem_U18405 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n19343), .ZN(MEM_stage_inst_dmem_n19334) );
NAND2_X1 MEM_stage_inst_dmem_U18404 ( .A1(MEM_stage_inst_dmem_ram_3556), .A2(MEM_stage_inst_dmem_n19342), .ZN(MEM_stage_inst_dmem_n19335) );
NAND2_X1 MEM_stage_inst_dmem_U18403 ( .A1(MEM_stage_inst_dmem_n19333), .A2(MEM_stage_inst_dmem_n19332), .ZN(MEM_stage_inst_dmem_n9760) );
NAND2_X1 MEM_stage_inst_dmem_U18402 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n19343), .ZN(MEM_stage_inst_dmem_n19332) );
NAND2_X1 MEM_stage_inst_dmem_U18401 ( .A1(MEM_stage_inst_dmem_ram_3557), .A2(MEM_stage_inst_dmem_n19342), .ZN(MEM_stage_inst_dmem_n19333) );
NAND2_X1 MEM_stage_inst_dmem_U18400 ( .A1(MEM_stage_inst_dmem_n19331), .A2(MEM_stage_inst_dmem_n19330), .ZN(MEM_stage_inst_dmem_n9761) );
NAND2_X1 MEM_stage_inst_dmem_U18399 ( .A1(MEM_stage_inst_dmem_n21340), .A2(MEM_stage_inst_dmem_n19343), .ZN(MEM_stage_inst_dmem_n19330) );
NAND2_X1 MEM_stage_inst_dmem_U18398 ( .A1(MEM_stage_inst_dmem_ram_3558), .A2(MEM_stage_inst_dmem_n19342), .ZN(MEM_stage_inst_dmem_n19331) );
NAND2_X1 MEM_stage_inst_dmem_U18397 ( .A1(MEM_stage_inst_dmem_n19329), .A2(MEM_stage_inst_dmem_n19328), .ZN(MEM_stage_inst_dmem_n9762) );
NAND2_X1 MEM_stage_inst_dmem_U18396 ( .A1(MEM_stage_inst_dmem_n16361), .A2(MEM_stage_inst_dmem_n19343), .ZN(MEM_stage_inst_dmem_n19328) );
NAND2_X1 MEM_stage_inst_dmem_U18395 ( .A1(MEM_stage_inst_dmem_ram_3559), .A2(MEM_stage_inst_dmem_n19342), .ZN(MEM_stage_inst_dmem_n19329) );
NAND2_X1 MEM_stage_inst_dmem_U18394 ( .A1(MEM_stage_inst_dmem_n19327), .A2(MEM_stage_inst_dmem_n19326), .ZN(MEM_stage_inst_dmem_n9763) );
NAND2_X1 MEM_stage_inst_dmem_U18393 ( .A1(MEM_stage_inst_dmem_n13051), .A2(MEM_stage_inst_dmem_n19343), .ZN(MEM_stage_inst_dmem_n19326) );
NAND2_X1 MEM_stage_inst_dmem_U18392 ( .A1(MEM_stage_inst_dmem_ram_3560), .A2(MEM_stage_inst_dmem_n19342), .ZN(MEM_stage_inst_dmem_n19327) );
NAND2_X1 MEM_stage_inst_dmem_U18391 ( .A1(MEM_stage_inst_dmem_n19325), .A2(MEM_stage_inst_dmem_n19324), .ZN(MEM_stage_inst_dmem_n9764) );
NAND2_X1 MEM_stage_inst_dmem_U18390 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n19343), .ZN(MEM_stage_inst_dmem_n19324) );
NAND2_X1 MEM_stage_inst_dmem_U18389 ( .A1(MEM_stage_inst_dmem_ram_3561), .A2(MEM_stage_inst_dmem_n19342), .ZN(MEM_stage_inst_dmem_n19325) );
NAND2_X1 MEM_stage_inst_dmem_U18388 ( .A1(MEM_stage_inst_dmem_n19323), .A2(MEM_stage_inst_dmem_n19322), .ZN(MEM_stage_inst_dmem_n9765) );
NAND2_X1 MEM_stage_inst_dmem_U18387 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n19343), .ZN(MEM_stage_inst_dmem_n19322) );
NAND2_X1 MEM_stage_inst_dmem_U18386 ( .A1(MEM_stage_inst_dmem_ram_3562), .A2(MEM_stage_inst_dmem_n19342), .ZN(MEM_stage_inst_dmem_n19323) );
NAND2_X1 MEM_stage_inst_dmem_U18385 ( .A1(MEM_stage_inst_dmem_n19321), .A2(MEM_stage_inst_dmem_n19320), .ZN(MEM_stage_inst_dmem_n9766) );
NAND2_X1 MEM_stage_inst_dmem_U18384 ( .A1(EX_pipeline_reg_out_16), .A2(MEM_stage_inst_dmem_n19343), .ZN(MEM_stage_inst_dmem_n19320) );
NAND2_X1 MEM_stage_inst_dmem_U18383 ( .A1(MEM_stage_inst_dmem_ram_3563), .A2(MEM_stage_inst_dmem_n19342), .ZN(MEM_stage_inst_dmem_n19321) );
NAND2_X1 MEM_stage_inst_dmem_U18382 ( .A1(MEM_stage_inst_dmem_n19319), .A2(MEM_stage_inst_dmem_n19318), .ZN(MEM_stage_inst_dmem_n9767) );
NAND2_X1 MEM_stage_inst_dmem_U18381 ( .A1(EX_pipeline_reg_out_17), .A2(MEM_stage_inst_dmem_n19343), .ZN(MEM_stage_inst_dmem_n19318) );
NAND2_X1 MEM_stage_inst_dmem_U18380 ( .A1(MEM_stage_inst_dmem_ram_3564), .A2(MEM_stage_inst_dmem_n19342), .ZN(MEM_stage_inst_dmem_n19319) );
NAND2_X1 MEM_stage_inst_dmem_U18379 ( .A1(MEM_stage_inst_dmem_n19317), .A2(MEM_stage_inst_dmem_n19316), .ZN(MEM_stage_inst_dmem_n9768) );
NAND2_X1 MEM_stage_inst_dmem_U18378 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n19343), .ZN(MEM_stage_inst_dmem_n19316) );
NAND2_X1 MEM_stage_inst_dmem_U18377 ( .A1(MEM_stage_inst_dmem_ram_3565), .A2(MEM_stage_inst_dmem_n19342), .ZN(MEM_stage_inst_dmem_n19317) );
NAND2_X1 MEM_stage_inst_dmem_U18376 ( .A1(MEM_stage_inst_dmem_n19315), .A2(MEM_stage_inst_dmem_n19314), .ZN(MEM_stage_inst_dmem_n9769) );
NAND2_X1 MEM_stage_inst_dmem_U18375 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n19343), .ZN(MEM_stage_inst_dmem_n19314) );
NAND2_X1 MEM_stage_inst_dmem_U18374 ( .A1(MEM_stage_inst_dmem_ram_3566), .A2(MEM_stage_inst_dmem_n19342), .ZN(MEM_stage_inst_dmem_n19315) );
NAND2_X1 MEM_stage_inst_dmem_U18373 ( .A1(MEM_stage_inst_dmem_n19313), .A2(MEM_stage_inst_dmem_n19312), .ZN(MEM_stage_inst_dmem_n9770) );
NAND2_X1 MEM_stage_inst_dmem_U18372 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n19343), .ZN(MEM_stage_inst_dmem_n19312) );
INV_X1 MEM_stage_inst_dmem_U18371 ( .A(MEM_stage_inst_dmem_n19342), .ZN(MEM_stage_inst_dmem_n19343) );
NAND2_X1 MEM_stage_inst_dmem_U18370 ( .A1(MEM_stage_inst_dmem_ram_3567), .A2(MEM_stage_inst_dmem_n19342), .ZN(MEM_stage_inst_dmem_n19313) );
NAND2_X1 MEM_stage_inst_dmem_U18369 ( .A1(MEM_stage_inst_dmem_n20969), .A2(MEM_stage_inst_dmem_n19788), .ZN(MEM_stage_inst_dmem_n19342) );
NAND2_X1 MEM_stage_inst_dmem_U18368 ( .A1(MEM_stage_inst_dmem_n19311), .A2(MEM_stage_inst_dmem_n19310), .ZN(MEM_stage_inst_dmem_n9771) );
NAND2_X1 MEM_stage_inst_dmem_U18367 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n19309), .ZN(MEM_stage_inst_dmem_n19310) );
BUF_X2 MEM_stage_inst_dmem_U18366 ( .A(MEM_stage_inst_dmem_n20551), .Z(MEM_stage_inst_dmem_n21501) );
NAND2_X1 MEM_stage_inst_dmem_U18365 ( .A1(MEM_stage_inst_dmem_ram_3568), .A2(MEM_stage_inst_dmem_n19308), .ZN(MEM_stage_inst_dmem_n19311) );
NAND2_X1 MEM_stage_inst_dmem_U18364 ( .A1(MEM_stage_inst_dmem_n19307), .A2(MEM_stage_inst_dmem_n19306), .ZN(MEM_stage_inst_dmem_n9772) );
NAND2_X1 MEM_stage_inst_dmem_U18363 ( .A1(MEM_stage_inst_dmem_n20547), .A2(MEM_stage_inst_dmem_n19309), .ZN(MEM_stage_inst_dmem_n19306) );
NAND2_X1 MEM_stage_inst_dmem_U18362 ( .A1(MEM_stage_inst_dmem_ram_3569), .A2(MEM_stage_inst_dmem_n19308), .ZN(MEM_stage_inst_dmem_n19307) );
NAND2_X1 MEM_stage_inst_dmem_U18361 ( .A1(MEM_stage_inst_dmem_n19305), .A2(MEM_stage_inst_dmem_n19304), .ZN(MEM_stage_inst_dmem_n9773) );
NAND2_X1 MEM_stage_inst_dmem_U18360 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n19309), .ZN(MEM_stage_inst_dmem_n19304) );
NAND2_X1 MEM_stage_inst_dmem_U18359 ( .A1(MEM_stage_inst_dmem_ram_3570), .A2(MEM_stage_inst_dmem_n19308), .ZN(MEM_stage_inst_dmem_n19305) );
NAND2_X1 MEM_stage_inst_dmem_U18358 ( .A1(MEM_stage_inst_dmem_n19303), .A2(MEM_stage_inst_dmem_n19302), .ZN(MEM_stage_inst_dmem_n9774) );
NAND2_X1 MEM_stage_inst_dmem_U18357 ( .A1(EX_pipeline_reg_out_8), .A2(MEM_stage_inst_dmem_n19309), .ZN(MEM_stage_inst_dmem_n19302) );
NAND2_X1 MEM_stage_inst_dmem_U18356 ( .A1(MEM_stage_inst_dmem_ram_3571), .A2(MEM_stage_inst_dmem_n19308), .ZN(MEM_stage_inst_dmem_n19303) );
NAND2_X1 MEM_stage_inst_dmem_U18355 ( .A1(MEM_stage_inst_dmem_n19301), .A2(MEM_stage_inst_dmem_n19300), .ZN(MEM_stage_inst_dmem_n9775) );
NAND2_X1 MEM_stage_inst_dmem_U18354 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n19309), .ZN(MEM_stage_inst_dmem_n19300) );
NAND2_X1 MEM_stage_inst_dmem_U18353 ( .A1(MEM_stage_inst_dmem_ram_3572), .A2(MEM_stage_inst_dmem_n19308), .ZN(MEM_stage_inst_dmem_n19301) );
NAND2_X1 MEM_stage_inst_dmem_U18352 ( .A1(MEM_stage_inst_dmem_n19299), .A2(MEM_stage_inst_dmem_n19298), .ZN(MEM_stage_inst_dmem_n9776) );
NAND2_X1 MEM_stage_inst_dmem_U18351 ( .A1(EX_pipeline_reg_out_10), .A2(MEM_stage_inst_dmem_n19309), .ZN(MEM_stage_inst_dmem_n19298) );
NAND2_X1 MEM_stage_inst_dmem_U18350 ( .A1(MEM_stage_inst_dmem_ram_3573), .A2(MEM_stage_inst_dmem_n19308), .ZN(MEM_stage_inst_dmem_n19299) );
NAND2_X1 MEM_stage_inst_dmem_U18349 ( .A1(MEM_stage_inst_dmem_n19297), .A2(MEM_stage_inst_dmem_n19296), .ZN(MEM_stage_inst_dmem_n9777) );
NAND2_X1 MEM_stage_inst_dmem_U18348 ( .A1(EX_pipeline_reg_out_11), .A2(MEM_stage_inst_dmem_n19309), .ZN(MEM_stage_inst_dmem_n19296) );
NAND2_X1 MEM_stage_inst_dmem_U18347 ( .A1(MEM_stage_inst_dmem_ram_3574), .A2(MEM_stage_inst_dmem_n19308), .ZN(MEM_stage_inst_dmem_n19297) );
NAND2_X1 MEM_stage_inst_dmem_U18346 ( .A1(MEM_stage_inst_dmem_n19295), .A2(MEM_stage_inst_dmem_n19294), .ZN(MEM_stage_inst_dmem_n9778) );
NAND2_X1 MEM_stage_inst_dmem_U18345 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n19309), .ZN(MEM_stage_inst_dmem_n19294) );
NAND2_X1 MEM_stage_inst_dmem_U18344 ( .A1(MEM_stage_inst_dmem_ram_3575), .A2(MEM_stage_inst_dmem_n19308), .ZN(MEM_stage_inst_dmem_n19295) );
NAND2_X1 MEM_stage_inst_dmem_U18343 ( .A1(MEM_stage_inst_dmem_n19293), .A2(MEM_stage_inst_dmem_n19292), .ZN(MEM_stage_inst_dmem_n9779) );
NAND2_X1 MEM_stage_inst_dmem_U18342 ( .A1(MEM_stage_inst_dmem_n13051), .A2(MEM_stage_inst_dmem_n19309), .ZN(MEM_stage_inst_dmem_n19292) );
NAND2_X1 MEM_stage_inst_dmem_U18341 ( .A1(MEM_stage_inst_dmem_ram_3576), .A2(MEM_stage_inst_dmem_n19308), .ZN(MEM_stage_inst_dmem_n19293) );
NAND2_X1 MEM_stage_inst_dmem_U18340 ( .A1(MEM_stage_inst_dmem_n19291), .A2(MEM_stage_inst_dmem_n19290), .ZN(MEM_stage_inst_dmem_n9780) );
NAND2_X1 MEM_stage_inst_dmem_U18339 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n19309), .ZN(MEM_stage_inst_dmem_n19290) );
NAND2_X1 MEM_stage_inst_dmem_U18338 ( .A1(MEM_stage_inst_dmem_ram_3577), .A2(MEM_stage_inst_dmem_n19308), .ZN(MEM_stage_inst_dmem_n19291) );
NAND2_X1 MEM_stage_inst_dmem_U18337 ( .A1(MEM_stage_inst_dmem_n19289), .A2(MEM_stage_inst_dmem_n19288), .ZN(MEM_stage_inst_dmem_n9781) );
NAND2_X1 MEM_stage_inst_dmem_U18336 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n19309), .ZN(MEM_stage_inst_dmem_n19288) );
NAND2_X1 MEM_stage_inst_dmem_U18335 ( .A1(MEM_stage_inst_dmem_ram_3578), .A2(MEM_stage_inst_dmem_n19308), .ZN(MEM_stage_inst_dmem_n19289) );
NAND2_X1 MEM_stage_inst_dmem_U18334 ( .A1(MEM_stage_inst_dmem_n19287), .A2(MEM_stage_inst_dmem_n19286), .ZN(MEM_stage_inst_dmem_n9782) );
NAND2_X1 MEM_stage_inst_dmem_U18333 ( .A1(MEM_stage_inst_dmem_n14705), .A2(MEM_stage_inst_dmem_n19309), .ZN(MEM_stage_inst_dmem_n19286) );
NAND2_X1 MEM_stage_inst_dmem_U18332 ( .A1(MEM_stage_inst_dmem_ram_3579), .A2(MEM_stage_inst_dmem_n19308), .ZN(MEM_stage_inst_dmem_n19287) );
NAND2_X1 MEM_stage_inst_dmem_U18331 ( .A1(MEM_stage_inst_dmem_n19285), .A2(MEM_stage_inst_dmem_n19284), .ZN(MEM_stage_inst_dmem_n9783) );
NAND2_X1 MEM_stage_inst_dmem_U18330 ( .A1(MEM_stage_inst_dmem_n21474), .A2(MEM_stage_inst_dmem_n19309), .ZN(MEM_stage_inst_dmem_n19284) );
NAND2_X1 MEM_stage_inst_dmem_U18329 ( .A1(MEM_stage_inst_dmem_ram_3580), .A2(MEM_stage_inst_dmem_n19308), .ZN(MEM_stage_inst_dmem_n19285) );
NAND2_X1 MEM_stage_inst_dmem_U18328 ( .A1(MEM_stage_inst_dmem_n19283), .A2(MEM_stage_inst_dmem_n19282), .ZN(MEM_stage_inst_dmem_n9784) );
NAND2_X1 MEM_stage_inst_dmem_U18327 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n19309), .ZN(MEM_stage_inst_dmem_n19282) );
BUF_X2 MEM_stage_inst_dmem_U18326 ( .A(MEM_stage_inst_dmem_n20512), .Z(MEM_stage_inst_dmem_n21471) );
NAND2_X1 MEM_stage_inst_dmem_U18325 ( .A1(MEM_stage_inst_dmem_ram_3581), .A2(MEM_stage_inst_dmem_n19308), .ZN(MEM_stage_inst_dmem_n19283) );
NAND2_X1 MEM_stage_inst_dmem_U18324 ( .A1(MEM_stage_inst_dmem_n19281), .A2(MEM_stage_inst_dmem_n19280), .ZN(MEM_stage_inst_dmem_n9785) );
NAND2_X1 MEM_stage_inst_dmem_U18323 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n19309), .ZN(MEM_stage_inst_dmem_n19280) );
BUF_X2 MEM_stage_inst_dmem_U18322 ( .A(MEM_stage_inst_dmem_n20509), .Z(MEM_stage_inst_dmem_n21468) );
NAND2_X1 MEM_stage_inst_dmem_U18321 ( .A1(MEM_stage_inst_dmem_ram_3582), .A2(MEM_stage_inst_dmem_n19308), .ZN(MEM_stage_inst_dmem_n19281) );
NAND2_X1 MEM_stage_inst_dmem_U18320 ( .A1(MEM_stage_inst_dmem_n19279), .A2(MEM_stage_inst_dmem_n19278), .ZN(MEM_stage_inst_dmem_n9786) );
NAND2_X1 MEM_stage_inst_dmem_U18319 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n19309), .ZN(MEM_stage_inst_dmem_n19278) );
INV_X1 MEM_stage_inst_dmem_U18318 ( .A(MEM_stage_inst_dmem_n19308), .ZN(MEM_stage_inst_dmem_n19309) );
NAND2_X1 MEM_stage_inst_dmem_U18317 ( .A1(MEM_stage_inst_dmem_ram_3583), .A2(MEM_stage_inst_dmem_n19308), .ZN(MEM_stage_inst_dmem_n19279) );
NAND2_X1 MEM_stage_inst_dmem_U18316 ( .A1(MEM_stage_inst_dmem_n20934), .A2(MEM_stage_inst_dmem_n19788), .ZN(MEM_stage_inst_dmem_n19308) );
NOR2_X2 MEM_stage_inst_dmem_U18315 ( .A1(MEM_stage_inst_dmem_n19823), .A2(MEM_stage_inst_dmem_n20369), .ZN(MEM_stage_inst_dmem_n19788) );
NAND2_X1 MEM_stage_inst_dmem_U18314 ( .A1(MEM_stage_inst_dmem_n19277), .A2(MEM_stage_inst_dmem_n19276), .ZN(MEM_stage_inst_dmem_n9787) );
NAND2_X1 MEM_stage_inst_dmem_U18313 ( .A1(MEM_stage_inst_dmem_n19275), .A2(MEM_stage_inst_dmem_n19274), .ZN(MEM_stage_inst_dmem_n19276) );
NAND2_X1 MEM_stage_inst_dmem_U18312 ( .A1(MEM_stage_inst_dmem_ram_2560), .A2(MEM_stage_inst_dmem_n19273), .ZN(MEM_stage_inst_dmem_n19277) );
NAND2_X1 MEM_stage_inst_dmem_U18311 ( .A1(MEM_stage_inst_dmem_n19272), .A2(MEM_stage_inst_dmem_n19271), .ZN(MEM_stage_inst_dmem_n9788) );
NAND2_X1 MEM_stage_inst_dmem_U18310 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n19274), .ZN(MEM_stage_inst_dmem_n19271) );
NAND2_X1 MEM_stage_inst_dmem_U18309 ( .A1(MEM_stage_inst_dmem_ram_2561), .A2(MEM_stage_inst_dmem_n19273), .ZN(MEM_stage_inst_dmem_n19272) );
NAND2_X1 MEM_stage_inst_dmem_U18308 ( .A1(MEM_stage_inst_dmem_n19270), .A2(MEM_stage_inst_dmem_n19269), .ZN(MEM_stage_inst_dmem_n9789) );
NAND2_X1 MEM_stage_inst_dmem_U18307 ( .A1(EX_pipeline_reg_out_7), .A2(MEM_stage_inst_dmem_n19274), .ZN(MEM_stage_inst_dmem_n19269) );
NAND2_X1 MEM_stage_inst_dmem_U18306 ( .A1(MEM_stage_inst_dmem_ram_2562), .A2(MEM_stage_inst_dmem_n19273), .ZN(MEM_stage_inst_dmem_n19270) );
NAND2_X1 MEM_stage_inst_dmem_U18305 ( .A1(MEM_stage_inst_dmem_n19268), .A2(MEM_stage_inst_dmem_n19267), .ZN(MEM_stage_inst_dmem_n9790) );
NAND2_X1 MEM_stage_inst_dmem_U18304 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n19274), .ZN(MEM_stage_inst_dmem_n19267) );
NAND2_X1 MEM_stage_inst_dmem_U18303 ( .A1(MEM_stage_inst_dmem_ram_2563), .A2(MEM_stage_inst_dmem_n19273), .ZN(MEM_stage_inst_dmem_n19268) );
NAND2_X1 MEM_stage_inst_dmem_U18302 ( .A1(MEM_stage_inst_dmem_n19265), .A2(MEM_stage_inst_dmem_n19264), .ZN(MEM_stage_inst_dmem_n9791) );
NAND2_X1 MEM_stage_inst_dmem_U18301 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n19274), .ZN(MEM_stage_inst_dmem_n19264) );
NAND2_X1 MEM_stage_inst_dmem_U18300 ( .A1(MEM_stage_inst_dmem_ram_2564), .A2(MEM_stage_inst_dmem_n19273), .ZN(MEM_stage_inst_dmem_n19265) );
NAND2_X1 MEM_stage_inst_dmem_U18299 ( .A1(MEM_stage_inst_dmem_n19262), .A2(MEM_stage_inst_dmem_n19261), .ZN(MEM_stage_inst_dmem_n9792) );
NAND2_X1 MEM_stage_inst_dmem_U18298 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n19274), .ZN(MEM_stage_inst_dmem_n19261) );
NAND2_X1 MEM_stage_inst_dmem_U18297 ( .A1(MEM_stage_inst_dmem_ram_2565), .A2(MEM_stage_inst_dmem_n19273), .ZN(MEM_stage_inst_dmem_n19262) );
NAND2_X1 MEM_stage_inst_dmem_U18296 ( .A1(MEM_stage_inst_dmem_n19259), .A2(MEM_stage_inst_dmem_n19258), .ZN(MEM_stage_inst_dmem_n9793) );
NAND2_X1 MEM_stage_inst_dmem_U18295 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n19274), .ZN(MEM_stage_inst_dmem_n19258) );
NAND2_X1 MEM_stage_inst_dmem_U18294 ( .A1(MEM_stage_inst_dmem_ram_2566), .A2(MEM_stage_inst_dmem_n19273), .ZN(MEM_stage_inst_dmem_n19259) );
NAND2_X1 MEM_stage_inst_dmem_U18293 ( .A1(MEM_stage_inst_dmem_n19257), .A2(MEM_stage_inst_dmem_n19256), .ZN(MEM_stage_inst_dmem_n9794) );
NAND2_X1 MEM_stage_inst_dmem_U18292 ( .A1(MEM_stage_inst_dmem_n18875), .A2(MEM_stage_inst_dmem_n19274), .ZN(MEM_stage_inst_dmem_n19256) );
NAND2_X1 MEM_stage_inst_dmem_U18291 ( .A1(MEM_stage_inst_dmem_ram_2567), .A2(MEM_stage_inst_dmem_n19273), .ZN(MEM_stage_inst_dmem_n19257) );
NAND2_X1 MEM_stage_inst_dmem_U18290 ( .A1(MEM_stage_inst_dmem_n19255), .A2(MEM_stage_inst_dmem_n19254), .ZN(MEM_stage_inst_dmem_n9795) );
NAND2_X1 MEM_stage_inst_dmem_U18289 ( .A1(EX_pipeline_reg_out_13), .A2(MEM_stage_inst_dmem_n19274), .ZN(MEM_stage_inst_dmem_n19254) );
NAND2_X1 MEM_stage_inst_dmem_U18288 ( .A1(MEM_stage_inst_dmem_ram_2568), .A2(MEM_stage_inst_dmem_n19273), .ZN(MEM_stage_inst_dmem_n19255) );
NAND2_X1 MEM_stage_inst_dmem_U18287 ( .A1(MEM_stage_inst_dmem_n19253), .A2(MEM_stage_inst_dmem_n19252), .ZN(MEM_stage_inst_dmem_n9796) );
NAND2_X1 MEM_stage_inst_dmem_U18286 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n19274), .ZN(MEM_stage_inst_dmem_n19252) );
NAND2_X1 MEM_stage_inst_dmem_U18285 ( .A1(MEM_stage_inst_dmem_ram_2569), .A2(MEM_stage_inst_dmem_n19273), .ZN(MEM_stage_inst_dmem_n19253) );
NAND2_X1 MEM_stage_inst_dmem_U18284 ( .A1(MEM_stage_inst_dmem_n19250), .A2(MEM_stage_inst_dmem_n19249), .ZN(MEM_stage_inst_dmem_n9797) );
NAND2_X1 MEM_stage_inst_dmem_U18283 ( .A1(EX_pipeline_reg_out_15), .A2(MEM_stage_inst_dmem_n19274), .ZN(MEM_stage_inst_dmem_n19249) );
NAND2_X1 MEM_stage_inst_dmem_U18282 ( .A1(MEM_stage_inst_dmem_ram_2570), .A2(MEM_stage_inst_dmem_n19273), .ZN(MEM_stage_inst_dmem_n19250) );
NAND2_X1 MEM_stage_inst_dmem_U18281 ( .A1(MEM_stage_inst_dmem_n19248), .A2(MEM_stage_inst_dmem_n19247), .ZN(MEM_stage_inst_dmem_n9798) );
NAND2_X1 MEM_stage_inst_dmem_U18280 ( .A1(MEM_stage_inst_dmem_n20904), .A2(MEM_stage_inst_dmem_n19274), .ZN(MEM_stage_inst_dmem_n19247) );
NAND2_X1 MEM_stage_inst_dmem_U18279 ( .A1(MEM_stage_inst_dmem_ram_2571), .A2(MEM_stage_inst_dmem_n19273), .ZN(MEM_stage_inst_dmem_n19248) );
NAND2_X1 MEM_stage_inst_dmem_U18278 ( .A1(MEM_stage_inst_dmem_n19246), .A2(MEM_stage_inst_dmem_n19245), .ZN(MEM_stage_inst_dmem_n9799) );
NAND2_X1 MEM_stage_inst_dmem_U18277 ( .A1(MEM_stage_inst_dmem_n21474), .A2(MEM_stage_inst_dmem_n19274), .ZN(MEM_stage_inst_dmem_n19245) );
NAND2_X1 MEM_stage_inst_dmem_U18276 ( .A1(MEM_stage_inst_dmem_ram_2572), .A2(MEM_stage_inst_dmem_n19273), .ZN(MEM_stage_inst_dmem_n19246) );
NAND2_X1 MEM_stage_inst_dmem_U18275 ( .A1(MEM_stage_inst_dmem_n19244), .A2(MEM_stage_inst_dmem_n19243), .ZN(MEM_stage_inst_dmem_n9800) );
NAND2_X1 MEM_stage_inst_dmem_U18274 ( .A1(MEM_stage_inst_dmem_n19242), .A2(MEM_stage_inst_dmem_n19274), .ZN(MEM_stage_inst_dmem_n19243) );
NAND2_X1 MEM_stage_inst_dmem_U18273 ( .A1(MEM_stage_inst_dmem_ram_2573), .A2(MEM_stage_inst_dmem_n19273), .ZN(MEM_stage_inst_dmem_n19244) );
NAND2_X1 MEM_stage_inst_dmem_U18272 ( .A1(MEM_stage_inst_dmem_n19241), .A2(MEM_stage_inst_dmem_n19240), .ZN(MEM_stage_inst_dmem_n9801) );
NAND2_X1 MEM_stage_inst_dmem_U18271 ( .A1(MEM_stage_inst_dmem_n115), .A2(MEM_stage_inst_dmem_n19274), .ZN(MEM_stage_inst_dmem_n19240) );
NAND2_X1 MEM_stage_inst_dmem_U18270 ( .A1(MEM_stage_inst_dmem_ram_2574), .A2(MEM_stage_inst_dmem_n19273), .ZN(MEM_stage_inst_dmem_n19241) );
NAND2_X1 MEM_stage_inst_dmem_U18269 ( .A1(MEM_stage_inst_dmem_n19238), .A2(MEM_stage_inst_dmem_n19237), .ZN(MEM_stage_inst_dmem_n9802) );
NAND2_X1 MEM_stage_inst_dmem_U18268 ( .A1(EX_pipeline_reg_out_20), .A2(MEM_stage_inst_dmem_n19274), .ZN(MEM_stage_inst_dmem_n19237) );
INV_X1 MEM_stage_inst_dmem_U18267 ( .A(MEM_stage_inst_dmem_n19273), .ZN(MEM_stage_inst_dmem_n19274) );
NAND2_X1 MEM_stage_inst_dmem_U18266 ( .A1(MEM_stage_inst_dmem_ram_2575), .A2(MEM_stage_inst_dmem_n19273), .ZN(MEM_stage_inst_dmem_n19238) );
NAND2_X1 MEM_stage_inst_dmem_U18265 ( .A1(MEM_stage_inst_dmem_n21465), .A2(MEM_stage_inst_dmem_n19236), .ZN(MEM_stage_inst_dmem_n19273) );
NAND2_X1 MEM_stage_inst_dmem_U18264 ( .A1(MEM_stage_inst_dmem_n19235), .A2(MEM_stage_inst_dmem_n19234), .ZN(MEM_stage_inst_dmem_n9803) );
NAND2_X1 MEM_stage_inst_dmem_U18263 ( .A1(MEM_stage_inst_dmem_n19275), .A2(MEM_stage_inst_dmem_n19233), .ZN(MEM_stage_inst_dmem_n19234) );
NAND2_X1 MEM_stage_inst_dmem_U18262 ( .A1(MEM_stage_inst_dmem_ram_2576), .A2(MEM_stage_inst_dmem_n19232), .ZN(MEM_stage_inst_dmem_n19235) );
NAND2_X1 MEM_stage_inst_dmem_U18261 ( .A1(MEM_stage_inst_dmem_n19231), .A2(MEM_stage_inst_dmem_n19230), .ZN(MEM_stage_inst_dmem_n9804) );
NAND2_X1 MEM_stage_inst_dmem_U18260 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n19233), .ZN(MEM_stage_inst_dmem_n19230) );
NAND2_X1 MEM_stage_inst_dmem_U18259 ( .A1(MEM_stage_inst_dmem_ram_2577), .A2(MEM_stage_inst_dmem_n19232), .ZN(MEM_stage_inst_dmem_n19231) );
NAND2_X1 MEM_stage_inst_dmem_U18258 ( .A1(MEM_stage_inst_dmem_n19229), .A2(MEM_stage_inst_dmem_n19228), .ZN(MEM_stage_inst_dmem_n9805) );
NAND2_X1 MEM_stage_inst_dmem_U18257 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n19233), .ZN(MEM_stage_inst_dmem_n19228) );
NAND2_X1 MEM_stage_inst_dmem_U18256 ( .A1(MEM_stage_inst_dmem_ram_2578), .A2(MEM_stage_inst_dmem_n19232), .ZN(MEM_stage_inst_dmem_n19229) );
NAND2_X1 MEM_stage_inst_dmem_U18255 ( .A1(MEM_stage_inst_dmem_n19227), .A2(MEM_stage_inst_dmem_n19226), .ZN(MEM_stage_inst_dmem_n9806) );
NAND2_X1 MEM_stage_inst_dmem_U18254 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n19233), .ZN(MEM_stage_inst_dmem_n19226) );
NAND2_X1 MEM_stage_inst_dmem_U18253 ( .A1(MEM_stage_inst_dmem_ram_2579), .A2(MEM_stage_inst_dmem_n19232), .ZN(MEM_stage_inst_dmem_n19227) );
NAND2_X1 MEM_stage_inst_dmem_U18252 ( .A1(MEM_stage_inst_dmem_n19225), .A2(MEM_stage_inst_dmem_n19224), .ZN(MEM_stage_inst_dmem_n9807) );
NAND2_X1 MEM_stage_inst_dmem_U18251 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n19233), .ZN(MEM_stage_inst_dmem_n19224) );
NAND2_X1 MEM_stage_inst_dmem_U18250 ( .A1(MEM_stage_inst_dmem_ram_2580), .A2(MEM_stage_inst_dmem_n19232), .ZN(MEM_stage_inst_dmem_n19225) );
NAND2_X1 MEM_stage_inst_dmem_U18249 ( .A1(MEM_stage_inst_dmem_n19223), .A2(MEM_stage_inst_dmem_n19222), .ZN(MEM_stage_inst_dmem_n9808) );
NAND2_X1 MEM_stage_inst_dmem_U18248 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n19233), .ZN(MEM_stage_inst_dmem_n19222) );
NAND2_X1 MEM_stage_inst_dmem_U18247 ( .A1(MEM_stage_inst_dmem_ram_2581), .A2(MEM_stage_inst_dmem_n19232), .ZN(MEM_stage_inst_dmem_n19223) );
NAND2_X1 MEM_stage_inst_dmem_U18246 ( .A1(MEM_stage_inst_dmem_n19221), .A2(MEM_stage_inst_dmem_n19220), .ZN(MEM_stage_inst_dmem_n9809) );
NAND2_X1 MEM_stage_inst_dmem_U18245 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n19233), .ZN(MEM_stage_inst_dmem_n19220) );
NAND2_X1 MEM_stage_inst_dmem_U18244 ( .A1(MEM_stage_inst_dmem_ram_2582), .A2(MEM_stage_inst_dmem_n19232), .ZN(MEM_stage_inst_dmem_n19221) );
NAND2_X1 MEM_stage_inst_dmem_U18243 ( .A1(MEM_stage_inst_dmem_n19219), .A2(MEM_stage_inst_dmem_n19218), .ZN(MEM_stage_inst_dmem_n9810) );
NAND2_X1 MEM_stage_inst_dmem_U18242 ( .A1(MEM_stage_inst_dmem_n20530), .A2(MEM_stage_inst_dmem_n19233), .ZN(MEM_stage_inst_dmem_n19218) );
NAND2_X1 MEM_stage_inst_dmem_U18241 ( .A1(MEM_stage_inst_dmem_ram_2583), .A2(MEM_stage_inst_dmem_n19232), .ZN(MEM_stage_inst_dmem_n19219) );
NAND2_X1 MEM_stage_inst_dmem_U18240 ( .A1(MEM_stage_inst_dmem_n19217), .A2(MEM_stage_inst_dmem_n19216), .ZN(MEM_stage_inst_dmem_n9811) );
NAND2_X1 MEM_stage_inst_dmem_U18239 ( .A1(MEM_stage_inst_dmem_n20527), .A2(MEM_stage_inst_dmem_n19233), .ZN(MEM_stage_inst_dmem_n19216) );
NAND2_X1 MEM_stage_inst_dmem_U18238 ( .A1(MEM_stage_inst_dmem_ram_2584), .A2(MEM_stage_inst_dmem_n19232), .ZN(MEM_stage_inst_dmem_n19217) );
NAND2_X1 MEM_stage_inst_dmem_U18237 ( .A1(MEM_stage_inst_dmem_n19215), .A2(MEM_stage_inst_dmem_n19214), .ZN(MEM_stage_inst_dmem_n9812) );
NAND2_X1 MEM_stage_inst_dmem_U18236 ( .A1(MEM_stage_inst_dmem_n19251), .A2(MEM_stage_inst_dmem_n19233), .ZN(MEM_stage_inst_dmem_n19214) );
NAND2_X1 MEM_stage_inst_dmem_U18235 ( .A1(MEM_stage_inst_dmem_ram_2585), .A2(MEM_stage_inst_dmem_n19232), .ZN(MEM_stage_inst_dmem_n19215) );
NAND2_X1 MEM_stage_inst_dmem_U18234 ( .A1(MEM_stage_inst_dmem_n19213), .A2(MEM_stage_inst_dmem_n19212), .ZN(MEM_stage_inst_dmem_n9813) );
NAND2_X1 MEM_stage_inst_dmem_U18233 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n19233), .ZN(MEM_stage_inst_dmem_n19212) );
NAND2_X1 MEM_stage_inst_dmem_U18232 ( .A1(MEM_stage_inst_dmem_ram_2586), .A2(MEM_stage_inst_dmem_n19232), .ZN(MEM_stage_inst_dmem_n19213) );
NAND2_X1 MEM_stage_inst_dmem_U18231 ( .A1(MEM_stage_inst_dmem_n19211), .A2(MEM_stage_inst_dmem_n19210), .ZN(MEM_stage_inst_dmem_n9814) );
NAND2_X1 MEM_stage_inst_dmem_U18230 ( .A1(MEM_stage_inst_dmem_n14705), .A2(MEM_stage_inst_dmem_n19233), .ZN(MEM_stage_inst_dmem_n19210) );
NAND2_X1 MEM_stage_inst_dmem_U18229 ( .A1(MEM_stage_inst_dmem_ram_2587), .A2(MEM_stage_inst_dmem_n19232), .ZN(MEM_stage_inst_dmem_n19211) );
NAND2_X1 MEM_stage_inst_dmem_U18228 ( .A1(MEM_stage_inst_dmem_n19209), .A2(MEM_stage_inst_dmem_n19208), .ZN(MEM_stage_inst_dmem_n9815) );
NAND2_X1 MEM_stage_inst_dmem_U18227 ( .A1(MEM_stage_inst_dmem_n14702), .A2(MEM_stage_inst_dmem_n19233), .ZN(MEM_stage_inst_dmem_n19208) );
NAND2_X1 MEM_stage_inst_dmem_U18226 ( .A1(MEM_stage_inst_dmem_ram_2588), .A2(MEM_stage_inst_dmem_n19232), .ZN(MEM_stage_inst_dmem_n19209) );
NAND2_X1 MEM_stage_inst_dmem_U18225 ( .A1(MEM_stage_inst_dmem_n19207), .A2(MEM_stage_inst_dmem_n19206), .ZN(MEM_stage_inst_dmem_n9816) );
NAND2_X1 MEM_stage_inst_dmem_U18224 ( .A1(MEM_stage_inst_dmem_n19242), .A2(MEM_stage_inst_dmem_n19233), .ZN(MEM_stage_inst_dmem_n19206) );
NAND2_X1 MEM_stage_inst_dmem_U18223 ( .A1(MEM_stage_inst_dmem_ram_2589), .A2(MEM_stage_inst_dmem_n19232), .ZN(MEM_stage_inst_dmem_n19207) );
NAND2_X1 MEM_stage_inst_dmem_U18222 ( .A1(MEM_stage_inst_dmem_n19205), .A2(MEM_stage_inst_dmem_n19204), .ZN(MEM_stage_inst_dmem_n9817) );
NAND2_X1 MEM_stage_inst_dmem_U18221 ( .A1(MEM_stage_inst_dmem_n20509), .A2(MEM_stage_inst_dmem_n19233), .ZN(MEM_stage_inst_dmem_n19204) );
NAND2_X1 MEM_stage_inst_dmem_U18220 ( .A1(MEM_stage_inst_dmem_ram_2590), .A2(MEM_stage_inst_dmem_n19232), .ZN(MEM_stage_inst_dmem_n19205) );
NAND2_X1 MEM_stage_inst_dmem_U18219 ( .A1(MEM_stage_inst_dmem_n19203), .A2(MEM_stage_inst_dmem_n19202), .ZN(MEM_stage_inst_dmem_n9818) );
NAND2_X1 MEM_stage_inst_dmem_U18218 ( .A1(MEM_stage_inst_dmem_n20506), .A2(MEM_stage_inst_dmem_n19233), .ZN(MEM_stage_inst_dmem_n19202) );
INV_X1 MEM_stage_inst_dmem_U18217 ( .A(MEM_stage_inst_dmem_n19232), .ZN(MEM_stage_inst_dmem_n19233) );
NAND2_X1 MEM_stage_inst_dmem_U18216 ( .A1(MEM_stage_inst_dmem_ram_2591), .A2(MEM_stage_inst_dmem_n19232), .ZN(MEM_stage_inst_dmem_n19203) );
NAND2_X1 MEM_stage_inst_dmem_U18215 ( .A1(MEM_stage_inst_dmem_n21429), .A2(MEM_stage_inst_dmem_n19236), .ZN(MEM_stage_inst_dmem_n19232) );
NAND2_X1 MEM_stage_inst_dmem_U18214 ( .A1(MEM_stage_inst_dmem_n19201), .A2(MEM_stage_inst_dmem_n19200), .ZN(MEM_stage_inst_dmem_n9819) );
NAND2_X1 MEM_stage_inst_dmem_U18213 ( .A1(MEM_stage_inst_dmem_n19275), .A2(MEM_stage_inst_dmem_n19199), .ZN(MEM_stage_inst_dmem_n19200) );
NAND2_X1 MEM_stage_inst_dmem_U18212 ( .A1(MEM_stage_inst_dmem_ram_2592), .A2(MEM_stage_inst_dmem_n19198), .ZN(MEM_stage_inst_dmem_n19201) );
NAND2_X1 MEM_stage_inst_dmem_U18211 ( .A1(MEM_stage_inst_dmem_n19197), .A2(MEM_stage_inst_dmem_n19196), .ZN(MEM_stage_inst_dmem_n9820) );
NAND2_X1 MEM_stage_inst_dmem_U18210 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n19199), .ZN(MEM_stage_inst_dmem_n19196) );
NAND2_X1 MEM_stage_inst_dmem_U18209 ( .A1(MEM_stage_inst_dmem_ram_2593), .A2(MEM_stage_inst_dmem_n19198), .ZN(MEM_stage_inst_dmem_n19197) );
NAND2_X1 MEM_stage_inst_dmem_U18208 ( .A1(MEM_stage_inst_dmem_n19195), .A2(MEM_stage_inst_dmem_n19194), .ZN(MEM_stage_inst_dmem_n9821) );
NAND2_X1 MEM_stage_inst_dmem_U18207 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n19199), .ZN(MEM_stage_inst_dmem_n19194) );
NAND2_X1 MEM_stage_inst_dmem_U18206 ( .A1(MEM_stage_inst_dmem_ram_2594), .A2(MEM_stage_inst_dmem_n19198), .ZN(MEM_stage_inst_dmem_n19195) );
NAND2_X1 MEM_stage_inst_dmem_U18205 ( .A1(MEM_stage_inst_dmem_n19193), .A2(MEM_stage_inst_dmem_n19192), .ZN(MEM_stage_inst_dmem_n9822) );
NAND2_X1 MEM_stage_inst_dmem_U18204 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n19199), .ZN(MEM_stage_inst_dmem_n19192) );
NAND2_X1 MEM_stage_inst_dmem_U18203 ( .A1(MEM_stage_inst_dmem_ram_2595), .A2(MEM_stage_inst_dmem_n19198), .ZN(MEM_stage_inst_dmem_n19193) );
NAND2_X1 MEM_stage_inst_dmem_U18202 ( .A1(MEM_stage_inst_dmem_n19191), .A2(MEM_stage_inst_dmem_n19190), .ZN(MEM_stage_inst_dmem_n9823) );
NAND2_X1 MEM_stage_inst_dmem_U18201 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n19199), .ZN(MEM_stage_inst_dmem_n19190) );
NAND2_X1 MEM_stage_inst_dmem_U18200 ( .A1(MEM_stage_inst_dmem_ram_2596), .A2(MEM_stage_inst_dmem_n19198), .ZN(MEM_stage_inst_dmem_n19191) );
NAND2_X1 MEM_stage_inst_dmem_U18199 ( .A1(MEM_stage_inst_dmem_n19189), .A2(MEM_stage_inst_dmem_n19188), .ZN(MEM_stage_inst_dmem_n9824) );
NAND2_X1 MEM_stage_inst_dmem_U18198 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n19199), .ZN(MEM_stage_inst_dmem_n19188) );
NAND2_X1 MEM_stage_inst_dmem_U18197 ( .A1(MEM_stage_inst_dmem_ram_2597), .A2(MEM_stage_inst_dmem_n19198), .ZN(MEM_stage_inst_dmem_n19189) );
NAND2_X1 MEM_stage_inst_dmem_U18196 ( .A1(MEM_stage_inst_dmem_n19187), .A2(MEM_stage_inst_dmem_n19186), .ZN(MEM_stage_inst_dmem_n9825) );
NAND2_X1 MEM_stage_inst_dmem_U18195 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n19199), .ZN(MEM_stage_inst_dmem_n19186) );
NAND2_X1 MEM_stage_inst_dmem_U18194 ( .A1(MEM_stage_inst_dmem_ram_2598), .A2(MEM_stage_inst_dmem_n19198), .ZN(MEM_stage_inst_dmem_n19187) );
NAND2_X1 MEM_stage_inst_dmem_U18193 ( .A1(MEM_stage_inst_dmem_n19185), .A2(MEM_stage_inst_dmem_n19184), .ZN(MEM_stage_inst_dmem_n9826) );
NAND2_X1 MEM_stage_inst_dmem_U18192 ( .A1(EX_pipeline_reg_out_12), .A2(MEM_stage_inst_dmem_n19199), .ZN(MEM_stage_inst_dmem_n19184) );
NAND2_X1 MEM_stage_inst_dmem_U18191 ( .A1(MEM_stage_inst_dmem_ram_2599), .A2(MEM_stage_inst_dmem_n19198), .ZN(MEM_stage_inst_dmem_n19185) );
NAND2_X1 MEM_stage_inst_dmem_U18190 ( .A1(MEM_stage_inst_dmem_n19183), .A2(MEM_stage_inst_dmem_n19182), .ZN(MEM_stage_inst_dmem_n9827) );
NAND2_X1 MEM_stage_inst_dmem_U18189 ( .A1(MEM_stage_inst_dmem_n13883), .A2(MEM_stage_inst_dmem_n19199), .ZN(MEM_stage_inst_dmem_n19182) );
NAND2_X1 MEM_stage_inst_dmem_U18188 ( .A1(MEM_stage_inst_dmem_ram_2600), .A2(MEM_stage_inst_dmem_n19198), .ZN(MEM_stage_inst_dmem_n19183) );
NAND2_X1 MEM_stage_inst_dmem_U18187 ( .A1(MEM_stage_inst_dmem_n19181), .A2(MEM_stage_inst_dmem_n19180), .ZN(MEM_stage_inst_dmem_n9828) );
NAND2_X1 MEM_stage_inst_dmem_U18186 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n19199), .ZN(MEM_stage_inst_dmem_n19180) );
NAND2_X1 MEM_stage_inst_dmem_U18185 ( .A1(MEM_stage_inst_dmem_ram_2601), .A2(MEM_stage_inst_dmem_n19198), .ZN(MEM_stage_inst_dmem_n19181) );
NAND2_X1 MEM_stage_inst_dmem_U18184 ( .A1(MEM_stage_inst_dmem_n19179), .A2(MEM_stage_inst_dmem_n19178), .ZN(MEM_stage_inst_dmem_n9829) );
NAND2_X1 MEM_stage_inst_dmem_U18183 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n19199), .ZN(MEM_stage_inst_dmem_n19178) );
NAND2_X1 MEM_stage_inst_dmem_U18182 ( .A1(MEM_stage_inst_dmem_ram_2602), .A2(MEM_stage_inst_dmem_n19198), .ZN(MEM_stage_inst_dmem_n19179) );
NAND2_X1 MEM_stage_inst_dmem_U18181 ( .A1(MEM_stage_inst_dmem_n19177), .A2(MEM_stage_inst_dmem_n19176), .ZN(MEM_stage_inst_dmem_n9830) );
NAND2_X1 MEM_stage_inst_dmem_U18180 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n19199), .ZN(MEM_stage_inst_dmem_n19176) );
NAND2_X1 MEM_stage_inst_dmem_U18179 ( .A1(MEM_stage_inst_dmem_ram_2603), .A2(MEM_stage_inst_dmem_n19198), .ZN(MEM_stage_inst_dmem_n19177) );
NAND2_X1 MEM_stage_inst_dmem_U18178 ( .A1(MEM_stage_inst_dmem_n19175), .A2(MEM_stage_inst_dmem_n19174), .ZN(MEM_stage_inst_dmem_n9831) );
NAND2_X1 MEM_stage_inst_dmem_U18177 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n19199), .ZN(MEM_stage_inst_dmem_n19174) );
NAND2_X1 MEM_stage_inst_dmem_U18176 ( .A1(MEM_stage_inst_dmem_ram_2604), .A2(MEM_stage_inst_dmem_n19198), .ZN(MEM_stage_inst_dmem_n19175) );
NAND2_X1 MEM_stage_inst_dmem_U18175 ( .A1(MEM_stage_inst_dmem_n19173), .A2(MEM_stage_inst_dmem_n19172), .ZN(MEM_stage_inst_dmem_n9832) );
NAND2_X1 MEM_stage_inst_dmem_U18174 ( .A1(MEM_stage_inst_dmem_n19242), .A2(MEM_stage_inst_dmem_n19199), .ZN(MEM_stage_inst_dmem_n19172) );
NAND2_X1 MEM_stage_inst_dmem_U18173 ( .A1(MEM_stage_inst_dmem_ram_2605), .A2(MEM_stage_inst_dmem_n19198), .ZN(MEM_stage_inst_dmem_n19173) );
NAND2_X1 MEM_stage_inst_dmem_U18172 ( .A1(MEM_stage_inst_dmem_n19171), .A2(MEM_stage_inst_dmem_n19170), .ZN(MEM_stage_inst_dmem_n9833) );
NAND2_X1 MEM_stage_inst_dmem_U18171 ( .A1(MEM_stage_inst_dmem_n115), .A2(MEM_stage_inst_dmem_n19199), .ZN(MEM_stage_inst_dmem_n19170) );
NAND2_X1 MEM_stage_inst_dmem_U18170 ( .A1(MEM_stage_inst_dmem_ram_2606), .A2(MEM_stage_inst_dmem_n19198), .ZN(MEM_stage_inst_dmem_n19171) );
NAND2_X1 MEM_stage_inst_dmem_U18169 ( .A1(MEM_stage_inst_dmem_n19169), .A2(MEM_stage_inst_dmem_n19168), .ZN(MEM_stage_inst_dmem_n9834) );
NAND2_X1 MEM_stage_inst_dmem_U18168 ( .A1(MEM_stage_inst_dmem_n15110), .A2(MEM_stage_inst_dmem_n19199), .ZN(MEM_stage_inst_dmem_n19168) );
INV_X1 MEM_stage_inst_dmem_U18167 ( .A(MEM_stage_inst_dmem_n19198), .ZN(MEM_stage_inst_dmem_n19199) );
NAND2_X1 MEM_stage_inst_dmem_U18166 ( .A1(MEM_stage_inst_dmem_ram_2607), .A2(MEM_stage_inst_dmem_n19198), .ZN(MEM_stage_inst_dmem_n19169) );
NAND2_X1 MEM_stage_inst_dmem_U18165 ( .A1(MEM_stage_inst_dmem_n21394), .A2(MEM_stage_inst_dmem_n19236), .ZN(MEM_stage_inst_dmem_n19198) );
NAND2_X1 MEM_stage_inst_dmem_U18164 ( .A1(MEM_stage_inst_dmem_n19167), .A2(MEM_stage_inst_dmem_n19166), .ZN(MEM_stage_inst_dmem_n9835) );
NAND2_X1 MEM_stage_inst_dmem_U18163 ( .A1(MEM_stage_inst_dmem_n19275), .A2(MEM_stage_inst_dmem_n19165), .ZN(MEM_stage_inst_dmem_n19166) );
NAND2_X1 MEM_stage_inst_dmem_U18162 ( .A1(MEM_stage_inst_dmem_ram_2608), .A2(MEM_stage_inst_dmem_n19164), .ZN(MEM_stage_inst_dmem_n19167) );
NAND2_X1 MEM_stage_inst_dmem_U18161 ( .A1(MEM_stage_inst_dmem_n19163), .A2(MEM_stage_inst_dmem_n19162), .ZN(MEM_stage_inst_dmem_n9836) );
NAND2_X1 MEM_stage_inst_dmem_U18160 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n19165), .ZN(MEM_stage_inst_dmem_n19162) );
NAND2_X1 MEM_stage_inst_dmem_U18159 ( .A1(MEM_stage_inst_dmem_ram_2609), .A2(MEM_stage_inst_dmem_n19164), .ZN(MEM_stage_inst_dmem_n19163) );
NAND2_X1 MEM_stage_inst_dmem_U18158 ( .A1(MEM_stage_inst_dmem_n19161), .A2(MEM_stage_inst_dmem_n19160), .ZN(MEM_stage_inst_dmem_n9837) );
NAND2_X1 MEM_stage_inst_dmem_U18157 ( .A1(MEM_stage_inst_dmem_n20544), .A2(MEM_stage_inst_dmem_n19165), .ZN(MEM_stage_inst_dmem_n19160) );
NAND2_X1 MEM_stage_inst_dmem_U18156 ( .A1(MEM_stage_inst_dmem_ram_2610), .A2(MEM_stage_inst_dmem_n19164), .ZN(MEM_stage_inst_dmem_n19161) );
NAND2_X1 MEM_stage_inst_dmem_U18155 ( .A1(MEM_stage_inst_dmem_n19159), .A2(MEM_stage_inst_dmem_n19158), .ZN(MEM_stage_inst_dmem_n9838) );
NAND2_X1 MEM_stage_inst_dmem_U18154 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n19165), .ZN(MEM_stage_inst_dmem_n19158) );
NAND2_X1 MEM_stage_inst_dmem_U18153 ( .A1(MEM_stage_inst_dmem_ram_2611), .A2(MEM_stage_inst_dmem_n19164), .ZN(MEM_stage_inst_dmem_n19159) );
NAND2_X1 MEM_stage_inst_dmem_U18152 ( .A1(MEM_stage_inst_dmem_n19157), .A2(MEM_stage_inst_dmem_n19156), .ZN(MEM_stage_inst_dmem_n9839) );
NAND2_X1 MEM_stage_inst_dmem_U18151 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n19165), .ZN(MEM_stage_inst_dmem_n19156) );
NAND2_X1 MEM_stage_inst_dmem_U18150 ( .A1(MEM_stage_inst_dmem_ram_2612), .A2(MEM_stage_inst_dmem_n19164), .ZN(MEM_stage_inst_dmem_n19157) );
NAND2_X1 MEM_stage_inst_dmem_U18149 ( .A1(MEM_stage_inst_dmem_n19155), .A2(MEM_stage_inst_dmem_n19154), .ZN(MEM_stage_inst_dmem_n9840) );
NAND2_X1 MEM_stage_inst_dmem_U18148 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n19165), .ZN(MEM_stage_inst_dmem_n19154) );
NAND2_X1 MEM_stage_inst_dmem_U18147 ( .A1(MEM_stage_inst_dmem_ram_2613), .A2(MEM_stage_inst_dmem_n19164), .ZN(MEM_stage_inst_dmem_n19155) );
NAND2_X1 MEM_stage_inst_dmem_U18146 ( .A1(MEM_stage_inst_dmem_n19153), .A2(MEM_stage_inst_dmem_n19152), .ZN(MEM_stage_inst_dmem_n9841) );
NAND2_X1 MEM_stage_inst_dmem_U18145 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n19165), .ZN(MEM_stage_inst_dmem_n19152) );
NAND2_X1 MEM_stage_inst_dmem_U18144 ( .A1(MEM_stage_inst_dmem_ram_2614), .A2(MEM_stage_inst_dmem_n19164), .ZN(MEM_stage_inst_dmem_n19153) );
NAND2_X1 MEM_stage_inst_dmem_U18143 ( .A1(MEM_stage_inst_dmem_n19151), .A2(MEM_stage_inst_dmem_n19150), .ZN(MEM_stage_inst_dmem_n9842) );
NAND2_X1 MEM_stage_inst_dmem_U18142 ( .A1(MEM_stage_inst_dmem_n16361), .A2(MEM_stage_inst_dmem_n19165), .ZN(MEM_stage_inst_dmem_n19150) );
NAND2_X1 MEM_stage_inst_dmem_U18141 ( .A1(MEM_stage_inst_dmem_ram_2615), .A2(MEM_stage_inst_dmem_n19164), .ZN(MEM_stage_inst_dmem_n19151) );
NAND2_X1 MEM_stage_inst_dmem_U18140 ( .A1(MEM_stage_inst_dmem_n19149), .A2(MEM_stage_inst_dmem_n19148), .ZN(MEM_stage_inst_dmem_n9843) );
NAND2_X1 MEM_stage_inst_dmem_U18139 ( .A1(MEM_stage_inst_dmem_n20527), .A2(MEM_stage_inst_dmem_n19165), .ZN(MEM_stage_inst_dmem_n19148) );
NAND2_X1 MEM_stage_inst_dmem_U18138 ( .A1(MEM_stage_inst_dmem_ram_2616), .A2(MEM_stage_inst_dmem_n19164), .ZN(MEM_stage_inst_dmem_n19149) );
NAND2_X1 MEM_stage_inst_dmem_U18137 ( .A1(MEM_stage_inst_dmem_n19147), .A2(MEM_stage_inst_dmem_n19146), .ZN(MEM_stage_inst_dmem_n9844) );
NAND2_X1 MEM_stage_inst_dmem_U18136 ( .A1(MEM_stage_inst_dmem_n19251), .A2(MEM_stage_inst_dmem_n19165), .ZN(MEM_stage_inst_dmem_n19146) );
NAND2_X1 MEM_stage_inst_dmem_U18135 ( .A1(MEM_stage_inst_dmem_ram_2617), .A2(MEM_stage_inst_dmem_n19164), .ZN(MEM_stage_inst_dmem_n19147) );
NAND2_X1 MEM_stage_inst_dmem_U18134 ( .A1(MEM_stage_inst_dmem_n19145), .A2(MEM_stage_inst_dmem_n19144), .ZN(MEM_stage_inst_dmem_n9845) );
NAND2_X1 MEM_stage_inst_dmem_U18133 ( .A1(MEM_stage_inst_dmem_n20521), .A2(MEM_stage_inst_dmem_n19165), .ZN(MEM_stage_inst_dmem_n19144) );
NAND2_X1 MEM_stage_inst_dmem_U18132 ( .A1(MEM_stage_inst_dmem_ram_2618), .A2(MEM_stage_inst_dmem_n19164), .ZN(MEM_stage_inst_dmem_n19145) );
NAND2_X1 MEM_stage_inst_dmem_U18131 ( .A1(MEM_stage_inst_dmem_n19143), .A2(MEM_stage_inst_dmem_n19142), .ZN(MEM_stage_inst_dmem_n9846) );
NAND2_X1 MEM_stage_inst_dmem_U18130 ( .A1(MEM_stage_inst_dmem_n20904), .A2(MEM_stage_inst_dmem_n19165), .ZN(MEM_stage_inst_dmem_n19142) );
NAND2_X1 MEM_stage_inst_dmem_U18129 ( .A1(MEM_stage_inst_dmem_ram_2619), .A2(MEM_stage_inst_dmem_n19164), .ZN(MEM_stage_inst_dmem_n19143) );
NAND2_X1 MEM_stage_inst_dmem_U18128 ( .A1(MEM_stage_inst_dmem_n19141), .A2(MEM_stage_inst_dmem_n19140), .ZN(MEM_stage_inst_dmem_n9847) );
NAND2_X1 MEM_stage_inst_dmem_U18127 ( .A1(MEM_stage_inst_dmem_n21474), .A2(MEM_stage_inst_dmem_n19165), .ZN(MEM_stage_inst_dmem_n19140) );
NAND2_X1 MEM_stage_inst_dmem_U18126 ( .A1(MEM_stage_inst_dmem_ram_2620), .A2(MEM_stage_inst_dmem_n19164), .ZN(MEM_stage_inst_dmem_n19141) );
NAND2_X1 MEM_stage_inst_dmem_U18125 ( .A1(MEM_stage_inst_dmem_n19139), .A2(MEM_stage_inst_dmem_n19138), .ZN(MEM_stage_inst_dmem_n9848) );
NAND2_X1 MEM_stage_inst_dmem_U18124 ( .A1(MEM_stage_inst_dmem_n19242), .A2(MEM_stage_inst_dmem_n19165), .ZN(MEM_stage_inst_dmem_n19138) );
NAND2_X1 MEM_stage_inst_dmem_U18123 ( .A1(MEM_stage_inst_dmem_ram_2621), .A2(MEM_stage_inst_dmem_n19164), .ZN(MEM_stage_inst_dmem_n19139) );
NAND2_X1 MEM_stage_inst_dmem_U18122 ( .A1(MEM_stage_inst_dmem_n19137), .A2(MEM_stage_inst_dmem_n19136), .ZN(MEM_stage_inst_dmem_n9849) );
NAND2_X1 MEM_stage_inst_dmem_U18121 ( .A1(MEM_stage_inst_dmem_n115), .A2(MEM_stage_inst_dmem_n19165), .ZN(MEM_stage_inst_dmem_n19136) );
NAND2_X1 MEM_stage_inst_dmem_U18120 ( .A1(MEM_stage_inst_dmem_ram_2622), .A2(MEM_stage_inst_dmem_n19164), .ZN(MEM_stage_inst_dmem_n19137) );
NAND2_X1 MEM_stage_inst_dmem_U18119 ( .A1(MEM_stage_inst_dmem_n19135), .A2(MEM_stage_inst_dmem_n19134), .ZN(MEM_stage_inst_dmem_n9850) );
NAND2_X1 MEM_stage_inst_dmem_U18118 ( .A1(MEM_stage_inst_dmem_n16343), .A2(MEM_stage_inst_dmem_n19165), .ZN(MEM_stage_inst_dmem_n19134) );
INV_X1 MEM_stage_inst_dmem_U18117 ( .A(MEM_stage_inst_dmem_n19164), .ZN(MEM_stage_inst_dmem_n19165) );
NAND2_X1 MEM_stage_inst_dmem_U18116 ( .A1(MEM_stage_inst_dmem_ram_2623), .A2(MEM_stage_inst_dmem_n19164), .ZN(MEM_stage_inst_dmem_n19135) );
NAND2_X1 MEM_stage_inst_dmem_U18115 ( .A1(MEM_stage_inst_dmem_n21359), .A2(MEM_stage_inst_dmem_n19236), .ZN(MEM_stage_inst_dmem_n19164) );
NAND2_X1 MEM_stage_inst_dmem_U18114 ( .A1(MEM_stage_inst_dmem_n19133), .A2(MEM_stage_inst_dmem_n19132), .ZN(MEM_stage_inst_dmem_n9851) );
NAND2_X1 MEM_stage_inst_dmem_U18113 ( .A1(MEM_stage_inst_dmem_n19275), .A2(MEM_stage_inst_dmem_n19131), .ZN(MEM_stage_inst_dmem_n19132) );
NAND2_X1 MEM_stage_inst_dmem_U18112 ( .A1(MEM_stage_inst_dmem_ram_2624), .A2(MEM_stage_inst_dmem_n19130), .ZN(MEM_stage_inst_dmem_n19133) );
NAND2_X1 MEM_stage_inst_dmem_U18111 ( .A1(MEM_stage_inst_dmem_n19129), .A2(MEM_stage_inst_dmem_n19128), .ZN(MEM_stage_inst_dmem_n9852) );
NAND2_X1 MEM_stage_inst_dmem_U18110 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n19131), .ZN(MEM_stage_inst_dmem_n19128) );
NAND2_X1 MEM_stage_inst_dmem_U18109 ( .A1(MEM_stage_inst_dmem_ram_2625), .A2(MEM_stage_inst_dmem_n19130), .ZN(MEM_stage_inst_dmem_n19129) );
NAND2_X1 MEM_stage_inst_dmem_U18108 ( .A1(MEM_stage_inst_dmem_n19127), .A2(MEM_stage_inst_dmem_n19126), .ZN(MEM_stage_inst_dmem_n9853) );
NAND2_X1 MEM_stage_inst_dmem_U18107 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n19131), .ZN(MEM_stage_inst_dmem_n19126) );
NAND2_X1 MEM_stage_inst_dmem_U18106 ( .A1(MEM_stage_inst_dmem_ram_2626), .A2(MEM_stage_inst_dmem_n19130), .ZN(MEM_stage_inst_dmem_n19127) );
NAND2_X1 MEM_stage_inst_dmem_U18105 ( .A1(MEM_stage_inst_dmem_n19125), .A2(MEM_stage_inst_dmem_n19124), .ZN(MEM_stage_inst_dmem_n9854) );
NAND2_X1 MEM_stage_inst_dmem_U18104 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n19131), .ZN(MEM_stage_inst_dmem_n19124) );
NAND2_X1 MEM_stage_inst_dmem_U18103 ( .A1(MEM_stage_inst_dmem_ram_2627), .A2(MEM_stage_inst_dmem_n19130), .ZN(MEM_stage_inst_dmem_n19125) );
NAND2_X1 MEM_stage_inst_dmem_U18102 ( .A1(MEM_stage_inst_dmem_n19123), .A2(MEM_stage_inst_dmem_n19122), .ZN(MEM_stage_inst_dmem_n9855) );
NAND2_X1 MEM_stage_inst_dmem_U18101 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n19131), .ZN(MEM_stage_inst_dmem_n19122) );
NAND2_X1 MEM_stage_inst_dmem_U18100 ( .A1(MEM_stage_inst_dmem_ram_2628), .A2(MEM_stage_inst_dmem_n19130), .ZN(MEM_stage_inst_dmem_n19123) );
NAND2_X1 MEM_stage_inst_dmem_U18099 ( .A1(MEM_stage_inst_dmem_n19121), .A2(MEM_stage_inst_dmem_n19120), .ZN(MEM_stage_inst_dmem_n9856) );
NAND2_X1 MEM_stage_inst_dmem_U18098 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n19131), .ZN(MEM_stage_inst_dmem_n19120) );
NAND2_X1 MEM_stage_inst_dmem_U18097 ( .A1(MEM_stage_inst_dmem_ram_2629), .A2(MEM_stage_inst_dmem_n19130), .ZN(MEM_stage_inst_dmem_n19121) );
NAND2_X1 MEM_stage_inst_dmem_U18096 ( .A1(MEM_stage_inst_dmem_n19119), .A2(MEM_stage_inst_dmem_n19118), .ZN(MEM_stage_inst_dmem_n9857) );
NAND2_X1 MEM_stage_inst_dmem_U18095 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n19131), .ZN(MEM_stage_inst_dmem_n19118) );
NAND2_X1 MEM_stage_inst_dmem_U18094 ( .A1(MEM_stage_inst_dmem_ram_2630), .A2(MEM_stage_inst_dmem_n19130), .ZN(MEM_stage_inst_dmem_n19119) );
NAND2_X1 MEM_stage_inst_dmem_U18093 ( .A1(MEM_stage_inst_dmem_n19117), .A2(MEM_stage_inst_dmem_n19116), .ZN(MEM_stage_inst_dmem_n9858) );
NAND2_X1 MEM_stage_inst_dmem_U18092 ( .A1(MEM_stage_inst_dmem_n112), .A2(MEM_stage_inst_dmem_n19131), .ZN(MEM_stage_inst_dmem_n19116) );
NAND2_X1 MEM_stage_inst_dmem_U18091 ( .A1(MEM_stage_inst_dmem_ram_2631), .A2(MEM_stage_inst_dmem_n19130), .ZN(MEM_stage_inst_dmem_n19117) );
NAND2_X1 MEM_stage_inst_dmem_U18090 ( .A1(MEM_stage_inst_dmem_n19115), .A2(MEM_stage_inst_dmem_n19114), .ZN(MEM_stage_inst_dmem_n9859) );
NAND2_X1 MEM_stage_inst_dmem_U18089 ( .A1(MEM_stage_inst_dmem_n13051), .A2(MEM_stage_inst_dmem_n19131), .ZN(MEM_stage_inst_dmem_n19114) );
NAND2_X1 MEM_stage_inst_dmem_U18088 ( .A1(MEM_stage_inst_dmem_ram_2632), .A2(MEM_stage_inst_dmem_n19130), .ZN(MEM_stage_inst_dmem_n19115) );
NAND2_X1 MEM_stage_inst_dmem_U18087 ( .A1(MEM_stage_inst_dmem_n19113), .A2(MEM_stage_inst_dmem_n19112), .ZN(MEM_stage_inst_dmem_n9860) );
NAND2_X1 MEM_stage_inst_dmem_U18086 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n19131), .ZN(MEM_stage_inst_dmem_n19112) );
NAND2_X1 MEM_stage_inst_dmem_U18085 ( .A1(MEM_stage_inst_dmem_ram_2633), .A2(MEM_stage_inst_dmem_n19130), .ZN(MEM_stage_inst_dmem_n19113) );
NAND2_X1 MEM_stage_inst_dmem_U18084 ( .A1(MEM_stage_inst_dmem_n19111), .A2(MEM_stage_inst_dmem_n19110), .ZN(MEM_stage_inst_dmem_n9861) );
NAND2_X1 MEM_stage_inst_dmem_U18083 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n19131), .ZN(MEM_stage_inst_dmem_n19110) );
NAND2_X1 MEM_stage_inst_dmem_U18082 ( .A1(MEM_stage_inst_dmem_ram_2634), .A2(MEM_stage_inst_dmem_n19130), .ZN(MEM_stage_inst_dmem_n19111) );
NAND2_X1 MEM_stage_inst_dmem_U18081 ( .A1(MEM_stage_inst_dmem_n19109), .A2(MEM_stage_inst_dmem_n19108), .ZN(MEM_stage_inst_dmem_n9862) );
NAND2_X1 MEM_stage_inst_dmem_U18080 ( .A1(MEM_stage_inst_dmem_n14705), .A2(MEM_stage_inst_dmem_n19131), .ZN(MEM_stage_inst_dmem_n19108) );
NAND2_X1 MEM_stage_inst_dmem_U18079 ( .A1(MEM_stage_inst_dmem_ram_2635), .A2(MEM_stage_inst_dmem_n19130), .ZN(MEM_stage_inst_dmem_n19109) );
NAND2_X1 MEM_stage_inst_dmem_U18078 ( .A1(MEM_stage_inst_dmem_n19107), .A2(MEM_stage_inst_dmem_n19106), .ZN(MEM_stage_inst_dmem_n9863) );
NAND2_X1 MEM_stage_inst_dmem_U18077 ( .A1(MEM_stage_inst_dmem_n14702), .A2(MEM_stage_inst_dmem_n19131), .ZN(MEM_stage_inst_dmem_n19106) );
NAND2_X1 MEM_stage_inst_dmem_U18076 ( .A1(MEM_stage_inst_dmem_ram_2636), .A2(MEM_stage_inst_dmem_n19130), .ZN(MEM_stage_inst_dmem_n19107) );
NAND2_X1 MEM_stage_inst_dmem_U18075 ( .A1(MEM_stage_inst_dmem_n19105), .A2(MEM_stage_inst_dmem_n19104), .ZN(MEM_stage_inst_dmem_n9864) );
NAND2_X1 MEM_stage_inst_dmem_U18074 ( .A1(MEM_stage_inst_dmem_n19242), .A2(MEM_stage_inst_dmem_n19131), .ZN(MEM_stage_inst_dmem_n19104) );
NAND2_X1 MEM_stage_inst_dmem_U18073 ( .A1(MEM_stage_inst_dmem_ram_2637), .A2(MEM_stage_inst_dmem_n19130), .ZN(MEM_stage_inst_dmem_n19105) );
NAND2_X1 MEM_stage_inst_dmem_U18072 ( .A1(MEM_stage_inst_dmem_n19103), .A2(MEM_stage_inst_dmem_n19102), .ZN(MEM_stage_inst_dmem_n9865) );
NAND2_X1 MEM_stage_inst_dmem_U18071 ( .A1(MEM_stage_inst_dmem_n115), .A2(MEM_stage_inst_dmem_n19131), .ZN(MEM_stage_inst_dmem_n19102) );
NAND2_X1 MEM_stage_inst_dmem_U18070 ( .A1(MEM_stage_inst_dmem_ram_2638), .A2(MEM_stage_inst_dmem_n19130), .ZN(MEM_stage_inst_dmem_n19103) );
NAND2_X1 MEM_stage_inst_dmem_U18069 ( .A1(MEM_stage_inst_dmem_n19101), .A2(MEM_stage_inst_dmem_n19100), .ZN(MEM_stage_inst_dmem_n9866) );
NAND2_X1 MEM_stage_inst_dmem_U18068 ( .A1(MEM_stage_inst_dmem_n16758), .A2(MEM_stage_inst_dmem_n19131), .ZN(MEM_stage_inst_dmem_n19100) );
NAND2_X1 MEM_stage_inst_dmem_U18067 ( .A1(MEM_stage_inst_dmem_ram_2639), .A2(MEM_stage_inst_dmem_n19130), .ZN(MEM_stage_inst_dmem_n19101) );
NAND2_X1 MEM_stage_inst_dmem_U18066 ( .A1(MEM_stage_inst_dmem_n21319), .A2(MEM_stage_inst_dmem_n19236), .ZN(MEM_stage_inst_dmem_n19130) );
NAND2_X1 MEM_stage_inst_dmem_U18065 ( .A1(MEM_stage_inst_dmem_n19099), .A2(MEM_stage_inst_dmem_n19098), .ZN(MEM_stage_inst_dmem_n9867) );
NAND2_X1 MEM_stage_inst_dmem_U18064 ( .A1(MEM_stage_inst_dmem_n19275), .A2(MEM_stage_inst_dmem_n19097), .ZN(MEM_stage_inst_dmem_n19098) );
NAND2_X1 MEM_stage_inst_dmem_U18063 ( .A1(MEM_stage_inst_dmem_ram_2640), .A2(MEM_stage_inst_dmem_n19096), .ZN(MEM_stage_inst_dmem_n19099) );
NAND2_X1 MEM_stage_inst_dmem_U18062 ( .A1(MEM_stage_inst_dmem_n19095), .A2(MEM_stage_inst_dmem_n19094), .ZN(MEM_stage_inst_dmem_n9868) );
NAND2_X1 MEM_stage_inst_dmem_U18061 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n19097), .ZN(MEM_stage_inst_dmem_n19094) );
NAND2_X1 MEM_stage_inst_dmem_U18060 ( .A1(MEM_stage_inst_dmem_ram_2641), .A2(MEM_stage_inst_dmem_n19096), .ZN(MEM_stage_inst_dmem_n19095) );
NAND2_X1 MEM_stage_inst_dmem_U18059 ( .A1(MEM_stage_inst_dmem_n19093), .A2(MEM_stage_inst_dmem_n19092), .ZN(MEM_stage_inst_dmem_n9869) );
NAND2_X1 MEM_stage_inst_dmem_U18058 ( .A1(MEM_stage_inst_dmem_n16789), .A2(MEM_stage_inst_dmem_n19097), .ZN(MEM_stage_inst_dmem_n19092) );
NAND2_X1 MEM_stage_inst_dmem_U18057 ( .A1(MEM_stage_inst_dmem_ram_2642), .A2(MEM_stage_inst_dmem_n19096), .ZN(MEM_stage_inst_dmem_n19093) );
NAND2_X1 MEM_stage_inst_dmem_U18056 ( .A1(MEM_stage_inst_dmem_n19091), .A2(MEM_stage_inst_dmem_n19090), .ZN(MEM_stage_inst_dmem_n9870) );
NAND2_X1 MEM_stage_inst_dmem_U18055 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n19097), .ZN(MEM_stage_inst_dmem_n19090) );
NAND2_X1 MEM_stage_inst_dmem_U18054 ( .A1(MEM_stage_inst_dmem_ram_2643), .A2(MEM_stage_inst_dmem_n19096), .ZN(MEM_stage_inst_dmem_n19091) );
NAND2_X1 MEM_stage_inst_dmem_U18053 ( .A1(MEM_stage_inst_dmem_n19089), .A2(MEM_stage_inst_dmem_n19088), .ZN(MEM_stage_inst_dmem_n9871) );
NAND2_X1 MEM_stage_inst_dmem_U18052 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n19097), .ZN(MEM_stage_inst_dmem_n19088) );
NAND2_X1 MEM_stage_inst_dmem_U18051 ( .A1(MEM_stage_inst_dmem_ram_2644), .A2(MEM_stage_inst_dmem_n19096), .ZN(MEM_stage_inst_dmem_n19089) );
NAND2_X1 MEM_stage_inst_dmem_U18050 ( .A1(MEM_stage_inst_dmem_n19087), .A2(MEM_stage_inst_dmem_n19086), .ZN(MEM_stage_inst_dmem_n9872) );
NAND2_X1 MEM_stage_inst_dmem_U18049 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n19097), .ZN(MEM_stage_inst_dmem_n19086) );
NAND2_X1 MEM_stage_inst_dmem_U18048 ( .A1(MEM_stage_inst_dmem_ram_2645), .A2(MEM_stage_inst_dmem_n19096), .ZN(MEM_stage_inst_dmem_n19087) );
NAND2_X1 MEM_stage_inst_dmem_U18047 ( .A1(MEM_stage_inst_dmem_n19085), .A2(MEM_stage_inst_dmem_n19084), .ZN(MEM_stage_inst_dmem_n9873) );
NAND2_X1 MEM_stage_inst_dmem_U18046 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n19097), .ZN(MEM_stage_inst_dmem_n19084) );
NAND2_X1 MEM_stage_inst_dmem_U18045 ( .A1(MEM_stage_inst_dmem_ram_2646), .A2(MEM_stage_inst_dmem_n19096), .ZN(MEM_stage_inst_dmem_n19085) );
NAND2_X1 MEM_stage_inst_dmem_U18044 ( .A1(MEM_stage_inst_dmem_n19083), .A2(MEM_stage_inst_dmem_n19082), .ZN(MEM_stage_inst_dmem_n9874) );
NAND2_X1 MEM_stage_inst_dmem_U18043 ( .A1(MEM_stage_inst_dmem_n112), .A2(MEM_stage_inst_dmem_n19097), .ZN(MEM_stage_inst_dmem_n19082) );
NAND2_X1 MEM_stage_inst_dmem_U18042 ( .A1(MEM_stage_inst_dmem_ram_2647), .A2(MEM_stage_inst_dmem_n19096), .ZN(MEM_stage_inst_dmem_n19083) );
NAND2_X1 MEM_stage_inst_dmem_U18041 ( .A1(MEM_stage_inst_dmem_n19081), .A2(MEM_stage_inst_dmem_n19080), .ZN(MEM_stage_inst_dmem_n9875) );
NAND2_X1 MEM_stage_inst_dmem_U18040 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n19097), .ZN(MEM_stage_inst_dmem_n19080) );
NAND2_X1 MEM_stage_inst_dmem_U18039 ( .A1(MEM_stage_inst_dmem_ram_2648), .A2(MEM_stage_inst_dmem_n19096), .ZN(MEM_stage_inst_dmem_n19081) );
NAND2_X1 MEM_stage_inst_dmem_U18038 ( .A1(MEM_stage_inst_dmem_n19079), .A2(MEM_stage_inst_dmem_n19078), .ZN(MEM_stage_inst_dmem_n9876) );
NAND2_X1 MEM_stage_inst_dmem_U18037 ( .A1(MEM_stage_inst_dmem_n19251), .A2(MEM_stage_inst_dmem_n19097), .ZN(MEM_stage_inst_dmem_n19078) );
NAND2_X1 MEM_stage_inst_dmem_U18036 ( .A1(MEM_stage_inst_dmem_ram_2649), .A2(MEM_stage_inst_dmem_n19096), .ZN(MEM_stage_inst_dmem_n19079) );
NAND2_X1 MEM_stage_inst_dmem_U18035 ( .A1(MEM_stage_inst_dmem_n19077), .A2(MEM_stage_inst_dmem_n19076), .ZN(MEM_stage_inst_dmem_n9877) );
NAND2_X1 MEM_stage_inst_dmem_U18034 ( .A1(MEM_stage_inst_dmem_n16769), .A2(MEM_stage_inst_dmem_n19097), .ZN(MEM_stage_inst_dmem_n19076) );
NAND2_X1 MEM_stage_inst_dmem_U18033 ( .A1(MEM_stage_inst_dmem_ram_2650), .A2(MEM_stage_inst_dmem_n19096), .ZN(MEM_stage_inst_dmem_n19077) );
NAND2_X1 MEM_stage_inst_dmem_U18032 ( .A1(MEM_stage_inst_dmem_n19075), .A2(MEM_stage_inst_dmem_n19074), .ZN(MEM_stage_inst_dmem_n9878) );
NAND2_X1 MEM_stage_inst_dmem_U18031 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n19097), .ZN(MEM_stage_inst_dmem_n19074) );
NAND2_X1 MEM_stage_inst_dmem_U18030 ( .A1(MEM_stage_inst_dmem_ram_2651), .A2(MEM_stage_inst_dmem_n19096), .ZN(MEM_stage_inst_dmem_n19075) );
NAND2_X1 MEM_stage_inst_dmem_U18029 ( .A1(MEM_stage_inst_dmem_n19073), .A2(MEM_stage_inst_dmem_n19072), .ZN(MEM_stage_inst_dmem_n9879) );
NAND2_X1 MEM_stage_inst_dmem_U18028 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n19097), .ZN(MEM_stage_inst_dmem_n19072) );
NAND2_X1 MEM_stage_inst_dmem_U18027 ( .A1(MEM_stage_inst_dmem_ram_2652), .A2(MEM_stage_inst_dmem_n19096), .ZN(MEM_stage_inst_dmem_n19073) );
NAND2_X1 MEM_stage_inst_dmem_U18026 ( .A1(MEM_stage_inst_dmem_n19071), .A2(MEM_stage_inst_dmem_n19070), .ZN(MEM_stage_inst_dmem_n9880) );
NAND2_X1 MEM_stage_inst_dmem_U18025 ( .A1(MEM_stage_inst_dmem_n19242), .A2(MEM_stage_inst_dmem_n19097), .ZN(MEM_stage_inst_dmem_n19070) );
NAND2_X1 MEM_stage_inst_dmem_U18024 ( .A1(MEM_stage_inst_dmem_ram_2653), .A2(MEM_stage_inst_dmem_n19096), .ZN(MEM_stage_inst_dmem_n19071) );
NAND2_X1 MEM_stage_inst_dmem_U18023 ( .A1(MEM_stage_inst_dmem_n19069), .A2(MEM_stage_inst_dmem_n19068), .ZN(MEM_stage_inst_dmem_n9881) );
NAND2_X1 MEM_stage_inst_dmem_U18022 ( .A1(MEM_stage_inst_dmem_n115), .A2(MEM_stage_inst_dmem_n19097), .ZN(MEM_stage_inst_dmem_n19068) );
NAND2_X1 MEM_stage_inst_dmem_U18021 ( .A1(MEM_stage_inst_dmem_ram_2654), .A2(MEM_stage_inst_dmem_n19096), .ZN(MEM_stage_inst_dmem_n19069) );
NAND2_X1 MEM_stage_inst_dmem_U18020 ( .A1(MEM_stage_inst_dmem_n19067), .A2(MEM_stage_inst_dmem_n19066), .ZN(MEM_stage_inst_dmem_n9882) );
NAND2_X1 MEM_stage_inst_dmem_U18019 ( .A1(MEM_stage_inst_dmem_n16343), .A2(MEM_stage_inst_dmem_n19097), .ZN(MEM_stage_inst_dmem_n19066) );
INV_X1 MEM_stage_inst_dmem_U18018 ( .A(MEM_stage_inst_dmem_n19096), .ZN(MEM_stage_inst_dmem_n19097) );
NAND2_X1 MEM_stage_inst_dmem_U18017 ( .A1(MEM_stage_inst_dmem_ram_2655), .A2(MEM_stage_inst_dmem_n19096), .ZN(MEM_stage_inst_dmem_n19067) );
NAND2_X1 MEM_stage_inst_dmem_U18016 ( .A1(MEM_stage_inst_dmem_n21284), .A2(MEM_stage_inst_dmem_n19236), .ZN(MEM_stage_inst_dmem_n19096) );
NAND2_X1 MEM_stage_inst_dmem_U18015 ( .A1(MEM_stage_inst_dmem_n19065), .A2(MEM_stage_inst_dmem_n19064), .ZN(MEM_stage_inst_dmem_n9883) );
NAND2_X1 MEM_stage_inst_dmem_U18014 ( .A1(MEM_stage_inst_dmem_n19275), .A2(MEM_stage_inst_dmem_n19063), .ZN(MEM_stage_inst_dmem_n19064) );
NAND2_X1 MEM_stage_inst_dmem_U18013 ( .A1(MEM_stage_inst_dmem_ram_2656), .A2(MEM_stage_inst_dmem_n19062), .ZN(MEM_stage_inst_dmem_n19065) );
NAND2_X1 MEM_stage_inst_dmem_U18012 ( .A1(MEM_stage_inst_dmem_n19061), .A2(MEM_stage_inst_dmem_n19060), .ZN(MEM_stage_inst_dmem_n9884) );
NAND2_X1 MEM_stage_inst_dmem_U18011 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n19063), .ZN(MEM_stage_inst_dmem_n19060) );
NAND2_X1 MEM_stage_inst_dmem_U18010 ( .A1(MEM_stage_inst_dmem_ram_2657), .A2(MEM_stage_inst_dmem_n19062), .ZN(MEM_stage_inst_dmem_n19061) );
NAND2_X1 MEM_stage_inst_dmem_U18009 ( .A1(MEM_stage_inst_dmem_n19059), .A2(MEM_stage_inst_dmem_n19058), .ZN(MEM_stage_inst_dmem_n9885) );
NAND2_X1 MEM_stage_inst_dmem_U18008 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n19063), .ZN(MEM_stage_inst_dmem_n19058) );
NAND2_X1 MEM_stage_inst_dmem_U18007 ( .A1(MEM_stage_inst_dmem_ram_2658), .A2(MEM_stage_inst_dmem_n19062), .ZN(MEM_stage_inst_dmem_n19059) );
NAND2_X1 MEM_stage_inst_dmem_U18006 ( .A1(MEM_stage_inst_dmem_n19057), .A2(MEM_stage_inst_dmem_n19056), .ZN(MEM_stage_inst_dmem_n9886) );
NAND2_X1 MEM_stage_inst_dmem_U18005 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n19063), .ZN(MEM_stage_inst_dmem_n19056) );
NAND2_X1 MEM_stage_inst_dmem_U18004 ( .A1(MEM_stage_inst_dmem_ram_2659), .A2(MEM_stage_inst_dmem_n19062), .ZN(MEM_stage_inst_dmem_n19057) );
NAND2_X1 MEM_stage_inst_dmem_U18003 ( .A1(MEM_stage_inst_dmem_n19055), .A2(MEM_stage_inst_dmem_n19054), .ZN(MEM_stage_inst_dmem_n9887) );
NAND2_X1 MEM_stage_inst_dmem_U18002 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n19063), .ZN(MEM_stage_inst_dmem_n19054) );
NAND2_X1 MEM_stage_inst_dmem_U18001 ( .A1(MEM_stage_inst_dmem_ram_2660), .A2(MEM_stage_inst_dmem_n19062), .ZN(MEM_stage_inst_dmem_n19055) );
NAND2_X1 MEM_stage_inst_dmem_U18000 ( .A1(MEM_stage_inst_dmem_n19053), .A2(MEM_stage_inst_dmem_n19052), .ZN(MEM_stage_inst_dmem_n9888) );
NAND2_X1 MEM_stage_inst_dmem_U17999 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n19063), .ZN(MEM_stage_inst_dmem_n19052) );
NAND2_X1 MEM_stage_inst_dmem_U17998 ( .A1(MEM_stage_inst_dmem_ram_2661), .A2(MEM_stage_inst_dmem_n19062), .ZN(MEM_stage_inst_dmem_n19053) );
NAND2_X1 MEM_stage_inst_dmem_U17997 ( .A1(MEM_stage_inst_dmem_n19051), .A2(MEM_stage_inst_dmem_n19050), .ZN(MEM_stage_inst_dmem_n9889) );
NAND2_X1 MEM_stage_inst_dmem_U17996 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n19063), .ZN(MEM_stage_inst_dmem_n19050) );
NAND2_X1 MEM_stage_inst_dmem_U17995 ( .A1(MEM_stage_inst_dmem_ram_2662), .A2(MEM_stage_inst_dmem_n19062), .ZN(MEM_stage_inst_dmem_n19051) );
NAND2_X1 MEM_stage_inst_dmem_U17994 ( .A1(MEM_stage_inst_dmem_n19049), .A2(MEM_stage_inst_dmem_n19048), .ZN(MEM_stage_inst_dmem_n9890) );
NAND2_X1 MEM_stage_inst_dmem_U17993 ( .A1(MEM_stage_inst_dmem_n16777), .A2(MEM_stage_inst_dmem_n19063), .ZN(MEM_stage_inst_dmem_n19048) );
NAND2_X1 MEM_stage_inst_dmem_U17992 ( .A1(MEM_stage_inst_dmem_ram_2663), .A2(MEM_stage_inst_dmem_n19062), .ZN(MEM_stage_inst_dmem_n19049) );
NAND2_X1 MEM_stage_inst_dmem_U17991 ( .A1(MEM_stage_inst_dmem_n19047), .A2(MEM_stage_inst_dmem_n19046), .ZN(MEM_stage_inst_dmem_n9891) );
NAND2_X1 MEM_stage_inst_dmem_U17990 ( .A1(MEM_stage_inst_dmem_n18013), .A2(MEM_stage_inst_dmem_n19063), .ZN(MEM_stage_inst_dmem_n19046) );
NAND2_X1 MEM_stage_inst_dmem_U17989 ( .A1(MEM_stage_inst_dmem_ram_2664), .A2(MEM_stage_inst_dmem_n19062), .ZN(MEM_stage_inst_dmem_n19047) );
NAND2_X1 MEM_stage_inst_dmem_U17988 ( .A1(MEM_stage_inst_dmem_n19045), .A2(MEM_stage_inst_dmem_n19044), .ZN(MEM_stage_inst_dmem_n9892) );
NAND2_X1 MEM_stage_inst_dmem_U17987 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n19063), .ZN(MEM_stage_inst_dmem_n19044) );
NAND2_X1 MEM_stage_inst_dmem_U17986 ( .A1(MEM_stage_inst_dmem_ram_2665), .A2(MEM_stage_inst_dmem_n19062), .ZN(MEM_stage_inst_dmem_n19045) );
NAND2_X1 MEM_stage_inst_dmem_U17985 ( .A1(MEM_stage_inst_dmem_n19043), .A2(MEM_stage_inst_dmem_n19042), .ZN(MEM_stage_inst_dmem_n9893) );
NAND2_X1 MEM_stage_inst_dmem_U17984 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n19063), .ZN(MEM_stage_inst_dmem_n19042) );
NAND2_X1 MEM_stage_inst_dmem_U17983 ( .A1(MEM_stage_inst_dmem_ram_2666), .A2(MEM_stage_inst_dmem_n19062), .ZN(MEM_stage_inst_dmem_n19043) );
NAND2_X1 MEM_stage_inst_dmem_U17982 ( .A1(MEM_stage_inst_dmem_n19041), .A2(MEM_stage_inst_dmem_n19040), .ZN(MEM_stage_inst_dmem_n9894) );
NAND2_X1 MEM_stage_inst_dmem_U17981 ( .A1(MEM_stage_inst_dmem_n20904), .A2(MEM_stage_inst_dmem_n19063), .ZN(MEM_stage_inst_dmem_n19040) );
NAND2_X1 MEM_stage_inst_dmem_U17980 ( .A1(MEM_stage_inst_dmem_ram_2667), .A2(MEM_stage_inst_dmem_n19062), .ZN(MEM_stage_inst_dmem_n19041) );
NAND2_X1 MEM_stage_inst_dmem_U17979 ( .A1(MEM_stage_inst_dmem_n19039), .A2(MEM_stage_inst_dmem_n19038), .ZN(MEM_stage_inst_dmem_n9895) );
NAND2_X1 MEM_stage_inst_dmem_U17978 ( .A1(MEM_stage_inst_dmem_n21474), .A2(MEM_stage_inst_dmem_n19063), .ZN(MEM_stage_inst_dmem_n19038) );
NAND2_X1 MEM_stage_inst_dmem_U17977 ( .A1(MEM_stage_inst_dmem_ram_2668), .A2(MEM_stage_inst_dmem_n19062), .ZN(MEM_stage_inst_dmem_n19039) );
NAND2_X1 MEM_stage_inst_dmem_U17976 ( .A1(MEM_stage_inst_dmem_n19037), .A2(MEM_stage_inst_dmem_n19036), .ZN(MEM_stage_inst_dmem_n9896) );
NAND2_X1 MEM_stage_inst_dmem_U17975 ( .A1(MEM_stage_inst_dmem_n19242), .A2(MEM_stage_inst_dmem_n19063), .ZN(MEM_stage_inst_dmem_n19036) );
NAND2_X1 MEM_stage_inst_dmem_U17974 ( .A1(MEM_stage_inst_dmem_ram_2669), .A2(MEM_stage_inst_dmem_n19062), .ZN(MEM_stage_inst_dmem_n19037) );
NAND2_X1 MEM_stage_inst_dmem_U17973 ( .A1(MEM_stage_inst_dmem_n19035), .A2(MEM_stage_inst_dmem_n19034), .ZN(MEM_stage_inst_dmem_n9897) );
NAND2_X1 MEM_stage_inst_dmem_U17972 ( .A1(MEM_stage_inst_dmem_n115), .A2(MEM_stage_inst_dmem_n19063), .ZN(MEM_stage_inst_dmem_n19034) );
NAND2_X1 MEM_stage_inst_dmem_U17971 ( .A1(MEM_stage_inst_dmem_ram_2670), .A2(MEM_stage_inst_dmem_n19062), .ZN(MEM_stage_inst_dmem_n19035) );
NAND2_X1 MEM_stage_inst_dmem_U17970 ( .A1(MEM_stage_inst_dmem_n19033), .A2(MEM_stage_inst_dmem_n19032), .ZN(MEM_stage_inst_dmem_n9898) );
NAND2_X1 MEM_stage_inst_dmem_U17969 ( .A1(MEM_stage_inst_dmem_n21320), .A2(MEM_stage_inst_dmem_n19063), .ZN(MEM_stage_inst_dmem_n19032) );
INV_X1 MEM_stage_inst_dmem_U17968 ( .A(MEM_stage_inst_dmem_n19062), .ZN(MEM_stage_inst_dmem_n19063) );
NAND2_X1 MEM_stage_inst_dmem_U17967 ( .A1(MEM_stage_inst_dmem_ram_2671), .A2(MEM_stage_inst_dmem_n19062), .ZN(MEM_stage_inst_dmem_n19033) );
NAND2_X1 MEM_stage_inst_dmem_U17966 ( .A1(MEM_stage_inst_dmem_n21249), .A2(MEM_stage_inst_dmem_n19236), .ZN(MEM_stage_inst_dmem_n19062) );
NAND2_X1 MEM_stage_inst_dmem_U17965 ( .A1(MEM_stage_inst_dmem_n19031), .A2(MEM_stage_inst_dmem_n19030), .ZN(MEM_stage_inst_dmem_n9899) );
NAND2_X1 MEM_stage_inst_dmem_U17964 ( .A1(MEM_stage_inst_dmem_n19275), .A2(MEM_stage_inst_dmem_n19029), .ZN(MEM_stage_inst_dmem_n19030) );
NAND2_X1 MEM_stage_inst_dmem_U17963 ( .A1(MEM_stage_inst_dmem_ram_2672), .A2(MEM_stage_inst_dmem_n19028), .ZN(MEM_stage_inst_dmem_n19031) );
NAND2_X1 MEM_stage_inst_dmem_U17962 ( .A1(MEM_stage_inst_dmem_n19027), .A2(MEM_stage_inst_dmem_n19026), .ZN(MEM_stage_inst_dmem_n9900) );
NAND2_X1 MEM_stage_inst_dmem_U17961 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n19029), .ZN(MEM_stage_inst_dmem_n19026) );
NAND2_X1 MEM_stage_inst_dmem_U17960 ( .A1(MEM_stage_inst_dmem_ram_2673), .A2(MEM_stage_inst_dmem_n19028), .ZN(MEM_stage_inst_dmem_n19027) );
NAND2_X1 MEM_stage_inst_dmem_U17959 ( .A1(MEM_stage_inst_dmem_n19025), .A2(MEM_stage_inst_dmem_n19024), .ZN(MEM_stage_inst_dmem_n9901) );
NAND2_X1 MEM_stage_inst_dmem_U17958 ( .A1(MEM_stage_inst_dmem_n18027), .A2(MEM_stage_inst_dmem_n19029), .ZN(MEM_stage_inst_dmem_n19024) );
NAND2_X1 MEM_stage_inst_dmem_U17957 ( .A1(MEM_stage_inst_dmem_ram_2674), .A2(MEM_stage_inst_dmem_n19028), .ZN(MEM_stage_inst_dmem_n19025) );
NAND2_X1 MEM_stage_inst_dmem_U17956 ( .A1(MEM_stage_inst_dmem_n19023), .A2(MEM_stage_inst_dmem_n19022), .ZN(MEM_stage_inst_dmem_n9902) );
NAND2_X1 MEM_stage_inst_dmem_U17955 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n19029), .ZN(MEM_stage_inst_dmem_n19022) );
NAND2_X1 MEM_stage_inst_dmem_U17954 ( .A1(MEM_stage_inst_dmem_ram_2675), .A2(MEM_stage_inst_dmem_n19028), .ZN(MEM_stage_inst_dmem_n19023) );
NAND2_X1 MEM_stage_inst_dmem_U17953 ( .A1(MEM_stage_inst_dmem_n19021), .A2(MEM_stage_inst_dmem_n19020), .ZN(MEM_stage_inst_dmem_n9903) );
NAND2_X1 MEM_stage_inst_dmem_U17952 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n19029), .ZN(MEM_stage_inst_dmem_n19020) );
NAND2_X1 MEM_stage_inst_dmem_U17951 ( .A1(MEM_stage_inst_dmem_ram_2676), .A2(MEM_stage_inst_dmem_n19028), .ZN(MEM_stage_inst_dmem_n19021) );
NAND2_X1 MEM_stage_inst_dmem_U17950 ( .A1(MEM_stage_inst_dmem_n19019), .A2(MEM_stage_inst_dmem_n19018), .ZN(MEM_stage_inst_dmem_n9904) );
NAND2_X1 MEM_stage_inst_dmem_U17949 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n19029), .ZN(MEM_stage_inst_dmem_n19018) );
NAND2_X1 MEM_stage_inst_dmem_U17948 ( .A1(MEM_stage_inst_dmem_ram_2677), .A2(MEM_stage_inst_dmem_n19028), .ZN(MEM_stage_inst_dmem_n19019) );
NAND2_X1 MEM_stage_inst_dmem_U17947 ( .A1(MEM_stage_inst_dmem_n19017), .A2(MEM_stage_inst_dmem_n19016), .ZN(MEM_stage_inst_dmem_n9905) );
NAND2_X1 MEM_stage_inst_dmem_U17946 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n19029), .ZN(MEM_stage_inst_dmem_n19016) );
NAND2_X1 MEM_stage_inst_dmem_U17945 ( .A1(MEM_stage_inst_dmem_ram_2678), .A2(MEM_stage_inst_dmem_n19028), .ZN(MEM_stage_inst_dmem_n19017) );
NAND2_X1 MEM_stage_inst_dmem_U17944 ( .A1(MEM_stage_inst_dmem_n19015), .A2(MEM_stage_inst_dmem_n19014), .ZN(MEM_stage_inst_dmem_n9906) );
NAND2_X1 MEM_stage_inst_dmem_U17943 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n19029), .ZN(MEM_stage_inst_dmem_n19014) );
NAND2_X1 MEM_stage_inst_dmem_U17942 ( .A1(MEM_stage_inst_dmem_ram_2679), .A2(MEM_stage_inst_dmem_n19028), .ZN(MEM_stage_inst_dmem_n19015) );
NAND2_X1 MEM_stage_inst_dmem_U17941 ( .A1(MEM_stage_inst_dmem_n19013), .A2(MEM_stage_inst_dmem_n19012), .ZN(MEM_stage_inst_dmem_n9907) );
NAND2_X1 MEM_stage_inst_dmem_U17940 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n19029), .ZN(MEM_stage_inst_dmem_n19012) );
NAND2_X1 MEM_stage_inst_dmem_U17939 ( .A1(MEM_stage_inst_dmem_ram_2680), .A2(MEM_stage_inst_dmem_n19028), .ZN(MEM_stage_inst_dmem_n19013) );
NAND2_X1 MEM_stage_inst_dmem_U17938 ( .A1(MEM_stage_inst_dmem_n19011), .A2(MEM_stage_inst_dmem_n19010), .ZN(MEM_stage_inst_dmem_n9908) );
NAND2_X1 MEM_stage_inst_dmem_U17937 ( .A1(MEM_stage_inst_dmem_n19251), .A2(MEM_stage_inst_dmem_n19029), .ZN(MEM_stage_inst_dmem_n19010) );
NAND2_X1 MEM_stage_inst_dmem_U17936 ( .A1(MEM_stage_inst_dmem_ram_2681), .A2(MEM_stage_inst_dmem_n19028), .ZN(MEM_stage_inst_dmem_n19011) );
NAND2_X1 MEM_stage_inst_dmem_U17935 ( .A1(MEM_stage_inst_dmem_n19009), .A2(MEM_stage_inst_dmem_n19008), .ZN(MEM_stage_inst_dmem_n9909) );
NAND2_X1 MEM_stage_inst_dmem_U17934 ( .A1(MEM_stage_inst_dmem_n18007), .A2(MEM_stage_inst_dmem_n19029), .ZN(MEM_stage_inst_dmem_n19008) );
NAND2_X1 MEM_stage_inst_dmem_U17933 ( .A1(MEM_stage_inst_dmem_ram_2682), .A2(MEM_stage_inst_dmem_n19028), .ZN(MEM_stage_inst_dmem_n19009) );
NAND2_X1 MEM_stage_inst_dmem_U17932 ( .A1(MEM_stage_inst_dmem_n19007), .A2(MEM_stage_inst_dmem_n19006), .ZN(MEM_stage_inst_dmem_n9910) );
NAND2_X1 MEM_stage_inst_dmem_U17931 ( .A1(MEM_stage_inst_dmem_n14705), .A2(MEM_stage_inst_dmem_n19029), .ZN(MEM_stage_inst_dmem_n19006) );
NAND2_X1 MEM_stage_inst_dmem_U17930 ( .A1(MEM_stage_inst_dmem_ram_2683), .A2(MEM_stage_inst_dmem_n19028), .ZN(MEM_stage_inst_dmem_n19007) );
NAND2_X1 MEM_stage_inst_dmem_U17929 ( .A1(MEM_stage_inst_dmem_n19005), .A2(MEM_stage_inst_dmem_n19004), .ZN(MEM_stage_inst_dmem_n9911) );
NAND2_X1 MEM_stage_inst_dmem_U17928 ( .A1(MEM_stage_inst_dmem_n14702), .A2(MEM_stage_inst_dmem_n19029), .ZN(MEM_stage_inst_dmem_n19004) );
NAND2_X1 MEM_stage_inst_dmem_U17927 ( .A1(MEM_stage_inst_dmem_ram_2684), .A2(MEM_stage_inst_dmem_n19028), .ZN(MEM_stage_inst_dmem_n19005) );
NAND2_X1 MEM_stage_inst_dmem_U17926 ( .A1(MEM_stage_inst_dmem_n19003), .A2(MEM_stage_inst_dmem_n19002), .ZN(MEM_stage_inst_dmem_n9912) );
NAND2_X1 MEM_stage_inst_dmem_U17925 ( .A1(MEM_stage_inst_dmem_n19242), .A2(MEM_stage_inst_dmem_n19029), .ZN(MEM_stage_inst_dmem_n19002) );
NAND2_X1 MEM_stage_inst_dmem_U17924 ( .A1(MEM_stage_inst_dmem_ram_2685), .A2(MEM_stage_inst_dmem_n19028), .ZN(MEM_stage_inst_dmem_n19003) );
NAND2_X1 MEM_stage_inst_dmem_U17923 ( .A1(MEM_stage_inst_dmem_n19001), .A2(MEM_stage_inst_dmem_n19000), .ZN(MEM_stage_inst_dmem_n9913) );
NAND2_X1 MEM_stage_inst_dmem_U17922 ( .A1(MEM_stage_inst_dmem_n115), .A2(MEM_stage_inst_dmem_n19029), .ZN(MEM_stage_inst_dmem_n19000) );
NAND2_X1 MEM_stage_inst_dmem_U17921 ( .A1(MEM_stage_inst_dmem_ram_2686), .A2(MEM_stage_inst_dmem_n19028), .ZN(MEM_stage_inst_dmem_n19001) );
NAND2_X1 MEM_stage_inst_dmem_U17920 ( .A1(MEM_stage_inst_dmem_n18999), .A2(MEM_stage_inst_dmem_n18998), .ZN(MEM_stage_inst_dmem_n9914) );
NAND2_X1 MEM_stage_inst_dmem_U17919 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n19029), .ZN(MEM_stage_inst_dmem_n18998) );
INV_X1 MEM_stage_inst_dmem_U17918 ( .A(MEM_stage_inst_dmem_n19028), .ZN(MEM_stage_inst_dmem_n19029) );
NAND2_X1 MEM_stage_inst_dmem_U17917 ( .A1(MEM_stage_inst_dmem_ram_2687), .A2(MEM_stage_inst_dmem_n19028), .ZN(MEM_stage_inst_dmem_n18999) );
NAND2_X1 MEM_stage_inst_dmem_U17916 ( .A1(MEM_stage_inst_dmem_n21214), .A2(MEM_stage_inst_dmem_n19236), .ZN(MEM_stage_inst_dmem_n19028) );
NAND2_X1 MEM_stage_inst_dmem_U17915 ( .A1(MEM_stage_inst_dmem_n18997), .A2(MEM_stage_inst_dmem_n18996), .ZN(MEM_stage_inst_dmem_n9915) );
NAND2_X1 MEM_stage_inst_dmem_U17914 ( .A1(MEM_stage_inst_dmem_n19275), .A2(MEM_stage_inst_dmem_n18995), .ZN(MEM_stage_inst_dmem_n18996) );
NAND2_X1 MEM_stage_inst_dmem_U17913 ( .A1(MEM_stage_inst_dmem_ram_2688), .A2(MEM_stage_inst_dmem_n18994), .ZN(MEM_stage_inst_dmem_n18997) );
NAND2_X1 MEM_stage_inst_dmem_U17912 ( .A1(MEM_stage_inst_dmem_n18993), .A2(MEM_stage_inst_dmem_n18992), .ZN(MEM_stage_inst_dmem_n9916) );
NAND2_X1 MEM_stage_inst_dmem_U17911 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n18995), .ZN(MEM_stage_inst_dmem_n18992) );
NAND2_X1 MEM_stage_inst_dmem_U17910 ( .A1(MEM_stage_inst_dmem_ram_2689), .A2(MEM_stage_inst_dmem_n18994), .ZN(MEM_stage_inst_dmem_n18993) );
NAND2_X1 MEM_stage_inst_dmem_U17909 ( .A1(MEM_stage_inst_dmem_n18991), .A2(MEM_stage_inst_dmem_n18990), .ZN(MEM_stage_inst_dmem_n9917) );
NAND2_X1 MEM_stage_inst_dmem_U17908 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n18995), .ZN(MEM_stage_inst_dmem_n18990) );
NAND2_X1 MEM_stage_inst_dmem_U17907 ( .A1(MEM_stage_inst_dmem_ram_2690), .A2(MEM_stage_inst_dmem_n18994), .ZN(MEM_stage_inst_dmem_n18991) );
NAND2_X1 MEM_stage_inst_dmem_U17906 ( .A1(MEM_stage_inst_dmem_n18989), .A2(MEM_stage_inst_dmem_n18988), .ZN(MEM_stage_inst_dmem_n9918) );
NAND2_X1 MEM_stage_inst_dmem_U17905 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n18995), .ZN(MEM_stage_inst_dmem_n18988) );
NAND2_X1 MEM_stage_inst_dmem_U17904 ( .A1(MEM_stage_inst_dmem_ram_2691), .A2(MEM_stage_inst_dmem_n18994), .ZN(MEM_stage_inst_dmem_n18989) );
NAND2_X1 MEM_stage_inst_dmem_U17903 ( .A1(MEM_stage_inst_dmem_n18987), .A2(MEM_stage_inst_dmem_n18986), .ZN(MEM_stage_inst_dmem_n9919) );
NAND2_X1 MEM_stage_inst_dmem_U17902 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n18995), .ZN(MEM_stage_inst_dmem_n18986) );
NAND2_X1 MEM_stage_inst_dmem_U17901 ( .A1(MEM_stage_inst_dmem_ram_2692), .A2(MEM_stage_inst_dmem_n18994), .ZN(MEM_stage_inst_dmem_n18987) );
NAND2_X1 MEM_stage_inst_dmem_U17900 ( .A1(MEM_stage_inst_dmem_n18985), .A2(MEM_stage_inst_dmem_n18984), .ZN(MEM_stage_inst_dmem_n9920) );
NAND2_X1 MEM_stage_inst_dmem_U17899 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n18995), .ZN(MEM_stage_inst_dmem_n18984) );
NAND2_X1 MEM_stage_inst_dmem_U17898 ( .A1(MEM_stage_inst_dmem_ram_2693), .A2(MEM_stage_inst_dmem_n18994), .ZN(MEM_stage_inst_dmem_n18985) );
NAND2_X1 MEM_stage_inst_dmem_U17897 ( .A1(MEM_stage_inst_dmem_n18983), .A2(MEM_stage_inst_dmem_n18982), .ZN(MEM_stage_inst_dmem_n9921) );
NAND2_X1 MEM_stage_inst_dmem_U17896 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n18995), .ZN(MEM_stage_inst_dmem_n18982) );
NAND2_X1 MEM_stage_inst_dmem_U17895 ( .A1(MEM_stage_inst_dmem_ram_2694), .A2(MEM_stage_inst_dmem_n18994), .ZN(MEM_stage_inst_dmem_n18983) );
NAND2_X1 MEM_stage_inst_dmem_U17894 ( .A1(MEM_stage_inst_dmem_n18981), .A2(MEM_stage_inst_dmem_n18980), .ZN(MEM_stage_inst_dmem_n9922) );
NAND2_X1 MEM_stage_inst_dmem_U17893 ( .A1(MEM_stage_inst_dmem_n18), .A2(MEM_stage_inst_dmem_n18995), .ZN(MEM_stage_inst_dmem_n18980) );
NAND2_X1 MEM_stage_inst_dmem_U17892 ( .A1(MEM_stage_inst_dmem_ram_2695), .A2(MEM_stage_inst_dmem_n18994), .ZN(MEM_stage_inst_dmem_n18981) );
NAND2_X1 MEM_stage_inst_dmem_U17891 ( .A1(MEM_stage_inst_dmem_n18979), .A2(MEM_stage_inst_dmem_n18978), .ZN(MEM_stage_inst_dmem_n9923) );
NAND2_X1 MEM_stage_inst_dmem_U17890 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n18995), .ZN(MEM_stage_inst_dmem_n18978) );
NAND2_X1 MEM_stage_inst_dmem_U17889 ( .A1(MEM_stage_inst_dmem_ram_2696), .A2(MEM_stage_inst_dmem_n18994), .ZN(MEM_stage_inst_dmem_n18979) );
NAND2_X1 MEM_stage_inst_dmem_U17888 ( .A1(MEM_stage_inst_dmem_n18977), .A2(MEM_stage_inst_dmem_n18976), .ZN(MEM_stage_inst_dmem_n9924) );
NAND2_X1 MEM_stage_inst_dmem_U17887 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n18995), .ZN(MEM_stage_inst_dmem_n18976) );
NAND2_X1 MEM_stage_inst_dmem_U17886 ( .A1(MEM_stage_inst_dmem_ram_2697), .A2(MEM_stage_inst_dmem_n18994), .ZN(MEM_stage_inst_dmem_n18977) );
NAND2_X1 MEM_stage_inst_dmem_U17885 ( .A1(MEM_stage_inst_dmem_n18975), .A2(MEM_stage_inst_dmem_n18974), .ZN(MEM_stage_inst_dmem_n9925) );
NAND2_X1 MEM_stage_inst_dmem_U17884 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n18995), .ZN(MEM_stage_inst_dmem_n18974) );
NAND2_X1 MEM_stage_inst_dmem_U17883 ( .A1(MEM_stage_inst_dmem_ram_2698), .A2(MEM_stage_inst_dmem_n18994), .ZN(MEM_stage_inst_dmem_n18975) );
NAND2_X1 MEM_stage_inst_dmem_U17882 ( .A1(MEM_stage_inst_dmem_n18973), .A2(MEM_stage_inst_dmem_n18972), .ZN(MEM_stage_inst_dmem_n9926) );
NAND2_X1 MEM_stage_inst_dmem_U17881 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n18995), .ZN(MEM_stage_inst_dmem_n18972) );
NAND2_X1 MEM_stage_inst_dmem_U17880 ( .A1(MEM_stage_inst_dmem_ram_2699), .A2(MEM_stage_inst_dmem_n18994), .ZN(MEM_stage_inst_dmem_n18973) );
NAND2_X1 MEM_stage_inst_dmem_U17879 ( .A1(MEM_stage_inst_dmem_n18971), .A2(MEM_stage_inst_dmem_n18970), .ZN(MEM_stage_inst_dmem_n9927) );
NAND2_X1 MEM_stage_inst_dmem_U17878 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n18995), .ZN(MEM_stage_inst_dmem_n18970) );
NAND2_X1 MEM_stage_inst_dmem_U17877 ( .A1(MEM_stage_inst_dmem_ram_2700), .A2(MEM_stage_inst_dmem_n18994), .ZN(MEM_stage_inst_dmem_n18971) );
NAND2_X1 MEM_stage_inst_dmem_U17876 ( .A1(MEM_stage_inst_dmem_n18969), .A2(MEM_stage_inst_dmem_n18968), .ZN(MEM_stage_inst_dmem_n9928) );
NAND2_X1 MEM_stage_inst_dmem_U17875 ( .A1(MEM_stage_inst_dmem_n19242), .A2(MEM_stage_inst_dmem_n18995), .ZN(MEM_stage_inst_dmem_n18968) );
NAND2_X1 MEM_stage_inst_dmem_U17874 ( .A1(MEM_stage_inst_dmem_ram_2701), .A2(MEM_stage_inst_dmem_n18994), .ZN(MEM_stage_inst_dmem_n18969) );
NAND2_X1 MEM_stage_inst_dmem_U17873 ( .A1(MEM_stage_inst_dmem_n18967), .A2(MEM_stage_inst_dmem_n18966), .ZN(MEM_stage_inst_dmem_n9929) );
NAND2_X1 MEM_stage_inst_dmem_U17872 ( .A1(MEM_stage_inst_dmem_n115), .A2(MEM_stage_inst_dmem_n18995), .ZN(MEM_stage_inst_dmem_n18966) );
NAND2_X1 MEM_stage_inst_dmem_U17871 ( .A1(MEM_stage_inst_dmem_ram_2702), .A2(MEM_stage_inst_dmem_n18994), .ZN(MEM_stage_inst_dmem_n18967) );
NAND2_X1 MEM_stage_inst_dmem_U17870 ( .A1(MEM_stage_inst_dmem_n18965), .A2(MEM_stage_inst_dmem_n18964), .ZN(MEM_stage_inst_dmem_n9930) );
NAND2_X1 MEM_stage_inst_dmem_U17869 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n18995), .ZN(MEM_stage_inst_dmem_n18964) );
INV_X1 MEM_stage_inst_dmem_U17868 ( .A(MEM_stage_inst_dmem_n18994), .ZN(MEM_stage_inst_dmem_n18995) );
NAND2_X1 MEM_stage_inst_dmem_U17867 ( .A1(MEM_stage_inst_dmem_ram_2703), .A2(MEM_stage_inst_dmem_n18994), .ZN(MEM_stage_inst_dmem_n18965) );
NAND2_X1 MEM_stage_inst_dmem_U17866 ( .A1(MEM_stage_inst_dmem_n21179), .A2(MEM_stage_inst_dmem_n19236), .ZN(MEM_stage_inst_dmem_n18994) );
NAND2_X1 MEM_stage_inst_dmem_U17865 ( .A1(MEM_stage_inst_dmem_n18963), .A2(MEM_stage_inst_dmem_n18962), .ZN(MEM_stage_inst_dmem_n9931) );
NAND2_X1 MEM_stage_inst_dmem_U17864 ( .A1(MEM_stage_inst_dmem_n19275), .A2(MEM_stage_inst_dmem_n18961), .ZN(MEM_stage_inst_dmem_n18962) );
NAND2_X1 MEM_stage_inst_dmem_U17863 ( .A1(MEM_stage_inst_dmem_ram_2704), .A2(MEM_stage_inst_dmem_n18960), .ZN(MEM_stage_inst_dmem_n18963) );
NAND2_X1 MEM_stage_inst_dmem_U17862 ( .A1(MEM_stage_inst_dmem_n18959), .A2(MEM_stage_inst_dmem_n18958), .ZN(MEM_stage_inst_dmem_n9932) );
NAND2_X1 MEM_stage_inst_dmem_U17861 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n18961), .ZN(MEM_stage_inst_dmem_n18958) );
NAND2_X1 MEM_stage_inst_dmem_U17860 ( .A1(MEM_stage_inst_dmem_ram_2705), .A2(MEM_stage_inst_dmem_n18960), .ZN(MEM_stage_inst_dmem_n18959) );
NAND2_X1 MEM_stage_inst_dmem_U17859 ( .A1(MEM_stage_inst_dmem_n18957), .A2(MEM_stage_inst_dmem_n18956), .ZN(MEM_stage_inst_dmem_n9933) );
NAND2_X1 MEM_stage_inst_dmem_U17858 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n18961), .ZN(MEM_stage_inst_dmem_n18956) );
NAND2_X1 MEM_stage_inst_dmem_U17857 ( .A1(MEM_stage_inst_dmem_ram_2706), .A2(MEM_stage_inst_dmem_n18960), .ZN(MEM_stage_inst_dmem_n18957) );
NAND2_X1 MEM_stage_inst_dmem_U17856 ( .A1(MEM_stage_inst_dmem_n18955), .A2(MEM_stage_inst_dmem_n18954), .ZN(MEM_stage_inst_dmem_n9934) );
NAND2_X1 MEM_stage_inst_dmem_U17855 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n18961), .ZN(MEM_stage_inst_dmem_n18954) );
NAND2_X1 MEM_stage_inst_dmem_U17854 ( .A1(MEM_stage_inst_dmem_ram_2707), .A2(MEM_stage_inst_dmem_n18960), .ZN(MEM_stage_inst_dmem_n18955) );
NAND2_X1 MEM_stage_inst_dmem_U17853 ( .A1(MEM_stage_inst_dmem_n18953), .A2(MEM_stage_inst_dmem_n18952), .ZN(MEM_stage_inst_dmem_n9935) );
NAND2_X1 MEM_stage_inst_dmem_U17852 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n18961), .ZN(MEM_stage_inst_dmem_n18952) );
NAND2_X1 MEM_stage_inst_dmem_U17851 ( .A1(MEM_stage_inst_dmem_ram_2708), .A2(MEM_stage_inst_dmem_n18960), .ZN(MEM_stage_inst_dmem_n18953) );
NAND2_X1 MEM_stage_inst_dmem_U17850 ( .A1(MEM_stage_inst_dmem_n18951), .A2(MEM_stage_inst_dmem_n18950), .ZN(MEM_stage_inst_dmem_n9936) );
NAND2_X1 MEM_stage_inst_dmem_U17849 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n18961), .ZN(MEM_stage_inst_dmem_n18950) );
NAND2_X1 MEM_stage_inst_dmem_U17848 ( .A1(MEM_stage_inst_dmem_ram_2709), .A2(MEM_stage_inst_dmem_n18960), .ZN(MEM_stage_inst_dmem_n18951) );
NAND2_X1 MEM_stage_inst_dmem_U17847 ( .A1(MEM_stage_inst_dmem_n18949), .A2(MEM_stage_inst_dmem_n18948), .ZN(MEM_stage_inst_dmem_n9937) );
NAND2_X1 MEM_stage_inst_dmem_U17846 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n18961), .ZN(MEM_stage_inst_dmem_n18948) );
NAND2_X1 MEM_stage_inst_dmem_U17845 ( .A1(MEM_stage_inst_dmem_ram_2710), .A2(MEM_stage_inst_dmem_n18960), .ZN(MEM_stage_inst_dmem_n18949) );
NAND2_X1 MEM_stage_inst_dmem_U17844 ( .A1(MEM_stage_inst_dmem_n18947), .A2(MEM_stage_inst_dmem_n18946), .ZN(MEM_stage_inst_dmem_n9938) );
NAND2_X1 MEM_stage_inst_dmem_U17843 ( .A1(MEM_stage_inst_dmem_n17), .A2(MEM_stage_inst_dmem_n18961), .ZN(MEM_stage_inst_dmem_n18946) );
NAND2_X1 MEM_stage_inst_dmem_U17842 ( .A1(MEM_stage_inst_dmem_ram_2711), .A2(MEM_stage_inst_dmem_n18960), .ZN(MEM_stage_inst_dmem_n18947) );
NAND2_X1 MEM_stage_inst_dmem_U17841 ( .A1(MEM_stage_inst_dmem_n18945), .A2(MEM_stage_inst_dmem_n18944), .ZN(MEM_stage_inst_dmem_n9939) );
NAND2_X1 MEM_stage_inst_dmem_U17840 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n18961), .ZN(MEM_stage_inst_dmem_n18944) );
NAND2_X1 MEM_stage_inst_dmem_U17839 ( .A1(MEM_stage_inst_dmem_ram_2712), .A2(MEM_stage_inst_dmem_n18960), .ZN(MEM_stage_inst_dmem_n18945) );
NAND2_X1 MEM_stage_inst_dmem_U17838 ( .A1(MEM_stage_inst_dmem_n18943), .A2(MEM_stage_inst_dmem_n18942), .ZN(MEM_stage_inst_dmem_n9940) );
NAND2_X1 MEM_stage_inst_dmem_U17837 ( .A1(MEM_stage_inst_dmem_n19251), .A2(MEM_stage_inst_dmem_n18961), .ZN(MEM_stage_inst_dmem_n18942) );
NAND2_X1 MEM_stage_inst_dmem_U17836 ( .A1(MEM_stage_inst_dmem_ram_2713), .A2(MEM_stage_inst_dmem_n18960), .ZN(MEM_stage_inst_dmem_n18943) );
NAND2_X1 MEM_stage_inst_dmem_U17835 ( .A1(MEM_stage_inst_dmem_n18941), .A2(MEM_stage_inst_dmem_n18940), .ZN(MEM_stage_inst_dmem_n9941) );
NAND2_X1 MEM_stage_inst_dmem_U17834 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n18961), .ZN(MEM_stage_inst_dmem_n18940) );
NAND2_X1 MEM_stage_inst_dmem_U17833 ( .A1(MEM_stage_inst_dmem_ram_2714), .A2(MEM_stage_inst_dmem_n18960), .ZN(MEM_stage_inst_dmem_n18941) );
NAND2_X1 MEM_stage_inst_dmem_U17832 ( .A1(MEM_stage_inst_dmem_n18939), .A2(MEM_stage_inst_dmem_n18938), .ZN(MEM_stage_inst_dmem_n9942) );
NAND2_X1 MEM_stage_inst_dmem_U17831 ( .A1(MEM_stage_inst_dmem_n20904), .A2(MEM_stage_inst_dmem_n18961), .ZN(MEM_stage_inst_dmem_n18938) );
NAND2_X1 MEM_stage_inst_dmem_U17830 ( .A1(MEM_stage_inst_dmem_ram_2715), .A2(MEM_stage_inst_dmem_n18960), .ZN(MEM_stage_inst_dmem_n18939) );
NAND2_X1 MEM_stage_inst_dmem_U17829 ( .A1(MEM_stage_inst_dmem_n18937), .A2(MEM_stage_inst_dmem_n18936), .ZN(MEM_stage_inst_dmem_n9943) );
NAND2_X1 MEM_stage_inst_dmem_U17828 ( .A1(MEM_stage_inst_dmem_n21474), .A2(MEM_stage_inst_dmem_n18961), .ZN(MEM_stage_inst_dmem_n18936) );
NAND2_X1 MEM_stage_inst_dmem_U17827 ( .A1(MEM_stage_inst_dmem_ram_2716), .A2(MEM_stage_inst_dmem_n18960), .ZN(MEM_stage_inst_dmem_n18937) );
NAND2_X1 MEM_stage_inst_dmem_U17826 ( .A1(MEM_stage_inst_dmem_n18935), .A2(MEM_stage_inst_dmem_n18934), .ZN(MEM_stage_inst_dmem_n9944) );
NAND2_X1 MEM_stage_inst_dmem_U17825 ( .A1(MEM_stage_inst_dmem_n19242), .A2(MEM_stage_inst_dmem_n18961), .ZN(MEM_stage_inst_dmem_n18934) );
NAND2_X1 MEM_stage_inst_dmem_U17824 ( .A1(MEM_stage_inst_dmem_ram_2717), .A2(MEM_stage_inst_dmem_n18960), .ZN(MEM_stage_inst_dmem_n18935) );
NAND2_X1 MEM_stage_inst_dmem_U17823 ( .A1(MEM_stage_inst_dmem_n18933), .A2(MEM_stage_inst_dmem_n18932), .ZN(MEM_stage_inst_dmem_n9945) );
NAND2_X1 MEM_stage_inst_dmem_U17822 ( .A1(MEM_stage_inst_dmem_n115), .A2(MEM_stage_inst_dmem_n18961), .ZN(MEM_stage_inst_dmem_n18932) );
NAND2_X1 MEM_stage_inst_dmem_U17821 ( .A1(MEM_stage_inst_dmem_ram_2718), .A2(MEM_stage_inst_dmem_n18960), .ZN(MEM_stage_inst_dmem_n18933) );
NAND2_X1 MEM_stage_inst_dmem_U17820 ( .A1(MEM_stage_inst_dmem_n18931), .A2(MEM_stage_inst_dmem_n18930), .ZN(MEM_stage_inst_dmem_n9946) );
NAND2_X1 MEM_stage_inst_dmem_U17819 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n18961), .ZN(MEM_stage_inst_dmem_n18930) );
INV_X1 MEM_stage_inst_dmem_U17818 ( .A(MEM_stage_inst_dmem_n18960), .ZN(MEM_stage_inst_dmem_n18961) );
NAND2_X1 MEM_stage_inst_dmem_U17817 ( .A1(MEM_stage_inst_dmem_ram_2719), .A2(MEM_stage_inst_dmem_n18960), .ZN(MEM_stage_inst_dmem_n18931) );
NAND2_X1 MEM_stage_inst_dmem_U17816 ( .A1(MEM_stage_inst_dmem_n21144), .A2(MEM_stage_inst_dmem_n19236), .ZN(MEM_stage_inst_dmem_n18960) );
NAND2_X1 MEM_stage_inst_dmem_U17815 ( .A1(MEM_stage_inst_dmem_n18929), .A2(MEM_stage_inst_dmem_n18928), .ZN(MEM_stage_inst_dmem_n9947) );
NAND2_X1 MEM_stage_inst_dmem_U17814 ( .A1(MEM_stage_inst_dmem_n14732), .A2(MEM_stage_inst_dmem_n18927), .ZN(MEM_stage_inst_dmem_n18928) );
NAND2_X1 MEM_stage_inst_dmem_U17813 ( .A1(MEM_stage_inst_dmem_ram_2720), .A2(MEM_stage_inst_dmem_n18926), .ZN(MEM_stage_inst_dmem_n18929) );
NAND2_X1 MEM_stage_inst_dmem_U17812 ( .A1(MEM_stage_inst_dmem_n18925), .A2(MEM_stage_inst_dmem_n18924), .ZN(MEM_stage_inst_dmem_n9948) );
NAND2_X1 MEM_stage_inst_dmem_U17811 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n18927), .ZN(MEM_stage_inst_dmem_n18924) );
NAND2_X1 MEM_stage_inst_dmem_U17810 ( .A1(MEM_stage_inst_dmem_ram_2721), .A2(MEM_stage_inst_dmem_n18926), .ZN(MEM_stage_inst_dmem_n18925) );
NAND2_X1 MEM_stage_inst_dmem_U17809 ( .A1(MEM_stage_inst_dmem_n18923), .A2(MEM_stage_inst_dmem_n18922), .ZN(MEM_stage_inst_dmem_n9949) );
NAND2_X1 MEM_stage_inst_dmem_U17808 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n18927), .ZN(MEM_stage_inst_dmem_n18922) );
NAND2_X1 MEM_stage_inst_dmem_U17807 ( .A1(MEM_stage_inst_dmem_ram_2722), .A2(MEM_stage_inst_dmem_n18926), .ZN(MEM_stage_inst_dmem_n18923) );
NAND2_X1 MEM_stage_inst_dmem_U17806 ( .A1(MEM_stage_inst_dmem_n18921), .A2(MEM_stage_inst_dmem_n18920), .ZN(MEM_stage_inst_dmem_n9950) );
NAND2_X1 MEM_stage_inst_dmem_U17805 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n18927), .ZN(MEM_stage_inst_dmem_n18920) );
NAND2_X1 MEM_stage_inst_dmem_U17804 ( .A1(MEM_stage_inst_dmem_ram_2723), .A2(MEM_stage_inst_dmem_n18926), .ZN(MEM_stage_inst_dmem_n18921) );
NAND2_X1 MEM_stage_inst_dmem_U17803 ( .A1(MEM_stage_inst_dmem_n18919), .A2(MEM_stage_inst_dmem_n18918), .ZN(MEM_stage_inst_dmem_n9951) );
NAND2_X1 MEM_stage_inst_dmem_U17802 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n18927), .ZN(MEM_stage_inst_dmem_n18918) );
NAND2_X1 MEM_stage_inst_dmem_U17801 ( .A1(MEM_stage_inst_dmem_ram_2724), .A2(MEM_stage_inst_dmem_n18926), .ZN(MEM_stage_inst_dmem_n18919) );
NAND2_X1 MEM_stage_inst_dmem_U17800 ( .A1(MEM_stage_inst_dmem_n18917), .A2(MEM_stage_inst_dmem_n18916), .ZN(MEM_stage_inst_dmem_n9952) );
NAND2_X1 MEM_stage_inst_dmem_U17799 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n18927), .ZN(MEM_stage_inst_dmem_n18916) );
NAND2_X1 MEM_stage_inst_dmem_U17798 ( .A1(MEM_stage_inst_dmem_ram_2725), .A2(MEM_stage_inst_dmem_n18926), .ZN(MEM_stage_inst_dmem_n18917) );
NAND2_X1 MEM_stage_inst_dmem_U17797 ( .A1(MEM_stage_inst_dmem_n18915), .A2(MEM_stage_inst_dmem_n18914), .ZN(MEM_stage_inst_dmem_n9953) );
NAND2_X1 MEM_stage_inst_dmem_U17796 ( .A1(MEM_stage_inst_dmem_n21340), .A2(MEM_stage_inst_dmem_n18927), .ZN(MEM_stage_inst_dmem_n18914) );
NAND2_X1 MEM_stage_inst_dmem_U17795 ( .A1(MEM_stage_inst_dmem_ram_2726), .A2(MEM_stage_inst_dmem_n18926), .ZN(MEM_stage_inst_dmem_n18915) );
NAND2_X1 MEM_stage_inst_dmem_U17794 ( .A1(MEM_stage_inst_dmem_n18913), .A2(MEM_stage_inst_dmem_n18912), .ZN(MEM_stage_inst_dmem_n9954) );
NAND2_X1 MEM_stage_inst_dmem_U17793 ( .A1(MEM_stage_inst_dmem_n17), .A2(MEM_stage_inst_dmem_n18927), .ZN(MEM_stage_inst_dmem_n18912) );
NAND2_X1 MEM_stage_inst_dmem_U17792 ( .A1(MEM_stage_inst_dmem_ram_2727), .A2(MEM_stage_inst_dmem_n18926), .ZN(MEM_stage_inst_dmem_n18913) );
NAND2_X1 MEM_stage_inst_dmem_U17791 ( .A1(MEM_stage_inst_dmem_n18911), .A2(MEM_stage_inst_dmem_n18910), .ZN(MEM_stage_inst_dmem_n9955) );
NAND2_X1 MEM_stage_inst_dmem_U17790 ( .A1(MEM_stage_inst_dmem_n21335), .A2(MEM_stage_inst_dmem_n18927), .ZN(MEM_stage_inst_dmem_n18910) );
NAND2_X1 MEM_stage_inst_dmem_U17789 ( .A1(MEM_stage_inst_dmem_ram_2728), .A2(MEM_stage_inst_dmem_n18926), .ZN(MEM_stage_inst_dmem_n18911) );
NAND2_X1 MEM_stage_inst_dmem_U17788 ( .A1(MEM_stage_inst_dmem_n18909), .A2(MEM_stage_inst_dmem_n18908), .ZN(MEM_stage_inst_dmem_n9956) );
NAND2_X1 MEM_stage_inst_dmem_U17787 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n18927), .ZN(MEM_stage_inst_dmem_n18908) );
NAND2_X1 MEM_stage_inst_dmem_U17786 ( .A1(MEM_stage_inst_dmem_ram_2729), .A2(MEM_stage_inst_dmem_n18926), .ZN(MEM_stage_inst_dmem_n18909) );
NAND2_X1 MEM_stage_inst_dmem_U17785 ( .A1(MEM_stage_inst_dmem_n18907), .A2(MEM_stage_inst_dmem_n18906), .ZN(MEM_stage_inst_dmem_n9957) );
NAND2_X1 MEM_stage_inst_dmem_U17784 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n18927), .ZN(MEM_stage_inst_dmem_n18906) );
NAND2_X1 MEM_stage_inst_dmem_U17783 ( .A1(MEM_stage_inst_dmem_ram_2730), .A2(MEM_stage_inst_dmem_n18926), .ZN(MEM_stage_inst_dmem_n18907) );
NAND2_X1 MEM_stage_inst_dmem_U17782 ( .A1(MEM_stage_inst_dmem_n18905), .A2(MEM_stage_inst_dmem_n18904), .ZN(MEM_stage_inst_dmem_n9958) );
NAND2_X1 MEM_stage_inst_dmem_U17781 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n18927), .ZN(MEM_stage_inst_dmem_n18904) );
NAND2_X1 MEM_stage_inst_dmem_U17780 ( .A1(MEM_stage_inst_dmem_ram_2731), .A2(MEM_stage_inst_dmem_n18926), .ZN(MEM_stage_inst_dmem_n18905) );
NAND2_X1 MEM_stage_inst_dmem_U17779 ( .A1(MEM_stage_inst_dmem_n18903), .A2(MEM_stage_inst_dmem_n18902), .ZN(MEM_stage_inst_dmem_n9959) );
NAND2_X1 MEM_stage_inst_dmem_U17778 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n18927), .ZN(MEM_stage_inst_dmem_n18902) );
NAND2_X1 MEM_stage_inst_dmem_U17777 ( .A1(MEM_stage_inst_dmem_ram_2732), .A2(MEM_stage_inst_dmem_n18926), .ZN(MEM_stage_inst_dmem_n18903) );
NAND2_X1 MEM_stage_inst_dmem_U17776 ( .A1(MEM_stage_inst_dmem_n18901), .A2(MEM_stage_inst_dmem_n18900), .ZN(MEM_stage_inst_dmem_n9960) );
NAND2_X1 MEM_stage_inst_dmem_U17775 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n18927), .ZN(MEM_stage_inst_dmem_n18900) );
NAND2_X1 MEM_stage_inst_dmem_U17774 ( .A1(MEM_stage_inst_dmem_ram_2733), .A2(MEM_stage_inst_dmem_n18926), .ZN(MEM_stage_inst_dmem_n18901) );
NAND2_X1 MEM_stage_inst_dmem_U17773 ( .A1(MEM_stage_inst_dmem_n18899), .A2(MEM_stage_inst_dmem_n18898), .ZN(MEM_stage_inst_dmem_n9961) );
NAND2_X1 MEM_stage_inst_dmem_U17772 ( .A1(MEM_stage_inst_dmem_n14696), .A2(MEM_stage_inst_dmem_n18927), .ZN(MEM_stage_inst_dmem_n18898) );
NAND2_X1 MEM_stage_inst_dmem_U17771 ( .A1(MEM_stage_inst_dmem_ram_2734), .A2(MEM_stage_inst_dmem_n18926), .ZN(MEM_stage_inst_dmem_n18899) );
NAND2_X1 MEM_stage_inst_dmem_U17770 ( .A1(MEM_stage_inst_dmem_n18897), .A2(MEM_stage_inst_dmem_n18896), .ZN(MEM_stage_inst_dmem_n9962) );
NAND2_X1 MEM_stage_inst_dmem_U17769 ( .A1(MEM_stage_inst_dmem_n21320), .A2(MEM_stage_inst_dmem_n18927), .ZN(MEM_stage_inst_dmem_n18896) );
INV_X1 MEM_stage_inst_dmem_U17768 ( .A(MEM_stage_inst_dmem_n18926), .ZN(MEM_stage_inst_dmem_n18927) );
NAND2_X1 MEM_stage_inst_dmem_U17767 ( .A1(MEM_stage_inst_dmem_ram_2735), .A2(MEM_stage_inst_dmem_n18926), .ZN(MEM_stage_inst_dmem_n18897) );
NAND2_X1 MEM_stage_inst_dmem_U17766 ( .A1(MEM_stage_inst_dmem_n21109), .A2(MEM_stage_inst_dmem_n19236), .ZN(MEM_stage_inst_dmem_n18926) );
NAND2_X1 MEM_stage_inst_dmem_U17765 ( .A1(MEM_stage_inst_dmem_n18895), .A2(MEM_stage_inst_dmem_n18894), .ZN(MEM_stage_inst_dmem_n9963) );
NAND2_X1 MEM_stage_inst_dmem_U17764 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n18893), .ZN(MEM_stage_inst_dmem_n18894) );
NAND2_X1 MEM_stage_inst_dmem_U17763 ( .A1(MEM_stage_inst_dmem_ram_2736), .A2(MEM_stage_inst_dmem_n18892), .ZN(MEM_stage_inst_dmem_n18895) );
NAND2_X1 MEM_stage_inst_dmem_U17762 ( .A1(MEM_stage_inst_dmem_n18891), .A2(MEM_stage_inst_dmem_n18890), .ZN(MEM_stage_inst_dmem_n9964) );
NAND2_X1 MEM_stage_inst_dmem_U17761 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n18893), .ZN(MEM_stage_inst_dmem_n18890) );
NAND2_X1 MEM_stage_inst_dmem_U17760 ( .A1(MEM_stage_inst_dmem_ram_2737), .A2(MEM_stage_inst_dmem_n18892), .ZN(MEM_stage_inst_dmem_n18891) );
NAND2_X1 MEM_stage_inst_dmem_U17759 ( .A1(MEM_stage_inst_dmem_n18889), .A2(MEM_stage_inst_dmem_n18888), .ZN(MEM_stage_inst_dmem_n9965) );
NAND2_X1 MEM_stage_inst_dmem_U17758 ( .A1(MEM_stage_inst_dmem_n18887), .A2(MEM_stage_inst_dmem_n18893), .ZN(MEM_stage_inst_dmem_n18888) );
NAND2_X1 MEM_stage_inst_dmem_U17757 ( .A1(MEM_stage_inst_dmem_ram_2738), .A2(MEM_stage_inst_dmem_n18892), .ZN(MEM_stage_inst_dmem_n18889) );
NAND2_X1 MEM_stage_inst_dmem_U17756 ( .A1(MEM_stage_inst_dmem_n18886), .A2(MEM_stage_inst_dmem_n18885), .ZN(MEM_stage_inst_dmem_n9966) );
NAND2_X1 MEM_stage_inst_dmem_U17755 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n18893), .ZN(MEM_stage_inst_dmem_n18885) );
NAND2_X1 MEM_stage_inst_dmem_U17754 ( .A1(MEM_stage_inst_dmem_ram_2739), .A2(MEM_stage_inst_dmem_n18892), .ZN(MEM_stage_inst_dmem_n18886) );
NAND2_X1 MEM_stage_inst_dmem_U17753 ( .A1(MEM_stage_inst_dmem_n18884), .A2(MEM_stage_inst_dmem_n18883), .ZN(MEM_stage_inst_dmem_n9967) );
NAND2_X1 MEM_stage_inst_dmem_U17752 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n18893), .ZN(MEM_stage_inst_dmem_n18883) );
NAND2_X1 MEM_stage_inst_dmem_U17751 ( .A1(MEM_stage_inst_dmem_ram_2740), .A2(MEM_stage_inst_dmem_n18892), .ZN(MEM_stage_inst_dmem_n18884) );
NAND2_X1 MEM_stage_inst_dmem_U17750 ( .A1(MEM_stage_inst_dmem_n18882), .A2(MEM_stage_inst_dmem_n18881), .ZN(MEM_stage_inst_dmem_n9968) );
NAND2_X1 MEM_stage_inst_dmem_U17749 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n18893), .ZN(MEM_stage_inst_dmem_n18881) );
NAND2_X1 MEM_stage_inst_dmem_U17748 ( .A1(MEM_stage_inst_dmem_ram_2741), .A2(MEM_stage_inst_dmem_n18892), .ZN(MEM_stage_inst_dmem_n18882) );
NAND2_X1 MEM_stage_inst_dmem_U17747 ( .A1(MEM_stage_inst_dmem_n18880), .A2(MEM_stage_inst_dmem_n18879), .ZN(MEM_stage_inst_dmem_n9969) );
NAND2_X1 MEM_stage_inst_dmem_U17746 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n18893), .ZN(MEM_stage_inst_dmem_n18879) );
NAND2_X1 MEM_stage_inst_dmem_U17745 ( .A1(MEM_stage_inst_dmem_ram_2742), .A2(MEM_stage_inst_dmem_n18892), .ZN(MEM_stage_inst_dmem_n18880) );
NAND2_X1 MEM_stage_inst_dmem_U17744 ( .A1(MEM_stage_inst_dmem_n18877), .A2(MEM_stage_inst_dmem_n18876), .ZN(MEM_stage_inst_dmem_n9970) );
NAND2_X1 MEM_stage_inst_dmem_U17743 ( .A1(MEM_stage_inst_dmem_n18875), .A2(MEM_stage_inst_dmem_n18893), .ZN(MEM_stage_inst_dmem_n18876) );
NAND2_X1 MEM_stage_inst_dmem_U17742 ( .A1(MEM_stage_inst_dmem_ram_2743), .A2(MEM_stage_inst_dmem_n18892), .ZN(MEM_stage_inst_dmem_n18877) );
NAND2_X1 MEM_stage_inst_dmem_U17741 ( .A1(MEM_stage_inst_dmem_n18874), .A2(MEM_stage_inst_dmem_n18873), .ZN(MEM_stage_inst_dmem_n9971) );
NAND2_X1 MEM_stage_inst_dmem_U17740 ( .A1(MEM_stage_inst_dmem_n111), .A2(MEM_stage_inst_dmem_n18893), .ZN(MEM_stage_inst_dmem_n18873) );
NAND2_X1 MEM_stage_inst_dmem_U17739 ( .A1(MEM_stage_inst_dmem_ram_2744), .A2(MEM_stage_inst_dmem_n18892), .ZN(MEM_stage_inst_dmem_n18874) );
NAND2_X1 MEM_stage_inst_dmem_U17738 ( .A1(MEM_stage_inst_dmem_n18871), .A2(MEM_stage_inst_dmem_n18870), .ZN(MEM_stage_inst_dmem_n9972) );
NAND2_X1 MEM_stage_inst_dmem_U17737 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n18893), .ZN(MEM_stage_inst_dmem_n18870) );
NAND2_X1 MEM_stage_inst_dmem_U17736 ( .A1(MEM_stage_inst_dmem_ram_2745), .A2(MEM_stage_inst_dmem_n18892), .ZN(MEM_stage_inst_dmem_n18871) );
NAND2_X1 MEM_stage_inst_dmem_U17735 ( .A1(MEM_stage_inst_dmem_n18869), .A2(MEM_stage_inst_dmem_n18868), .ZN(MEM_stage_inst_dmem_n9973) );
NAND2_X1 MEM_stage_inst_dmem_U17734 ( .A1(MEM_stage_inst_dmem_n18867), .A2(MEM_stage_inst_dmem_n18893), .ZN(MEM_stage_inst_dmem_n18868) );
NAND2_X1 MEM_stage_inst_dmem_U17733 ( .A1(MEM_stage_inst_dmem_ram_2746), .A2(MEM_stage_inst_dmem_n18892), .ZN(MEM_stage_inst_dmem_n18869) );
NAND2_X1 MEM_stage_inst_dmem_U17732 ( .A1(MEM_stage_inst_dmem_n18866), .A2(MEM_stage_inst_dmem_n18865), .ZN(MEM_stage_inst_dmem_n9974) );
NAND2_X1 MEM_stage_inst_dmem_U17731 ( .A1(MEM_stage_inst_dmem_n18864), .A2(MEM_stage_inst_dmem_n18893), .ZN(MEM_stage_inst_dmem_n18865) );
NAND2_X1 MEM_stage_inst_dmem_U17730 ( .A1(MEM_stage_inst_dmem_ram_2747), .A2(MEM_stage_inst_dmem_n18892), .ZN(MEM_stage_inst_dmem_n18866) );
NAND2_X1 MEM_stage_inst_dmem_U17729 ( .A1(MEM_stage_inst_dmem_n18863), .A2(MEM_stage_inst_dmem_n18862), .ZN(MEM_stage_inst_dmem_n9975) );
NAND2_X1 MEM_stage_inst_dmem_U17728 ( .A1(MEM_stage_inst_dmem_n18861), .A2(MEM_stage_inst_dmem_n18893), .ZN(MEM_stage_inst_dmem_n18862) );
NAND2_X1 MEM_stage_inst_dmem_U17727 ( .A1(MEM_stage_inst_dmem_ram_2748), .A2(MEM_stage_inst_dmem_n18892), .ZN(MEM_stage_inst_dmem_n18863) );
NAND2_X1 MEM_stage_inst_dmem_U17726 ( .A1(MEM_stage_inst_dmem_n18860), .A2(MEM_stage_inst_dmem_n18859), .ZN(MEM_stage_inst_dmem_n9976) );
NAND2_X1 MEM_stage_inst_dmem_U17725 ( .A1(EX_pipeline_reg_out_18), .A2(MEM_stage_inst_dmem_n18893), .ZN(MEM_stage_inst_dmem_n18859) );
NAND2_X1 MEM_stage_inst_dmem_U17724 ( .A1(MEM_stage_inst_dmem_ram_2749), .A2(MEM_stage_inst_dmem_n18892), .ZN(MEM_stage_inst_dmem_n18860) );
NAND2_X1 MEM_stage_inst_dmem_U17723 ( .A1(MEM_stage_inst_dmem_n18858), .A2(MEM_stage_inst_dmem_n18857), .ZN(MEM_stage_inst_dmem_n9977) );
NAND2_X1 MEM_stage_inst_dmem_U17722 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n18893), .ZN(MEM_stage_inst_dmem_n18857) );
NAND2_X1 MEM_stage_inst_dmem_U17721 ( .A1(MEM_stage_inst_dmem_ram_2750), .A2(MEM_stage_inst_dmem_n18892), .ZN(MEM_stage_inst_dmem_n18858) );
NAND2_X1 MEM_stage_inst_dmem_U17720 ( .A1(MEM_stage_inst_dmem_n18856), .A2(MEM_stage_inst_dmem_n18855), .ZN(MEM_stage_inst_dmem_n9978) );
NAND2_X1 MEM_stage_inst_dmem_U17719 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n18893), .ZN(MEM_stage_inst_dmem_n18855) );
INV_X1 MEM_stage_inst_dmem_U17718 ( .A(MEM_stage_inst_dmem_n18892), .ZN(MEM_stage_inst_dmem_n18893) );
NAND2_X1 MEM_stage_inst_dmem_U17717 ( .A1(MEM_stage_inst_dmem_ram_2751), .A2(MEM_stage_inst_dmem_n18892), .ZN(MEM_stage_inst_dmem_n18856) );
NAND2_X1 MEM_stage_inst_dmem_U17716 ( .A1(MEM_stage_inst_dmem_n21074), .A2(MEM_stage_inst_dmem_n19236), .ZN(MEM_stage_inst_dmem_n18892) );
NAND2_X1 MEM_stage_inst_dmem_U17715 ( .A1(MEM_stage_inst_dmem_n18854), .A2(MEM_stage_inst_dmem_n18853), .ZN(MEM_stage_inst_dmem_n9979) );
NAND2_X1 MEM_stage_inst_dmem_U17714 ( .A1(MEM_stage_inst_dmem_n19275), .A2(MEM_stage_inst_dmem_n18852), .ZN(MEM_stage_inst_dmem_n18853) );
NAND2_X1 MEM_stage_inst_dmem_U17713 ( .A1(MEM_stage_inst_dmem_ram_2752), .A2(MEM_stage_inst_dmem_n18851), .ZN(MEM_stage_inst_dmem_n18854) );
NAND2_X1 MEM_stage_inst_dmem_U17712 ( .A1(MEM_stage_inst_dmem_n18850), .A2(MEM_stage_inst_dmem_n18849), .ZN(MEM_stage_inst_dmem_n9980) );
NAND2_X1 MEM_stage_inst_dmem_U17711 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n18852), .ZN(MEM_stage_inst_dmem_n18849) );
NAND2_X1 MEM_stage_inst_dmem_U17710 ( .A1(MEM_stage_inst_dmem_ram_2753), .A2(MEM_stage_inst_dmem_n18851), .ZN(MEM_stage_inst_dmem_n18850) );
NAND2_X1 MEM_stage_inst_dmem_U17709 ( .A1(MEM_stage_inst_dmem_n18848), .A2(MEM_stage_inst_dmem_n18847), .ZN(MEM_stage_inst_dmem_n9981) );
NAND2_X1 MEM_stage_inst_dmem_U17708 ( .A1(EX_pipeline_reg_out_7), .A2(MEM_stage_inst_dmem_n18852), .ZN(MEM_stage_inst_dmem_n18847) );
NAND2_X1 MEM_stage_inst_dmem_U17707 ( .A1(MEM_stage_inst_dmem_ram_2754), .A2(MEM_stage_inst_dmem_n18851), .ZN(MEM_stage_inst_dmem_n18848) );
NAND2_X1 MEM_stage_inst_dmem_U17706 ( .A1(MEM_stage_inst_dmem_n18846), .A2(MEM_stage_inst_dmem_n18845), .ZN(MEM_stage_inst_dmem_n9982) );
NAND2_X1 MEM_stage_inst_dmem_U17705 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n18852), .ZN(MEM_stage_inst_dmem_n18845) );
NAND2_X1 MEM_stage_inst_dmem_U17704 ( .A1(MEM_stage_inst_dmem_ram_2755), .A2(MEM_stage_inst_dmem_n18851), .ZN(MEM_stage_inst_dmem_n18846) );
NAND2_X1 MEM_stage_inst_dmem_U17703 ( .A1(MEM_stage_inst_dmem_n18844), .A2(MEM_stage_inst_dmem_n18843), .ZN(MEM_stage_inst_dmem_n9983) );
NAND2_X1 MEM_stage_inst_dmem_U17702 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n18852), .ZN(MEM_stage_inst_dmem_n18843) );
NAND2_X1 MEM_stage_inst_dmem_U17701 ( .A1(MEM_stage_inst_dmem_ram_2756), .A2(MEM_stage_inst_dmem_n18851), .ZN(MEM_stage_inst_dmem_n18844) );
NAND2_X1 MEM_stage_inst_dmem_U17700 ( .A1(MEM_stage_inst_dmem_n18842), .A2(MEM_stage_inst_dmem_n18841), .ZN(MEM_stage_inst_dmem_n9984) );
NAND2_X1 MEM_stage_inst_dmem_U17699 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n18852), .ZN(MEM_stage_inst_dmem_n18841) );
NAND2_X1 MEM_stage_inst_dmem_U17698 ( .A1(MEM_stage_inst_dmem_ram_2757), .A2(MEM_stage_inst_dmem_n18851), .ZN(MEM_stage_inst_dmem_n18842) );
NAND2_X1 MEM_stage_inst_dmem_U17697 ( .A1(MEM_stage_inst_dmem_n18840), .A2(MEM_stage_inst_dmem_n18839), .ZN(MEM_stage_inst_dmem_n9985) );
NAND2_X1 MEM_stage_inst_dmem_U17696 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n18852), .ZN(MEM_stage_inst_dmem_n18839) );
NAND2_X1 MEM_stage_inst_dmem_U17695 ( .A1(MEM_stage_inst_dmem_ram_2758), .A2(MEM_stage_inst_dmem_n18851), .ZN(MEM_stage_inst_dmem_n18840) );
NAND2_X1 MEM_stage_inst_dmem_U17694 ( .A1(MEM_stage_inst_dmem_n18838), .A2(MEM_stage_inst_dmem_n18837), .ZN(MEM_stage_inst_dmem_n9986) );
NAND2_X1 MEM_stage_inst_dmem_U17693 ( .A1(MEM_stage_inst_dmem_n13886), .A2(MEM_stage_inst_dmem_n18852), .ZN(MEM_stage_inst_dmem_n18837) );
NAND2_X1 MEM_stage_inst_dmem_U17692 ( .A1(MEM_stage_inst_dmem_ram_2759), .A2(MEM_stage_inst_dmem_n18851), .ZN(MEM_stage_inst_dmem_n18838) );
NAND2_X1 MEM_stage_inst_dmem_U17691 ( .A1(MEM_stage_inst_dmem_n18836), .A2(MEM_stage_inst_dmem_n18835), .ZN(MEM_stage_inst_dmem_n9987) );
NAND2_X1 MEM_stage_inst_dmem_U17690 ( .A1(MEM_stage_inst_dmem_n20527), .A2(MEM_stage_inst_dmem_n18852), .ZN(MEM_stage_inst_dmem_n18835) );
NAND2_X1 MEM_stage_inst_dmem_U17689 ( .A1(MEM_stage_inst_dmem_ram_2760), .A2(MEM_stage_inst_dmem_n18851), .ZN(MEM_stage_inst_dmem_n18836) );
NAND2_X1 MEM_stage_inst_dmem_U17688 ( .A1(MEM_stage_inst_dmem_n18834), .A2(MEM_stage_inst_dmem_n18833), .ZN(MEM_stage_inst_dmem_n9988) );
NAND2_X1 MEM_stage_inst_dmem_U17687 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n18852), .ZN(MEM_stage_inst_dmem_n18833) );
NAND2_X1 MEM_stage_inst_dmem_U17686 ( .A1(MEM_stage_inst_dmem_ram_2761), .A2(MEM_stage_inst_dmem_n18851), .ZN(MEM_stage_inst_dmem_n18834) );
NAND2_X1 MEM_stage_inst_dmem_U17685 ( .A1(MEM_stage_inst_dmem_n18832), .A2(MEM_stage_inst_dmem_n18831), .ZN(MEM_stage_inst_dmem_n9989) );
NAND2_X1 MEM_stage_inst_dmem_U17684 ( .A1(EX_pipeline_reg_out_15), .A2(MEM_stage_inst_dmem_n18852), .ZN(MEM_stage_inst_dmem_n18831) );
NAND2_X1 MEM_stage_inst_dmem_U17683 ( .A1(MEM_stage_inst_dmem_ram_2762), .A2(MEM_stage_inst_dmem_n18851), .ZN(MEM_stage_inst_dmem_n18832) );
NAND2_X1 MEM_stage_inst_dmem_U17682 ( .A1(MEM_stage_inst_dmem_n18830), .A2(MEM_stage_inst_dmem_n18829), .ZN(MEM_stage_inst_dmem_n9990) );
NAND2_X1 MEM_stage_inst_dmem_U17681 ( .A1(MEM_stage_inst_dmem_n14705), .A2(MEM_stage_inst_dmem_n18852), .ZN(MEM_stage_inst_dmem_n18829) );
NAND2_X1 MEM_stage_inst_dmem_U17680 ( .A1(MEM_stage_inst_dmem_ram_2763), .A2(MEM_stage_inst_dmem_n18851), .ZN(MEM_stage_inst_dmem_n18830) );
NAND2_X1 MEM_stage_inst_dmem_U17679 ( .A1(MEM_stage_inst_dmem_n18828), .A2(MEM_stage_inst_dmem_n18827), .ZN(MEM_stage_inst_dmem_n9991) );
NAND2_X1 MEM_stage_inst_dmem_U17678 ( .A1(MEM_stage_inst_dmem_n14702), .A2(MEM_stage_inst_dmem_n18852), .ZN(MEM_stage_inst_dmem_n18827) );
NAND2_X1 MEM_stage_inst_dmem_U17677 ( .A1(MEM_stage_inst_dmem_ram_2764), .A2(MEM_stage_inst_dmem_n18851), .ZN(MEM_stage_inst_dmem_n18828) );
NAND2_X1 MEM_stage_inst_dmem_U17676 ( .A1(MEM_stage_inst_dmem_n18826), .A2(MEM_stage_inst_dmem_n18825), .ZN(MEM_stage_inst_dmem_n9992) );
NAND2_X1 MEM_stage_inst_dmem_U17675 ( .A1(MEM_stage_inst_dmem_n19242), .A2(MEM_stage_inst_dmem_n18852), .ZN(MEM_stage_inst_dmem_n18825) );
NAND2_X1 MEM_stage_inst_dmem_U17674 ( .A1(MEM_stage_inst_dmem_ram_2765), .A2(MEM_stage_inst_dmem_n18851), .ZN(MEM_stage_inst_dmem_n18826) );
NAND2_X1 MEM_stage_inst_dmem_U17673 ( .A1(MEM_stage_inst_dmem_n18824), .A2(MEM_stage_inst_dmem_n18823), .ZN(MEM_stage_inst_dmem_n9993) );
NAND2_X1 MEM_stage_inst_dmem_U17672 ( .A1(MEM_stage_inst_dmem_n115), .A2(MEM_stage_inst_dmem_n18852), .ZN(MEM_stage_inst_dmem_n18823) );
NAND2_X1 MEM_stage_inst_dmem_U17671 ( .A1(MEM_stage_inst_dmem_ram_2766), .A2(MEM_stage_inst_dmem_n18851), .ZN(MEM_stage_inst_dmem_n18824) );
NAND2_X1 MEM_stage_inst_dmem_U17670 ( .A1(MEM_stage_inst_dmem_n18822), .A2(MEM_stage_inst_dmem_n18821), .ZN(MEM_stage_inst_dmem_n9994) );
NAND2_X1 MEM_stage_inst_dmem_U17669 ( .A1(EX_pipeline_reg_out_20), .A2(MEM_stage_inst_dmem_n18852), .ZN(MEM_stage_inst_dmem_n18821) );
NAND2_X1 MEM_stage_inst_dmem_U17668 ( .A1(MEM_stage_inst_dmem_ram_2767), .A2(MEM_stage_inst_dmem_n18851), .ZN(MEM_stage_inst_dmem_n18822) );
NAND2_X1 MEM_stage_inst_dmem_U17667 ( .A1(MEM_stage_inst_dmem_n21039), .A2(MEM_stage_inst_dmem_n19236), .ZN(MEM_stage_inst_dmem_n18851) );
NAND2_X1 MEM_stage_inst_dmem_U17666 ( .A1(MEM_stage_inst_dmem_n18820), .A2(MEM_stage_inst_dmem_n18819), .ZN(MEM_stage_inst_dmem_n9995) );
NAND2_X1 MEM_stage_inst_dmem_U17665 ( .A1(MEM_stage_inst_dmem_n19275), .A2(MEM_stage_inst_dmem_n18818), .ZN(MEM_stage_inst_dmem_n18819) );
NAND2_X1 MEM_stage_inst_dmem_U17664 ( .A1(MEM_stage_inst_dmem_ram_2768), .A2(MEM_stage_inst_dmem_n18817), .ZN(MEM_stage_inst_dmem_n18820) );
NAND2_X1 MEM_stage_inst_dmem_U17663 ( .A1(MEM_stage_inst_dmem_n18816), .A2(MEM_stage_inst_dmem_n18815), .ZN(MEM_stage_inst_dmem_n9996) );
NAND2_X1 MEM_stage_inst_dmem_U17662 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n18818), .ZN(MEM_stage_inst_dmem_n18815) );
NAND2_X1 MEM_stage_inst_dmem_U17661 ( .A1(MEM_stage_inst_dmem_ram_2769), .A2(MEM_stage_inst_dmem_n18817), .ZN(MEM_stage_inst_dmem_n18816) );
NAND2_X1 MEM_stage_inst_dmem_U17660 ( .A1(MEM_stage_inst_dmem_n18814), .A2(MEM_stage_inst_dmem_n18813), .ZN(MEM_stage_inst_dmem_n9997) );
NAND2_X1 MEM_stage_inst_dmem_U17659 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n18818), .ZN(MEM_stage_inst_dmem_n18813) );
NAND2_X1 MEM_stage_inst_dmem_U17658 ( .A1(MEM_stage_inst_dmem_ram_2770), .A2(MEM_stage_inst_dmem_n18817), .ZN(MEM_stage_inst_dmem_n18814) );
NAND2_X1 MEM_stage_inst_dmem_U17657 ( .A1(MEM_stage_inst_dmem_n18812), .A2(MEM_stage_inst_dmem_n18811), .ZN(MEM_stage_inst_dmem_n9998) );
NAND2_X1 MEM_stage_inst_dmem_U17656 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n18818), .ZN(MEM_stage_inst_dmem_n18811) );
NAND2_X1 MEM_stage_inst_dmem_U17655 ( .A1(MEM_stage_inst_dmem_ram_2771), .A2(MEM_stage_inst_dmem_n18817), .ZN(MEM_stage_inst_dmem_n18812) );
NAND2_X1 MEM_stage_inst_dmem_U17654 ( .A1(MEM_stage_inst_dmem_n18810), .A2(MEM_stage_inst_dmem_n18809), .ZN(MEM_stage_inst_dmem_n9999) );
NAND2_X1 MEM_stage_inst_dmem_U17653 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n18818), .ZN(MEM_stage_inst_dmem_n18809) );
NAND2_X1 MEM_stage_inst_dmem_U17652 ( .A1(MEM_stage_inst_dmem_ram_2772), .A2(MEM_stage_inst_dmem_n18817), .ZN(MEM_stage_inst_dmem_n18810) );
NAND2_X1 MEM_stage_inst_dmem_U17651 ( .A1(MEM_stage_inst_dmem_n18808), .A2(MEM_stage_inst_dmem_n18807), .ZN(MEM_stage_inst_dmem_n10000) );
NAND2_X1 MEM_stage_inst_dmem_U17650 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n18818), .ZN(MEM_stage_inst_dmem_n18807) );
NAND2_X1 MEM_stage_inst_dmem_U17649 ( .A1(MEM_stage_inst_dmem_ram_2773), .A2(MEM_stage_inst_dmem_n18817), .ZN(MEM_stage_inst_dmem_n18808) );
NAND2_X1 MEM_stage_inst_dmem_U17648 ( .A1(MEM_stage_inst_dmem_n18806), .A2(MEM_stage_inst_dmem_n18805), .ZN(MEM_stage_inst_dmem_n10001) );
NAND2_X1 MEM_stage_inst_dmem_U17647 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n18818), .ZN(MEM_stage_inst_dmem_n18805) );
NAND2_X1 MEM_stage_inst_dmem_U17646 ( .A1(MEM_stage_inst_dmem_ram_2774), .A2(MEM_stage_inst_dmem_n18817), .ZN(MEM_stage_inst_dmem_n18806) );
NAND2_X1 MEM_stage_inst_dmem_U17645 ( .A1(MEM_stage_inst_dmem_n18804), .A2(MEM_stage_inst_dmem_n18803), .ZN(MEM_stage_inst_dmem_n10002) );
NAND2_X1 MEM_stage_inst_dmem_U17644 ( .A1(MEM_stage_inst_dmem_n20530), .A2(MEM_stage_inst_dmem_n18818), .ZN(MEM_stage_inst_dmem_n18803) );
NAND2_X1 MEM_stage_inst_dmem_U17643 ( .A1(MEM_stage_inst_dmem_ram_2775), .A2(MEM_stage_inst_dmem_n18817), .ZN(MEM_stage_inst_dmem_n18804) );
NAND2_X1 MEM_stage_inst_dmem_U17642 ( .A1(MEM_stage_inst_dmem_n18802), .A2(MEM_stage_inst_dmem_n18801), .ZN(MEM_stage_inst_dmem_n10003) );
NAND2_X1 MEM_stage_inst_dmem_U17641 ( .A1(MEM_stage_inst_dmem_n13883), .A2(MEM_stage_inst_dmem_n18818), .ZN(MEM_stage_inst_dmem_n18801) );
NAND2_X1 MEM_stage_inst_dmem_U17640 ( .A1(MEM_stage_inst_dmem_ram_2776), .A2(MEM_stage_inst_dmem_n18817), .ZN(MEM_stage_inst_dmem_n18802) );
NAND2_X1 MEM_stage_inst_dmem_U17639 ( .A1(MEM_stage_inst_dmem_n18800), .A2(MEM_stage_inst_dmem_n18799), .ZN(MEM_stage_inst_dmem_n10004) );
NAND2_X1 MEM_stage_inst_dmem_U17638 ( .A1(MEM_stage_inst_dmem_n19251), .A2(MEM_stage_inst_dmem_n18818), .ZN(MEM_stage_inst_dmem_n18799) );
NAND2_X1 MEM_stage_inst_dmem_U17637 ( .A1(MEM_stage_inst_dmem_ram_2777), .A2(MEM_stage_inst_dmem_n18817), .ZN(MEM_stage_inst_dmem_n18800) );
NAND2_X1 MEM_stage_inst_dmem_U17636 ( .A1(MEM_stage_inst_dmem_n18798), .A2(MEM_stage_inst_dmem_n18797), .ZN(MEM_stage_inst_dmem_n10005) );
NAND2_X1 MEM_stage_inst_dmem_U17635 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n18818), .ZN(MEM_stage_inst_dmem_n18797) );
NAND2_X1 MEM_stage_inst_dmem_U17634 ( .A1(MEM_stage_inst_dmem_ram_2778), .A2(MEM_stage_inst_dmem_n18817), .ZN(MEM_stage_inst_dmem_n18798) );
NAND2_X1 MEM_stage_inst_dmem_U17633 ( .A1(MEM_stage_inst_dmem_n18796), .A2(MEM_stage_inst_dmem_n18795), .ZN(MEM_stage_inst_dmem_n10006) );
NAND2_X1 MEM_stage_inst_dmem_U17632 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n18818), .ZN(MEM_stage_inst_dmem_n18795) );
NAND2_X1 MEM_stage_inst_dmem_U17631 ( .A1(MEM_stage_inst_dmem_ram_2779), .A2(MEM_stage_inst_dmem_n18817), .ZN(MEM_stage_inst_dmem_n18796) );
NAND2_X1 MEM_stage_inst_dmem_U17630 ( .A1(MEM_stage_inst_dmem_n18794), .A2(MEM_stage_inst_dmem_n18793), .ZN(MEM_stage_inst_dmem_n10007) );
NAND2_X1 MEM_stage_inst_dmem_U17629 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n18818), .ZN(MEM_stage_inst_dmem_n18793) );
NAND2_X1 MEM_stage_inst_dmem_U17628 ( .A1(MEM_stage_inst_dmem_ram_2780), .A2(MEM_stage_inst_dmem_n18817), .ZN(MEM_stage_inst_dmem_n18794) );
NAND2_X1 MEM_stage_inst_dmem_U17627 ( .A1(MEM_stage_inst_dmem_n18792), .A2(MEM_stage_inst_dmem_n18791), .ZN(MEM_stage_inst_dmem_n10008) );
NAND2_X1 MEM_stage_inst_dmem_U17626 ( .A1(MEM_stage_inst_dmem_n19242), .A2(MEM_stage_inst_dmem_n18818), .ZN(MEM_stage_inst_dmem_n18791) );
NAND2_X1 MEM_stage_inst_dmem_U17625 ( .A1(MEM_stage_inst_dmem_ram_2781), .A2(MEM_stage_inst_dmem_n18817), .ZN(MEM_stage_inst_dmem_n18792) );
NAND2_X1 MEM_stage_inst_dmem_U17624 ( .A1(MEM_stage_inst_dmem_n18790), .A2(MEM_stage_inst_dmem_n18789), .ZN(MEM_stage_inst_dmem_n10009) );
NAND2_X1 MEM_stage_inst_dmem_U17623 ( .A1(MEM_stage_inst_dmem_n115), .A2(MEM_stage_inst_dmem_n18818), .ZN(MEM_stage_inst_dmem_n18789) );
NAND2_X1 MEM_stage_inst_dmem_U17622 ( .A1(MEM_stage_inst_dmem_ram_2782), .A2(MEM_stage_inst_dmem_n18817), .ZN(MEM_stage_inst_dmem_n18790) );
NAND2_X1 MEM_stage_inst_dmem_U17621 ( .A1(MEM_stage_inst_dmem_n18788), .A2(MEM_stage_inst_dmem_n18787), .ZN(MEM_stage_inst_dmem_n10010) );
NAND2_X1 MEM_stage_inst_dmem_U17620 ( .A1(MEM_stage_inst_dmem_n20506), .A2(MEM_stage_inst_dmem_n18818), .ZN(MEM_stage_inst_dmem_n18787) );
INV_X1 MEM_stage_inst_dmem_U17619 ( .A(MEM_stage_inst_dmem_n18817), .ZN(MEM_stage_inst_dmem_n18818) );
NAND2_X1 MEM_stage_inst_dmem_U17618 ( .A1(MEM_stage_inst_dmem_ram_2783), .A2(MEM_stage_inst_dmem_n18817), .ZN(MEM_stage_inst_dmem_n18788) );
NAND2_X1 MEM_stage_inst_dmem_U17617 ( .A1(MEM_stage_inst_dmem_n21004), .A2(MEM_stage_inst_dmem_n19236), .ZN(MEM_stage_inst_dmem_n18817) );
NAND2_X1 MEM_stage_inst_dmem_U17616 ( .A1(MEM_stage_inst_dmem_n18786), .A2(MEM_stage_inst_dmem_n18785), .ZN(MEM_stage_inst_dmem_n10011) );
NAND2_X1 MEM_stage_inst_dmem_U17615 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n18784), .ZN(MEM_stage_inst_dmem_n18785) );
NAND2_X1 MEM_stage_inst_dmem_U17614 ( .A1(MEM_stage_inst_dmem_ram_2784), .A2(MEM_stage_inst_dmem_n18783), .ZN(MEM_stage_inst_dmem_n18786) );
NAND2_X1 MEM_stage_inst_dmem_U17613 ( .A1(MEM_stage_inst_dmem_n18782), .A2(MEM_stage_inst_dmem_n18781), .ZN(MEM_stage_inst_dmem_n10012) );
NAND2_X1 MEM_stage_inst_dmem_U17612 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n18784), .ZN(MEM_stage_inst_dmem_n18781) );
NAND2_X1 MEM_stage_inst_dmem_U17611 ( .A1(MEM_stage_inst_dmem_ram_2785), .A2(MEM_stage_inst_dmem_n18783), .ZN(MEM_stage_inst_dmem_n18782) );
NAND2_X1 MEM_stage_inst_dmem_U17610 ( .A1(MEM_stage_inst_dmem_n18780), .A2(MEM_stage_inst_dmem_n18779), .ZN(MEM_stage_inst_dmem_n10013) );
NAND2_X1 MEM_stage_inst_dmem_U17609 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n18784), .ZN(MEM_stage_inst_dmem_n18779) );
NAND2_X1 MEM_stage_inst_dmem_U17608 ( .A1(MEM_stage_inst_dmem_ram_2786), .A2(MEM_stage_inst_dmem_n18783), .ZN(MEM_stage_inst_dmem_n18780) );
NAND2_X1 MEM_stage_inst_dmem_U17607 ( .A1(MEM_stage_inst_dmem_n18778), .A2(MEM_stage_inst_dmem_n18777), .ZN(MEM_stage_inst_dmem_n10014) );
NAND2_X1 MEM_stage_inst_dmem_U17606 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n18784), .ZN(MEM_stage_inst_dmem_n18777) );
NAND2_X1 MEM_stage_inst_dmem_U17605 ( .A1(MEM_stage_inst_dmem_ram_2787), .A2(MEM_stage_inst_dmem_n18783), .ZN(MEM_stage_inst_dmem_n18778) );
NAND2_X1 MEM_stage_inst_dmem_U17604 ( .A1(MEM_stage_inst_dmem_n18776), .A2(MEM_stage_inst_dmem_n18775), .ZN(MEM_stage_inst_dmem_n10015) );
NAND2_X1 MEM_stage_inst_dmem_U17603 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n18784), .ZN(MEM_stage_inst_dmem_n18775) );
NAND2_X1 MEM_stage_inst_dmem_U17602 ( .A1(MEM_stage_inst_dmem_ram_2788), .A2(MEM_stage_inst_dmem_n18783), .ZN(MEM_stage_inst_dmem_n18776) );
NAND2_X1 MEM_stage_inst_dmem_U17601 ( .A1(MEM_stage_inst_dmem_n18774), .A2(MEM_stage_inst_dmem_n18773), .ZN(MEM_stage_inst_dmem_n10016) );
NAND2_X1 MEM_stage_inst_dmem_U17600 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n18784), .ZN(MEM_stage_inst_dmem_n18773) );
NAND2_X1 MEM_stage_inst_dmem_U17599 ( .A1(MEM_stage_inst_dmem_ram_2789), .A2(MEM_stage_inst_dmem_n18783), .ZN(MEM_stage_inst_dmem_n18774) );
NAND2_X1 MEM_stage_inst_dmem_U17598 ( .A1(MEM_stage_inst_dmem_n18772), .A2(MEM_stage_inst_dmem_n18771), .ZN(MEM_stage_inst_dmem_n10017) );
NAND2_X1 MEM_stage_inst_dmem_U17597 ( .A1(MEM_stage_inst_dmem_n21340), .A2(MEM_stage_inst_dmem_n18784), .ZN(MEM_stage_inst_dmem_n18771) );
NAND2_X1 MEM_stage_inst_dmem_U17596 ( .A1(MEM_stage_inst_dmem_ram_2790), .A2(MEM_stage_inst_dmem_n18783), .ZN(MEM_stage_inst_dmem_n18772) );
NAND2_X1 MEM_stage_inst_dmem_U17595 ( .A1(MEM_stage_inst_dmem_n18770), .A2(MEM_stage_inst_dmem_n18769), .ZN(MEM_stage_inst_dmem_n10018) );
NAND2_X1 MEM_stage_inst_dmem_U17594 ( .A1(MEM_stage_inst_dmem_n18), .A2(MEM_stage_inst_dmem_n18784), .ZN(MEM_stage_inst_dmem_n18769) );
NAND2_X1 MEM_stage_inst_dmem_U17593 ( .A1(MEM_stage_inst_dmem_ram_2791), .A2(MEM_stage_inst_dmem_n18783), .ZN(MEM_stage_inst_dmem_n18770) );
NAND2_X1 MEM_stage_inst_dmem_U17592 ( .A1(MEM_stage_inst_dmem_n18768), .A2(MEM_stage_inst_dmem_n18767), .ZN(MEM_stage_inst_dmem_n10019) );
NAND2_X1 MEM_stage_inst_dmem_U17591 ( .A1(MEM_stage_inst_dmem_n21335), .A2(MEM_stage_inst_dmem_n18784), .ZN(MEM_stage_inst_dmem_n18767) );
NAND2_X1 MEM_stage_inst_dmem_U17590 ( .A1(MEM_stage_inst_dmem_ram_2792), .A2(MEM_stage_inst_dmem_n18783), .ZN(MEM_stage_inst_dmem_n18768) );
NAND2_X1 MEM_stage_inst_dmem_U17589 ( .A1(MEM_stage_inst_dmem_n18766), .A2(MEM_stage_inst_dmem_n18765), .ZN(MEM_stage_inst_dmem_n10020) );
NAND2_X1 MEM_stage_inst_dmem_U17588 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n18784), .ZN(MEM_stage_inst_dmem_n18765) );
NAND2_X1 MEM_stage_inst_dmem_U17587 ( .A1(MEM_stage_inst_dmem_ram_2793), .A2(MEM_stage_inst_dmem_n18783), .ZN(MEM_stage_inst_dmem_n18766) );
NAND2_X1 MEM_stage_inst_dmem_U17586 ( .A1(MEM_stage_inst_dmem_n18764), .A2(MEM_stage_inst_dmem_n18763), .ZN(MEM_stage_inst_dmem_n10021) );
NAND2_X1 MEM_stage_inst_dmem_U17585 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n18784), .ZN(MEM_stage_inst_dmem_n18763) );
NAND2_X1 MEM_stage_inst_dmem_U17584 ( .A1(MEM_stage_inst_dmem_ram_2794), .A2(MEM_stage_inst_dmem_n18783), .ZN(MEM_stage_inst_dmem_n18764) );
NAND2_X1 MEM_stage_inst_dmem_U17583 ( .A1(MEM_stage_inst_dmem_n18762), .A2(MEM_stage_inst_dmem_n18761), .ZN(MEM_stage_inst_dmem_n10022) );
NAND2_X1 MEM_stage_inst_dmem_U17582 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n18784), .ZN(MEM_stage_inst_dmem_n18761) );
NAND2_X1 MEM_stage_inst_dmem_U17581 ( .A1(MEM_stage_inst_dmem_ram_2795), .A2(MEM_stage_inst_dmem_n18783), .ZN(MEM_stage_inst_dmem_n18762) );
NAND2_X1 MEM_stage_inst_dmem_U17580 ( .A1(MEM_stage_inst_dmem_n18760), .A2(MEM_stage_inst_dmem_n18759), .ZN(MEM_stage_inst_dmem_n10023) );
NAND2_X1 MEM_stage_inst_dmem_U17579 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n18784), .ZN(MEM_stage_inst_dmem_n18759) );
NAND2_X1 MEM_stage_inst_dmem_U17578 ( .A1(MEM_stage_inst_dmem_ram_2796), .A2(MEM_stage_inst_dmem_n18783), .ZN(MEM_stage_inst_dmem_n18760) );
NAND2_X1 MEM_stage_inst_dmem_U17577 ( .A1(MEM_stage_inst_dmem_n18758), .A2(MEM_stage_inst_dmem_n18757), .ZN(MEM_stage_inst_dmem_n10024) );
NAND2_X1 MEM_stage_inst_dmem_U17576 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n18784), .ZN(MEM_stage_inst_dmem_n18757) );
NAND2_X1 MEM_stage_inst_dmem_U17575 ( .A1(MEM_stage_inst_dmem_ram_2797), .A2(MEM_stage_inst_dmem_n18783), .ZN(MEM_stage_inst_dmem_n18758) );
NAND2_X1 MEM_stage_inst_dmem_U17574 ( .A1(MEM_stage_inst_dmem_n18756), .A2(MEM_stage_inst_dmem_n18755), .ZN(MEM_stage_inst_dmem_n10025) );
NAND2_X1 MEM_stage_inst_dmem_U17573 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n18784), .ZN(MEM_stage_inst_dmem_n18755) );
NAND2_X1 MEM_stage_inst_dmem_U17572 ( .A1(MEM_stage_inst_dmem_ram_2798), .A2(MEM_stage_inst_dmem_n18783), .ZN(MEM_stage_inst_dmem_n18756) );
NAND2_X1 MEM_stage_inst_dmem_U17571 ( .A1(MEM_stage_inst_dmem_n18754), .A2(MEM_stage_inst_dmem_n18753), .ZN(MEM_stage_inst_dmem_n10026) );
NAND2_X1 MEM_stage_inst_dmem_U17570 ( .A1(MEM_stage_inst_dmem_n21320), .A2(MEM_stage_inst_dmem_n18784), .ZN(MEM_stage_inst_dmem_n18753) );
INV_X1 MEM_stage_inst_dmem_U17569 ( .A(MEM_stage_inst_dmem_n18783), .ZN(MEM_stage_inst_dmem_n18784) );
NAND2_X1 MEM_stage_inst_dmem_U17568 ( .A1(MEM_stage_inst_dmem_ram_2799), .A2(MEM_stage_inst_dmem_n18783), .ZN(MEM_stage_inst_dmem_n18754) );
NAND2_X1 MEM_stage_inst_dmem_U17567 ( .A1(MEM_stage_inst_dmem_n20969), .A2(MEM_stage_inst_dmem_n19236), .ZN(MEM_stage_inst_dmem_n18783) );
NAND2_X1 MEM_stage_inst_dmem_U17566 ( .A1(MEM_stage_inst_dmem_n18752), .A2(MEM_stage_inst_dmem_n18751), .ZN(MEM_stage_inst_dmem_n10027) );
NAND2_X1 MEM_stage_inst_dmem_U17565 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n18750), .ZN(MEM_stage_inst_dmem_n18751) );
NAND2_X1 MEM_stage_inst_dmem_U17564 ( .A1(MEM_stage_inst_dmem_ram_2800), .A2(MEM_stage_inst_dmem_n18749), .ZN(MEM_stage_inst_dmem_n18752) );
NAND2_X1 MEM_stage_inst_dmem_U17563 ( .A1(MEM_stage_inst_dmem_n18748), .A2(MEM_stage_inst_dmem_n18747), .ZN(MEM_stage_inst_dmem_n10028) );
NAND2_X1 MEM_stage_inst_dmem_U17562 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n18750), .ZN(MEM_stage_inst_dmem_n18747) );
NAND2_X1 MEM_stage_inst_dmem_U17561 ( .A1(MEM_stage_inst_dmem_ram_2801), .A2(MEM_stage_inst_dmem_n18749), .ZN(MEM_stage_inst_dmem_n18748) );
NAND2_X1 MEM_stage_inst_dmem_U17560 ( .A1(MEM_stage_inst_dmem_n18746), .A2(MEM_stage_inst_dmem_n18745), .ZN(MEM_stage_inst_dmem_n10029) );
NAND2_X1 MEM_stage_inst_dmem_U17559 ( .A1(MEM_stage_inst_dmem_n18887), .A2(MEM_stage_inst_dmem_n18750), .ZN(MEM_stage_inst_dmem_n18745) );
NAND2_X1 MEM_stage_inst_dmem_U17558 ( .A1(MEM_stage_inst_dmem_ram_2802), .A2(MEM_stage_inst_dmem_n18749), .ZN(MEM_stage_inst_dmem_n18746) );
NAND2_X1 MEM_stage_inst_dmem_U17557 ( .A1(MEM_stage_inst_dmem_n18744), .A2(MEM_stage_inst_dmem_n18743), .ZN(MEM_stage_inst_dmem_n10030) );
NAND2_X1 MEM_stage_inst_dmem_U17556 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n18750), .ZN(MEM_stage_inst_dmem_n18743) );
NAND2_X1 MEM_stage_inst_dmem_U17555 ( .A1(MEM_stage_inst_dmem_ram_2803), .A2(MEM_stage_inst_dmem_n18749), .ZN(MEM_stage_inst_dmem_n18744) );
NAND2_X1 MEM_stage_inst_dmem_U17554 ( .A1(MEM_stage_inst_dmem_n18742), .A2(MEM_stage_inst_dmem_n18741), .ZN(MEM_stage_inst_dmem_n10031) );
NAND2_X1 MEM_stage_inst_dmem_U17553 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n18750), .ZN(MEM_stage_inst_dmem_n18741) );
NAND2_X1 MEM_stage_inst_dmem_U17552 ( .A1(MEM_stage_inst_dmem_ram_2804), .A2(MEM_stage_inst_dmem_n18749), .ZN(MEM_stage_inst_dmem_n18742) );
NAND2_X1 MEM_stage_inst_dmem_U17551 ( .A1(MEM_stage_inst_dmem_n18740), .A2(MEM_stage_inst_dmem_n18739), .ZN(MEM_stage_inst_dmem_n10032) );
NAND2_X1 MEM_stage_inst_dmem_U17550 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n18750), .ZN(MEM_stage_inst_dmem_n18739) );
NAND2_X1 MEM_stage_inst_dmem_U17549 ( .A1(MEM_stage_inst_dmem_ram_2805), .A2(MEM_stage_inst_dmem_n18749), .ZN(MEM_stage_inst_dmem_n18740) );
NAND2_X1 MEM_stage_inst_dmem_U17548 ( .A1(MEM_stage_inst_dmem_n18738), .A2(MEM_stage_inst_dmem_n18737), .ZN(MEM_stage_inst_dmem_n10033) );
NAND2_X1 MEM_stage_inst_dmem_U17547 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n18750), .ZN(MEM_stage_inst_dmem_n18737) );
NAND2_X1 MEM_stage_inst_dmem_U17546 ( .A1(MEM_stage_inst_dmem_ram_2806), .A2(MEM_stage_inst_dmem_n18749), .ZN(MEM_stage_inst_dmem_n18738) );
NAND2_X1 MEM_stage_inst_dmem_U17545 ( .A1(MEM_stage_inst_dmem_n18736), .A2(MEM_stage_inst_dmem_n18735), .ZN(MEM_stage_inst_dmem_n10034) );
NAND2_X1 MEM_stage_inst_dmem_U17544 ( .A1(MEM_stage_inst_dmem_n18875), .A2(MEM_stage_inst_dmem_n18750), .ZN(MEM_stage_inst_dmem_n18735) );
NAND2_X1 MEM_stage_inst_dmem_U17543 ( .A1(MEM_stage_inst_dmem_ram_2807), .A2(MEM_stage_inst_dmem_n18749), .ZN(MEM_stage_inst_dmem_n18736) );
NAND2_X1 MEM_stage_inst_dmem_U17542 ( .A1(MEM_stage_inst_dmem_n18734), .A2(MEM_stage_inst_dmem_n18733), .ZN(MEM_stage_inst_dmem_n10035) );
NAND2_X1 MEM_stage_inst_dmem_U17541 ( .A1(MEM_stage_inst_dmem_n111), .A2(MEM_stage_inst_dmem_n18750), .ZN(MEM_stage_inst_dmem_n18733) );
NAND2_X1 MEM_stage_inst_dmem_U17540 ( .A1(MEM_stage_inst_dmem_ram_2808), .A2(MEM_stage_inst_dmem_n18749), .ZN(MEM_stage_inst_dmem_n18734) );
NAND2_X1 MEM_stage_inst_dmem_U17539 ( .A1(MEM_stage_inst_dmem_n18732), .A2(MEM_stage_inst_dmem_n18731), .ZN(MEM_stage_inst_dmem_n10036) );
NAND2_X1 MEM_stage_inst_dmem_U17538 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n18750), .ZN(MEM_stage_inst_dmem_n18731) );
NAND2_X1 MEM_stage_inst_dmem_U17537 ( .A1(MEM_stage_inst_dmem_ram_2809), .A2(MEM_stage_inst_dmem_n18749), .ZN(MEM_stage_inst_dmem_n18732) );
NAND2_X1 MEM_stage_inst_dmem_U17536 ( .A1(MEM_stage_inst_dmem_n18730), .A2(MEM_stage_inst_dmem_n18729), .ZN(MEM_stage_inst_dmem_n10037) );
NAND2_X1 MEM_stage_inst_dmem_U17535 ( .A1(MEM_stage_inst_dmem_n18867), .A2(MEM_stage_inst_dmem_n18750), .ZN(MEM_stage_inst_dmem_n18729) );
NAND2_X1 MEM_stage_inst_dmem_U17534 ( .A1(MEM_stage_inst_dmem_ram_2810), .A2(MEM_stage_inst_dmem_n18749), .ZN(MEM_stage_inst_dmem_n18730) );
NAND2_X1 MEM_stage_inst_dmem_U17533 ( .A1(MEM_stage_inst_dmem_n18728), .A2(MEM_stage_inst_dmem_n18727), .ZN(MEM_stage_inst_dmem_n10038) );
NAND2_X1 MEM_stage_inst_dmem_U17532 ( .A1(MEM_stage_inst_dmem_n18864), .A2(MEM_stage_inst_dmem_n18750), .ZN(MEM_stage_inst_dmem_n18727) );
NAND2_X1 MEM_stage_inst_dmem_U17531 ( .A1(MEM_stage_inst_dmem_ram_2811), .A2(MEM_stage_inst_dmem_n18749), .ZN(MEM_stage_inst_dmem_n18728) );
NAND2_X1 MEM_stage_inst_dmem_U17530 ( .A1(MEM_stage_inst_dmem_n18726), .A2(MEM_stage_inst_dmem_n18725), .ZN(MEM_stage_inst_dmem_n10039) );
NAND2_X1 MEM_stage_inst_dmem_U17529 ( .A1(MEM_stage_inst_dmem_n18861), .A2(MEM_stage_inst_dmem_n18750), .ZN(MEM_stage_inst_dmem_n18725) );
NAND2_X1 MEM_stage_inst_dmem_U17528 ( .A1(MEM_stage_inst_dmem_ram_2812), .A2(MEM_stage_inst_dmem_n18749), .ZN(MEM_stage_inst_dmem_n18726) );
NAND2_X1 MEM_stage_inst_dmem_U17527 ( .A1(MEM_stage_inst_dmem_n18724), .A2(MEM_stage_inst_dmem_n18723), .ZN(MEM_stage_inst_dmem_n10040) );
NAND2_X1 MEM_stage_inst_dmem_U17526 ( .A1(MEM_stage_inst_dmem_n116), .A2(MEM_stage_inst_dmem_n18750), .ZN(MEM_stage_inst_dmem_n18723) );
NAND2_X1 MEM_stage_inst_dmem_U17525 ( .A1(MEM_stage_inst_dmem_ram_2813), .A2(MEM_stage_inst_dmem_n18749), .ZN(MEM_stage_inst_dmem_n18724) );
NAND2_X1 MEM_stage_inst_dmem_U17524 ( .A1(MEM_stage_inst_dmem_n18722), .A2(MEM_stage_inst_dmem_n18721), .ZN(MEM_stage_inst_dmem_n10041) );
NAND2_X1 MEM_stage_inst_dmem_U17523 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n18750), .ZN(MEM_stage_inst_dmem_n18721) );
NAND2_X1 MEM_stage_inst_dmem_U17522 ( .A1(MEM_stage_inst_dmem_ram_2814), .A2(MEM_stage_inst_dmem_n18749), .ZN(MEM_stage_inst_dmem_n18722) );
NAND2_X1 MEM_stage_inst_dmem_U17521 ( .A1(MEM_stage_inst_dmem_n18720), .A2(MEM_stage_inst_dmem_n18719), .ZN(MEM_stage_inst_dmem_n10042) );
NAND2_X1 MEM_stage_inst_dmem_U17520 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n18750), .ZN(MEM_stage_inst_dmem_n18719) );
INV_X1 MEM_stage_inst_dmem_U17519 ( .A(MEM_stage_inst_dmem_n18749), .ZN(MEM_stage_inst_dmem_n18750) );
NAND2_X1 MEM_stage_inst_dmem_U17518 ( .A1(MEM_stage_inst_dmem_ram_2815), .A2(MEM_stage_inst_dmem_n18749), .ZN(MEM_stage_inst_dmem_n18720) );
NAND2_X1 MEM_stage_inst_dmem_U17517 ( .A1(MEM_stage_inst_dmem_n20934), .A2(MEM_stage_inst_dmem_n19236), .ZN(MEM_stage_inst_dmem_n18749) );
NOR2_X2 MEM_stage_inst_dmem_U17516 ( .A1(MEM_stage_inst_dmem_n18718), .A2(MEM_stage_inst_dmem_n20932), .ZN(MEM_stage_inst_dmem_n19236) );
NAND2_X1 MEM_stage_inst_dmem_U17515 ( .A1(MEM_stage_inst_dmem_n18717), .A2(MEM_stage_inst_dmem_n18716), .ZN(MEM_stage_inst_dmem_n10043) );
NAND2_X1 MEM_stage_inst_dmem_U17514 ( .A1(MEM_stage_inst_dmem_n19275), .A2(MEM_stage_inst_dmem_n18715), .ZN(MEM_stage_inst_dmem_n18716) );
NAND2_X1 MEM_stage_inst_dmem_U17513 ( .A1(MEM_stage_inst_dmem_ram_2816), .A2(MEM_stage_inst_dmem_n18714), .ZN(MEM_stage_inst_dmem_n18717) );
NAND2_X1 MEM_stage_inst_dmem_U17512 ( .A1(MEM_stage_inst_dmem_n18713), .A2(MEM_stage_inst_dmem_n18712), .ZN(MEM_stage_inst_dmem_n10044) );
NAND2_X1 MEM_stage_inst_dmem_U17511 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n18715), .ZN(MEM_stage_inst_dmem_n18712) );
NAND2_X1 MEM_stage_inst_dmem_U17510 ( .A1(MEM_stage_inst_dmem_ram_2817), .A2(MEM_stage_inst_dmem_n18714), .ZN(MEM_stage_inst_dmem_n18713) );
NAND2_X1 MEM_stage_inst_dmem_U17509 ( .A1(MEM_stage_inst_dmem_n18711), .A2(MEM_stage_inst_dmem_n18710), .ZN(MEM_stage_inst_dmem_n10045) );
NAND2_X1 MEM_stage_inst_dmem_U17508 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n18715), .ZN(MEM_stage_inst_dmem_n18710) );
NAND2_X1 MEM_stage_inst_dmem_U17507 ( .A1(MEM_stage_inst_dmem_ram_2818), .A2(MEM_stage_inst_dmem_n18714), .ZN(MEM_stage_inst_dmem_n18711) );
NAND2_X1 MEM_stage_inst_dmem_U17506 ( .A1(MEM_stage_inst_dmem_n18709), .A2(MEM_stage_inst_dmem_n18708), .ZN(MEM_stage_inst_dmem_n10046) );
NAND2_X1 MEM_stage_inst_dmem_U17505 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n18715), .ZN(MEM_stage_inst_dmem_n18708) );
NAND2_X1 MEM_stage_inst_dmem_U17504 ( .A1(MEM_stage_inst_dmem_ram_2819), .A2(MEM_stage_inst_dmem_n18714), .ZN(MEM_stage_inst_dmem_n18709) );
NAND2_X1 MEM_stage_inst_dmem_U17503 ( .A1(MEM_stage_inst_dmem_n18707), .A2(MEM_stage_inst_dmem_n18706), .ZN(MEM_stage_inst_dmem_n10047) );
NAND2_X1 MEM_stage_inst_dmem_U17502 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n18715), .ZN(MEM_stage_inst_dmem_n18706) );
NAND2_X1 MEM_stage_inst_dmem_U17501 ( .A1(MEM_stage_inst_dmem_ram_2820), .A2(MEM_stage_inst_dmem_n18714), .ZN(MEM_stage_inst_dmem_n18707) );
NAND2_X1 MEM_stage_inst_dmem_U17500 ( .A1(MEM_stage_inst_dmem_n18705), .A2(MEM_stage_inst_dmem_n18704), .ZN(MEM_stage_inst_dmem_n10048) );
NAND2_X1 MEM_stage_inst_dmem_U17499 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n18715), .ZN(MEM_stage_inst_dmem_n18704) );
NAND2_X1 MEM_stage_inst_dmem_U17498 ( .A1(MEM_stage_inst_dmem_ram_2821), .A2(MEM_stage_inst_dmem_n18714), .ZN(MEM_stage_inst_dmem_n18705) );
NAND2_X1 MEM_stage_inst_dmem_U17497 ( .A1(MEM_stage_inst_dmem_n18703), .A2(MEM_stage_inst_dmem_n18702), .ZN(MEM_stage_inst_dmem_n10049) );
NAND2_X1 MEM_stage_inst_dmem_U17496 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n18715), .ZN(MEM_stage_inst_dmem_n18702) );
NAND2_X1 MEM_stage_inst_dmem_U17495 ( .A1(MEM_stage_inst_dmem_ram_2822), .A2(MEM_stage_inst_dmem_n18714), .ZN(MEM_stage_inst_dmem_n18703) );
NAND2_X1 MEM_stage_inst_dmem_U17494 ( .A1(MEM_stage_inst_dmem_n18701), .A2(MEM_stage_inst_dmem_n18700), .ZN(MEM_stage_inst_dmem_n10050) );
NAND2_X1 MEM_stage_inst_dmem_U17493 ( .A1(EX_pipeline_reg_out_12), .A2(MEM_stage_inst_dmem_n18715), .ZN(MEM_stage_inst_dmem_n18700) );
NAND2_X1 MEM_stage_inst_dmem_U17492 ( .A1(MEM_stage_inst_dmem_ram_2823), .A2(MEM_stage_inst_dmem_n18714), .ZN(MEM_stage_inst_dmem_n18701) );
NAND2_X1 MEM_stage_inst_dmem_U17491 ( .A1(MEM_stage_inst_dmem_n18699), .A2(MEM_stage_inst_dmem_n18698), .ZN(MEM_stage_inst_dmem_n10051) );
NAND2_X1 MEM_stage_inst_dmem_U17490 ( .A1(MEM_stage_inst_dmem_n13051), .A2(MEM_stage_inst_dmem_n18715), .ZN(MEM_stage_inst_dmem_n18698) );
NAND2_X1 MEM_stage_inst_dmem_U17489 ( .A1(MEM_stage_inst_dmem_ram_2824), .A2(MEM_stage_inst_dmem_n18714), .ZN(MEM_stage_inst_dmem_n18699) );
NAND2_X1 MEM_stage_inst_dmem_U17488 ( .A1(MEM_stage_inst_dmem_n18697), .A2(MEM_stage_inst_dmem_n18696), .ZN(MEM_stage_inst_dmem_n10052) );
NAND2_X1 MEM_stage_inst_dmem_U17487 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n18715), .ZN(MEM_stage_inst_dmem_n18696) );
NAND2_X1 MEM_stage_inst_dmem_U17486 ( .A1(MEM_stage_inst_dmem_ram_2825), .A2(MEM_stage_inst_dmem_n18714), .ZN(MEM_stage_inst_dmem_n18697) );
NAND2_X1 MEM_stage_inst_dmem_U17485 ( .A1(MEM_stage_inst_dmem_n18695), .A2(MEM_stage_inst_dmem_n18694), .ZN(MEM_stage_inst_dmem_n10053) );
NAND2_X1 MEM_stage_inst_dmem_U17484 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n18715), .ZN(MEM_stage_inst_dmem_n18694) );
NAND2_X1 MEM_stage_inst_dmem_U17483 ( .A1(MEM_stage_inst_dmem_ram_2826), .A2(MEM_stage_inst_dmem_n18714), .ZN(MEM_stage_inst_dmem_n18695) );
NAND2_X1 MEM_stage_inst_dmem_U17482 ( .A1(MEM_stage_inst_dmem_n18693), .A2(MEM_stage_inst_dmem_n18692), .ZN(MEM_stage_inst_dmem_n10054) );
NAND2_X1 MEM_stage_inst_dmem_U17481 ( .A1(MEM_stage_inst_dmem_n20904), .A2(MEM_stage_inst_dmem_n18715), .ZN(MEM_stage_inst_dmem_n18692) );
NAND2_X1 MEM_stage_inst_dmem_U17480 ( .A1(MEM_stage_inst_dmem_ram_2827), .A2(MEM_stage_inst_dmem_n18714), .ZN(MEM_stage_inst_dmem_n18693) );
NAND2_X1 MEM_stage_inst_dmem_U17479 ( .A1(MEM_stage_inst_dmem_n18691), .A2(MEM_stage_inst_dmem_n18690), .ZN(MEM_stage_inst_dmem_n10055) );
NAND2_X1 MEM_stage_inst_dmem_U17478 ( .A1(MEM_stage_inst_dmem_n21474), .A2(MEM_stage_inst_dmem_n18715), .ZN(MEM_stage_inst_dmem_n18690) );
NAND2_X1 MEM_stage_inst_dmem_U17477 ( .A1(MEM_stage_inst_dmem_ram_2828), .A2(MEM_stage_inst_dmem_n18714), .ZN(MEM_stage_inst_dmem_n18691) );
NAND2_X1 MEM_stage_inst_dmem_U17476 ( .A1(MEM_stage_inst_dmem_n18689), .A2(MEM_stage_inst_dmem_n18688), .ZN(MEM_stage_inst_dmem_n10056) );
NAND2_X1 MEM_stage_inst_dmem_U17475 ( .A1(MEM_stage_inst_dmem_n19242), .A2(MEM_stage_inst_dmem_n18715), .ZN(MEM_stage_inst_dmem_n18688) );
NAND2_X1 MEM_stage_inst_dmem_U17474 ( .A1(MEM_stage_inst_dmem_ram_2829), .A2(MEM_stage_inst_dmem_n18714), .ZN(MEM_stage_inst_dmem_n18689) );
NAND2_X1 MEM_stage_inst_dmem_U17473 ( .A1(MEM_stage_inst_dmem_n18687), .A2(MEM_stage_inst_dmem_n18686), .ZN(MEM_stage_inst_dmem_n10057) );
NAND2_X1 MEM_stage_inst_dmem_U17472 ( .A1(MEM_stage_inst_dmem_n115), .A2(MEM_stage_inst_dmem_n18715), .ZN(MEM_stage_inst_dmem_n18686) );
NAND2_X1 MEM_stage_inst_dmem_U17471 ( .A1(MEM_stage_inst_dmem_ram_2830), .A2(MEM_stage_inst_dmem_n18714), .ZN(MEM_stage_inst_dmem_n18687) );
NAND2_X1 MEM_stage_inst_dmem_U17470 ( .A1(MEM_stage_inst_dmem_n18685), .A2(MEM_stage_inst_dmem_n18684), .ZN(MEM_stage_inst_dmem_n10058) );
NAND2_X1 MEM_stage_inst_dmem_U17469 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n18715), .ZN(MEM_stage_inst_dmem_n18684) );
INV_X1 MEM_stage_inst_dmem_U17468 ( .A(MEM_stage_inst_dmem_n18714), .ZN(MEM_stage_inst_dmem_n18715) );
NAND2_X1 MEM_stage_inst_dmem_U17467 ( .A1(MEM_stage_inst_dmem_ram_2831), .A2(MEM_stage_inst_dmem_n18714), .ZN(MEM_stage_inst_dmem_n18685) );
NAND2_X1 MEM_stage_inst_dmem_U17466 ( .A1(MEM_stage_inst_dmem_n21465), .A2(MEM_stage_inst_dmem_n18683), .ZN(MEM_stage_inst_dmem_n18714) );
NAND2_X1 MEM_stage_inst_dmem_U17465 ( .A1(MEM_stage_inst_dmem_n18682), .A2(MEM_stage_inst_dmem_n18681), .ZN(MEM_stage_inst_dmem_n10059) );
NAND2_X1 MEM_stage_inst_dmem_U17464 ( .A1(MEM_stage_inst_dmem_n19275), .A2(MEM_stage_inst_dmem_n18680), .ZN(MEM_stage_inst_dmem_n18681) );
NAND2_X1 MEM_stage_inst_dmem_U17463 ( .A1(MEM_stage_inst_dmem_ram_2832), .A2(MEM_stage_inst_dmem_n18679), .ZN(MEM_stage_inst_dmem_n18682) );
NAND2_X1 MEM_stage_inst_dmem_U17462 ( .A1(MEM_stage_inst_dmem_n18678), .A2(MEM_stage_inst_dmem_n18677), .ZN(MEM_stage_inst_dmem_n10060) );
NAND2_X1 MEM_stage_inst_dmem_U17461 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n18680), .ZN(MEM_stage_inst_dmem_n18677) );
NAND2_X1 MEM_stage_inst_dmem_U17460 ( .A1(MEM_stage_inst_dmem_ram_2833), .A2(MEM_stage_inst_dmem_n18679), .ZN(MEM_stage_inst_dmem_n18678) );
NAND2_X1 MEM_stage_inst_dmem_U17459 ( .A1(MEM_stage_inst_dmem_n18676), .A2(MEM_stage_inst_dmem_n18675), .ZN(MEM_stage_inst_dmem_n10061) );
NAND2_X1 MEM_stage_inst_dmem_U17458 ( .A1(MEM_stage_inst_dmem_n20544), .A2(MEM_stage_inst_dmem_n18680), .ZN(MEM_stage_inst_dmem_n18675) );
NAND2_X1 MEM_stage_inst_dmem_U17457 ( .A1(MEM_stage_inst_dmem_ram_2834), .A2(MEM_stage_inst_dmem_n18679), .ZN(MEM_stage_inst_dmem_n18676) );
NAND2_X1 MEM_stage_inst_dmem_U17456 ( .A1(MEM_stage_inst_dmem_n18674), .A2(MEM_stage_inst_dmem_n18673), .ZN(MEM_stage_inst_dmem_n10062) );
NAND2_X1 MEM_stage_inst_dmem_U17455 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n18680), .ZN(MEM_stage_inst_dmem_n18673) );
NAND2_X1 MEM_stage_inst_dmem_U17454 ( .A1(MEM_stage_inst_dmem_ram_2835), .A2(MEM_stage_inst_dmem_n18679), .ZN(MEM_stage_inst_dmem_n18674) );
NAND2_X1 MEM_stage_inst_dmem_U17453 ( .A1(MEM_stage_inst_dmem_n18672), .A2(MEM_stage_inst_dmem_n18671), .ZN(MEM_stage_inst_dmem_n10063) );
NAND2_X1 MEM_stage_inst_dmem_U17452 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n18680), .ZN(MEM_stage_inst_dmem_n18671) );
NAND2_X1 MEM_stage_inst_dmem_U17451 ( .A1(MEM_stage_inst_dmem_ram_2836), .A2(MEM_stage_inst_dmem_n18679), .ZN(MEM_stage_inst_dmem_n18672) );
NAND2_X1 MEM_stage_inst_dmem_U17450 ( .A1(MEM_stage_inst_dmem_n18670), .A2(MEM_stage_inst_dmem_n18669), .ZN(MEM_stage_inst_dmem_n10064) );
NAND2_X1 MEM_stage_inst_dmem_U17449 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n18680), .ZN(MEM_stage_inst_dmem_n18669) );
NAND2_X1 MEM_stage_inst_dmem_U17448 ( .A1(MEM_stage_inst_dmem_ram_2837), .A2(MEM_stage_inst_dmem_n18679), .ZN(MEM_stage_inst_dmem_n18670) );
NAND2_X1 MEM_stage_inst_dmem_U17447 ( .A1(MEM_stage_inst_dmem_n18668), .A2(MEM_stage_inst_dmem_n18667), .ZN(MEM_stage_inst_dmem_n10065) );
NAND2_X1 MEM_stage_inst_dmem_U17446 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n18680), .ZN(MEM_stage_inst_dmem_n18667) );
NAND2_X1 MEM_stage_inst_dmem_U17445 ( .A1(MEM_stage_inst_dmem_ram_2838), .A2(MEM_stage_inst_dmem_n18679), .ZN(MEM_stage_inst_dmem_n18668) );
NAND2_X1 MEM_stage_inst_dmem_U17444 ( .A1(MEM_stage_inst_dmem_n18666), .A2(MEM_stage_inst_dmem_n18665), .ZN(MEM_stage_inst_dmem_n10066) );
NAND2_X1 MEM_stage_inst_dmem_U17443 ( .A1(MEM_stage_inst_dmem_n112), .A2(MEM_stage_inst_dmem_n18680), .ZN(MEM_stage_inst_dmem_n18665) );
NAND2_X1 MEM_stage_inst_dmem_U17442 ( .A1(MEM_stage_inst_dmem_ram_2839), .A2(MEM_stage_inst_dmem_n18679), .ZN(MEM_stage_inst_dmem_n18666) );
NAND2_X1 MEM_stage_inst_dmem_U17441 ( .A1(MEM_stage_inst_dmem_n18664), .A2(MEM_stage_inst_dmem_n18663), .ZN(MEM_stage_inst_dmem_n10067) );
NAND2_X1 MEM_stage_inst_dmem_U17440 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n18680), .ZN(MEM_stage_inst_dmem_n18663) );
NAND2_X1 MEM_stage_inst_dmem_U17439 ( .A1(MEM_stage_inst_dmem_ram_2840), .A2(MEM_stage_inst_dmem_n18679), .ZN(MEM_stage_inst_dmem_n18664) );
NAND2_X1 MEM_stage_inst_dmem_U17438 ( .A1(MEM_stage_inst_dmem_n18662), .A2(MEM_stage_inst_dmem_n18661), .ZN(MEM_stage_inst_dmem_n10068) );
NAND2_X1 MEM_stage_inst_dmem_U17437 ( .A1(MEM_stage_inst_dmem_n19251), .A2(MEM_stage_inst_dmem_n18680), .ZN(MEM_stage_inst_dmem_n18661) );
NAND2_X1 MEM_stage_inst_dmem_U17436 ( .A1(MEM_stage_inst_dmem_ram_2841), .A2(MEM_stage_inst_dmem_n18679), .ZN(MEM_stage_inst_dmem_n18662) );
NAND2_X1 MEM_stage_inst_dmem_U17435 ( .A1(MEM_stage_inst_dmem_n18660), .A2(MEM_stage_inst_dmem_n18659), .ZN(MEM_stage_inst_dmem_n10069) );
NAND2_X1 MEM_stage_inst_dmem_U17434 ( .A1(MEM_stage_inst_dmem_n20521), .A2(MEM_stage_inst_dmem_n18680), .ZN(MEM_stage_inst_dmem_n18659) );
NAND2_X1 MEM_stage_inst_dmem_U17433 ( .A1(MEM_stage_inst_dmem_ram_2842), .A2(MEM_stage_inst_dmem_n18679), .ZN(MEM_stage_inst_dmem_n18660) );
NAND2_X1 MEM_stage_inst_dmem_U17432 ( .A1(MEM_stage_inst_dmem_n18658), .A2(MEM_stage_inst_dmem_n18657), .ZN(MEM_stage_inst_dmem_n10070) );
NAND2_X1 MEM_stage_inst_dmem_U17431 ( .A1(MEM_stage_inst_dmem_n14705), .A2(MEM_stage_inst_dmem_n18680), .ZN(MEM_stage_inst_dmem_n18657) );
NAND2_X1 MEM_stage_inst_dmem_U17430 ( .A1(MEM_stage_inst_dmem_ram_2843), .A2(MEM_stage_inst_dmem_n18679), .ZN(MEM_stage_inst_dmem_n18658) );
NAND2_X1 MEM_stage_inst_dmem_U17429 ( .A1(MEM_stage_inst_dmem_n18656), .A2(MEM_stage_inst_dmem_n18655), .ZN(MEM_stage_inst_dmem_n10071) );
NAND2_X1 MEM_stage_inst_dmem_U17428 ( .A1(MEM_stage_inst_dmem_n14702), .A2(MEM_stage_inst_dmem_n18680), .ZN(MEM_stage_inst_dmem_n18655) );
NAND2_X1 MEM_stage_inst_dmem_U17427 ( .A1(MEM_stage_inst_dmem_ram_2844), .A2(MEM_stage_inst_dmem_n18679), .ZN(MEM_stage_inst_dmem_n18656) );
NAND2_X1 MEM_stage_inst_dmem_U17426 ( .A1(MEM_stage_inst_dmem_n18654), .A2(MEM_stage_inst_dmem_n18653), .ZN(MEM_stage_inst_dmem_n10072) );
NAND2_X1 MEM_stage_inst_dmem_U17425 ( .A1(MEM_stage_inst_dmem_n19242), .A2(MEM_stage_inst_dmem_n18680), .ZN(MEM_stage_inst_dmem_n18653) );
NAND2_X1 MEM_stage_inst_dmem_U17424 ( .A1(MEM_stage_inst_dmem_ram_2845), .A2(MEM_stage_inst_dmem_n18679), .ZN(MEM_stage_inst_dmem_n18654) );
NAND2_X1 MEM_stage_inst_dmem_U17423 ( .A1(MEM_stage_inst_dmem_n18652), .A2(MEM_stage_inst_dmem_n18651), .ZN(MEM_stage_inst_dmem_n10073) );
NAND2_X1 MEM_stage_inst_dmem_U17422 ( .A1(MEM_stage_inst_dmem_n115), .A2(MEM_stage_inst_dmem_n18680), .ZN(MEM_stage_inst_dmem_n18651) );
NAND2_X1 MEM_stage_inst_dmem_U17421 ( .A1(MEM_stage_inst_dmem_ram_2846), .A2(MEM_stage_inst_dmem_n18679), .ZN(MEM_stage_inst_dmem_n18652) );
NAND2_X1 MEM_stage_inst_dmem_U17420 ( .A1(MEM_stage_inst_dmem_n18650), .A2(MEM_stage_inst_dmem_n18649), .ZN(MEM_stage_inst_dmem_n10074) );
NAND2_X1 MEM_stage_inst_dmem_U17419 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n18680), .ZN(MEM_stage_inst_dmem_n18649) );
INV_X1 MEM_stage_inst_dmem_U17418 ( .A(MEM_stage_inst_dmem_n18679), .ZN(MEM_stage_inst_dmem_n18680) );
NAND2_X1 MEM_stage_inst_dmem_U17417 ( .A1(MEM_stage_inst_dmem_ram_2847), .A2(MEM_stage_inst_dmem_n18679), .ZN(MEM_stage_inst_dmem_n18650) );
NAND2_X1 MEM_stage_inst_dmem_U17416 ( .A1(MEM_stage_inst_dmem_n21429), .A2(MEM_stage_inst_dmem_n18683), .ZN(MEM_stage_inst_dmem_n18679) );
NAND2_X1 MEM_stage_inst_dmem_U17415 ( .A1(MEM_stage_inst_dmem_n18648), .A2(MEM_stage_inst_dmem_n18647), .ZN(MEM_stage_inst_dmem_n10075) );
NAND2_X1 MEM_stage_inst_dmem_U17414 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n18646), .ZN(MEM_stage_inst_dmem_n18647) );
NAND2_X1 MEM_stage_inst_dmem_U17413 ( .A1(MEM_stage_inst_dmem_ram_2848), .A2(MEM_stage_inst_dmem_n18645), .ZN(MEM_stage_inst_dmem_n18648) );
NAND2_X1 MEM_stage_inst_dmem_U17412 ( .A1(MEM_stage_inst_dmem_n18644), .A2(MEM_stage_inst_dmem_n18643), .ZN(MEM_stage_inst_dmem_n10076) );
NAND2_X1 MEM_stage_inst_dmem_U17411 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n18646), .ZN(MEM_stage_inst_dmem_n18643) );
NAND2_X1 MEM_stage_inst_dmem_U17410 ( .A1(MEM_stage_inst_dmem_ram_2849), .A2(MEM_stage_inst_dmem_n18645), .ZN(MEM_stage_inst_dmem_n18644) );
NAND2_X1 MEM_stage_inst_dmem_U17409 ( .A1(MEM_stage_inst_dmem_n18642), .A2(MEM_stage_inst_dmem_n18641), .ZN(MEM_stage_inst_dmem_n10077) );
NAND2_X1 MEM_stage_inst_dmem_U17408 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n18646), .ZN(MEM_stage_inst_dmem_n18641) );
NAND2_X1 MEM_stage_inst_dmem_U17407 ( .A1(MEM_stage_inst_dmem_ram_2850), .A2(MEM_stage_inst_dmem_n18645), .ZN(MEM_stage_inst_dmem_n18642) );
NAND2_X1 MEM_stage_inst_dmem_U17406 ( .A1(MEM_stage_inst_dmem_n18640), .A2(MEM_stage_inst_dmem_n18639), .ZN(MEM_stage_inst_dmem_n10078) );
NAND2_X1 MEM_stage_inst_dmem_U17405 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n18646), .ZN(MEM_stage_inst_dmem_n18639) );
NAND2_X1 MEM_stage_inst_dmem_U17404 ( .A1(MEM_stage_inst_dmem_ram_2851), .A2(MEM_stage_inst_dmem_n18645), .ZN(MEM_stage_inst_dmem_n18640) );
NAND2_X1 MEM_stage_inst_dmem_U17403 ( .A1(MEM_stage_inst_dmem_n18638), .A2(MEM_stage_inst_dmem_n18637), .ZN(MEM_stage_inst_dmem_n10079) );
NAND2_X1 MEM_stage_inst_dmem_U17402 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n18646), .ZN(MEM_stage_inst_dmem_n18637) );
NAND2_X1 MEM_stage_inst_dmem_U17401 ( .A1(MEM_stage_inst_dmem_ram_2852), .A2(MEM_stage_inst_dmem_n18645), .ZN(MEM_stage_inst_dmem_n18638) );
NAND2_X1 MEM_stage_inst_dmem_U17400 ( .A1(MEM_stage_inst_dmem_n18636), .A2(MEM_stage_inst_dmem_n18635), .ZN(MEM_stage_inst_dmem_n10080) );
NAND2_X1 MEM_stage_inst_dmem_U17399 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n18646), .ZN(MEM_stage_inst_dmem_n18635) );
NAND2_X1 MEM_stage_inst_dmem_U17398 ( .A1(MEM_stage_inst_dmem_ram_2853), .A2(MEM_stage_inst_dmem_n18645), .ZN(MEM_stage_inst_dmem_n18636) );
NAND2_X1 MEM_stage_inst_dmem_U17397 ( .A1(MEM_stage_inst_dmem_n18634), .A2(MEM_stage_inst_dmem_n18633), .ZN(MEM_stage_inst_dmem_n10081) );
NAND2_X1 MEM_stage_inst_dmem_U17396 ( .A1(MEM_stage_inst_dmem_n21340), .A2(MEM_stage_inst_dmem_n18646), .ZN(MEM_stage_inst_dmem_n18633) );
NAND2_X1 MEM_stage_inst_dmem_U17395 ( .A1(MEM_stage_inst_dmem_ram_2854), .A2(MEM_stage_inst_dmem_n18645), .ZN(MEM_stage_inst_dmem_n18634) );
NAND2_X1 MEM_stage_inst_dmem_U17394 ( .A1(MEM_stage_inst_dmem_n18632), .A2(MEM_stage_inst_dmem_n18631), .ZN(MEM_stage_inst_dmem_n10082) );
NAND2_X1 MEM_stage_inst_dmem_U17393 ( .A1(MEM_stage_inst_dmem_n17), .A2(MEM_stage_inst_dmem_n18646), .ZN(MEM_stage_inst_dmem_n18631) );
NAND2_X1 MEM_stage_inst_dmem_U17392 ( .A1(MEM_stage_inst_dmem_ram_2855), .A2(MEM_stage_inst_dmem_n18645), .ZN(MEM_stage_inst_dmem_n18632) );
NAND2_X1 MEM_stage_inst_dmem_U17391 ( .A1(MEM_stage_inst_dmem_n18630), .A2(MEM_stage_inst_dmem_n18629), .ZN(MEM_stage_inst_dmem_n10083) );
NAND2_X1 MEM_stage_inst_dmem_U17390 ( .A1(MEM_stage_inst_dmem_n21335), .A2(MEM_stage_inst_dmem_n18646), .ZN(MEM_stage_inst_dmem_n18629) );
NAND2_X1 MEM_stage_inst_dmem_U17389 ( .A1(MEM_stage_inst_dmem_ram_2856), .A2(MEM_stage_inst_dmem_n18645), .ZN(MEM_stage_inst_dmem_n18630) );
NAND2_X1 MEM_stage_inst_dmem_U17388 ( .A1(MEM_stage_inst_dmem_n18628), .A2(MEM_stage_inst_dmem_n18627), .ZN(MEM_stage_inst_dmem_n10084) );
NAND2_X1 MEM_stage_inst_dmem_U17387 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n18646), .ZN(MEM_stage_inst_dmem_n18627) );
NAND2_X1 MEM_stage_inst_dmem_U17386 ( .A1(MEM_stage_inst_dmem_ram_2857), .A2(MEM_stage_inst_dmem_n18645), .ZN(MEM_stage_inst_dmem_n18628) );
NAND2_X1 MEM_stage_inst_dmem_U17385 ( .A1(MEM_stage_inst_dmem_n18626), .A2(MEM_stage_inst_dmem_n18625), .ZN(MEM_stage_inst_dmem_n10085) );
NAND2_X1 MEM_stage_inst_dmem_U17384 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n18646), .ZN(MEM_stage_inst_dmem_n18625) );
NAND2_X1 MEM_stage_inst_dmem_U17383 ( .A1(MEM_stage_inst_dmem_ram_2858), .A2(MEM_stage_inst_dmem_n18645), .ZN(MEM_stage_inst_dmem_n18626) );
NAND2_X1 MEM_stage_inst_dmem_U17382 ( .A1(MEM_stage_inst_dmem_n18624), .A2(MEM_stage_inst_dmem_n18623), .ZN(MEM_stage_inst_dmem_n10086) );
NAND2_X1 MEM_stage_inst_dmem_U17381 ( .A1(MEM_stage_inst_dmem_n13044), .A2(MEM_stage_inst_dmem_n18646), .ZN(MEM_stage_inst_dmem_n18623) );
NAND2_X1 MEM_stage_inst_dmem_U17380 ( .A1(MEM_stage_inst_dmem_ram_2859), .A2(MEM_stage_inst_dmem_n18645), .ZN(MEM_stage_inst_dmem_n18624) );
NAND2_X1 MEM_stage_inst_dmem_U17379 ( .A1(MEM_stage_inst_dmem_n18622), .A2(MEM_stage_inst_dmem_n18621), .ZN(MEM_stage_inst_dmem_n10087) );
NAND2_X1 MEM_stage_inst_dmem_U17378 ( .A1(MEM_stage_inst_dmem_n13041), .A2(MEM_stage_inst_dmem_n18646), .ZN(MEM_stage_inst_dmem_n18621) );
NAND2_X1 MEM_stage_inst_dmem_U17377 ( .A1(MEM_stage_inst_dmem_ram_2860), .A2(MEM_stage_inst_dmem_n18645), .ZN(MEM_stage_inst_dmem_n18622) );
NAND2_X1 MEM_stage_inst_dmem_U17376 ( .A1(MEM_stage_inst_dmem_n18620), .A2(MEM_stage_inst_dmem_n18619), .ZN(MEM_stage_inst_dmem_n10088) );
NAND2_X1 MEM_stage_inst_dmem_U17375 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n18646), .ZN(MEM_stage_inst_dmem_n18619) );
NAND2_X1 MEM_stage_inst_dmem_U17374 ( .A1(MEM_stage_inst_dmem_ram_2861), .A2(MEM_stage_inst_dmem_n18645), .ZN(MEM_stage_inst_dmem_n18620) );
NAND2_X1 MEM_stage_inst_dmem_U17373 ( .A1(MEM_stage_inst_dmem_n18618), .A2(MEM_stage_inst_dmem_n18617), .ZN(MEM_stage_inst_dmem_n10089) );
NAND2_X1 MEM_stage_inst_dmem_U17372 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n18646), .ZN(MEM_stage_inst_dmem_n18617) );
NAND2_X1 MEM_stage_inst_dmem_U17371 ( .A1(MEM_stage_inst_dmem_ram_2862), .A2(MEM_stage_inst_dmem_n18645), .ZN(MEM_stage_inst_dmem_n18618) );
NAND2_X1 MEM_stage_inst_dmem_U17370 ( .A1(MEM_stage_inst_dmem_n18616), .A2(MEM_stage_inst_dmem_n18615), .ZN(MEM_stage_inst_dmem_n10090) );
NAND2_X1 MEM_stage_inst_dmem_U17369 ( .A1(MEM_stage_inst_dmem_n21320), .A2(MEM_stage_inst_dmem_n18646), .ZN(MEM_stage_inst_dmem_n18615) );
INV_X1 MEM_stage_inst_dmem_U17368 ( .A(MEM_stage_inst_dmem_n18645), .ZN(MEM_stage_inst_dmem_n18646) );
NAND2_X1 MEM_stage_inst_dmem_U17367 ( .A1(MEM_stage_inst_dmem_ram_2863), .A2(MEM_stage_inst_dmem_n18645), .ZN(MEM_stage_inst_dmem_n18616) );
NAND2_X1 MEM_stage_inst_dmem_U17366 ( .A1(MEM_stage_inst_dmem_n21394), .A2(MEM_stage_inst_dmem_n18683), .ZN(MEM_stage_inst_dmem_n18645) );
NAND2_X1 MEM_stage_inst_dmem_U17365 ( .A1(MEM_stage_inst_dmem_n18614), .A2(MEM_stage_inst_dmem_n18613), .ZN(MEM_stage_inst_dmem_n10091) );
NAND2_X1 MEM_stage_inst_dmem_U17364 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n18612), .ZN(MEM_stage_inst_dmem_n18613) );
NAND2_X1 MEM_stage_inst_dmem_U17363 ( .A1(MEM_stage_inst_dmem_ram_2864), .A2(MEM_stage_inst_dmem_n18611), .ZN(MEM_stage_inst_dmem_n18614) );
NAND2_X1 MEM_stage_inst_dmem_U17362 ( .A1(MEM_stage_inst_dmem_n18610), .A2(MEM_stage_inst_dmem_n18609), .ZN(MEM_stage_inst_dmem_n10092) );
NAND2_X1 MEM_stage_inst_dmem_U17361 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n18612), .ZN(MEM_stage_inst_dmem_n18609) );
NAND2_X1 MEM_stage_inst_dmem_U17360 ( .A1(MEM_stage_inst_dmem_ram_2865), .A2(MEM_stage_inst_dmem_n18611), .ZN(MEM_stage_inst_dmem_n18610) );
NAND2_X1 MEM_stage_inst_dmem_U17359 ( .A1(MEM_stage_inst_dmem_n18608), .A2(MEM_stage_inst_dmem_n18607), .ZN(MEM_stage_inst_dmem_n10093) );
NAND2_X1 MEM_stage_inst_dmem_U17358 ( .A1(MEM_stage_inst_dmem_n18887), .A2(MEM_stage_inst_dmem_n18612), .ZN(MEM_stage_inst_dmem_n18607) );
NAND2_X1 MEM_stage_inst_dmem_U17357 ( .A1(MEM_stage_inst_dmem_ram_2866), .A2(MEM_stage_inst_dmem_n18611), .ZN(MEM_stage_inst_dmem_n18608) );
NAND2_X1 MEM_stage_inst_dmem_U17356 ( .A1(MEM_stage_inst_dmem_n18606), .A2(MEM_stage_inst_dmem_n18605), .ZN(MEM_stage_inst_dmem_n10094) );
NAND2_X1 MEM_stage_inst_dmem_U17355 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n18612), .ZN(MEM_stage_inst_dmem_n18605) );
NAND2_X1 MEM_stage_inst_dmem_U17354 ( .A1(MEM_stage_inst_dmem_ram_2867), .A2(MEM_stage_inst_dmem_n18611), .ZN(MEM_stage_inst_dmem_n18606) );
NAND2_X1 MEM_stage_inst_dmem_U17353 ( .A1(MEM_stage_inst_dmem_n18604), .A2(MEM_stage_inst_dmem_n18603), .ZN(MEM_stage_inst_dmem_n10095) );
NAND2_X1 MEM_stage_inst_dmem_U17352 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n18612), .ZN(MEM_stage_inst_dmem_n18603) );
NAND2_X1 MEM_stage_inst_dmem_U17351 ( .A1(MEM_stage_inst_dmem_ram_2868), .A2(MEM_stage_inst_dmem_n18611), .ZN(MEM_stage_inst_dmem_n18604) );
NAND2_X1 MEM_stage_inst_dmem_U17350 ( .A1(MEM_stage_inst_dmem_n18602), .A2(MEM_stage_inst_dmem_n18601), .ZN(MEM_stage_inst_dmem_n10096) );
NAND2_X1 MEM_stage_inst_dmem_U17349 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n18612), .ZN(MEM_stage_inst_dmem_n18601) );
NAND2_X1 MEM_stage_inst_dmem_U17348 ( .A1(MEM_stage_inst_dmem_ram_2869), .A2(MEM_stage_inst_dmem_n18611), .ZN(MEM_stage_inst_dmem_n18602) );
NAND2_X1 MEM_stage_inst_dmem_U17347 ( .A1(MEM_stage_inst_dmem_n18600), .A2(MEM_stage_inst_dmem_n18599), .ZN(MEM_stage_inst_dmem_n10097) );
NAND2_X1 MEM_stage_inst_dmem_U17346 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n18612), .ZN(MEM_stage_inst_dmem_n18599) );
NAND2_X1 MEM_stage_inst_dmem_U17345 ( .A1(MEM_stage_inst_dmem_ram_2870), .A2(MEM_stage_inst_dmem_n18611), .ZN(MEM_stage_inst_dmem_n18600) );
NAND2_X1 MEM_stage_inst_dmem_U17344 ( .A1(MEM_stage_inst_dmem_n18598), .A2(MEM_stage_inst_dmem_n18597), .ZN(MEM_stage_inst_dmem_n10098) );
NAND2_X1 MEM_stage_inst_dmem_U17343 ( .A1(MEM_stage_inst_dmem_n18875), .A2(MEM_stage_inst_dmem_n18612), .ZN(MEM_stage_inst_dmem_n18597) );
NAND2_X1 MEM_stage_inst_dmem_U17342 ( .A1(MEM_stage_inst_dmem_ram_2871), .A2(MEM_stage_inst_dmem_n18611), .ZN(MEM_stage_inst_dmem_n18598) );
NAND2_X1 MEM_stage_inst_dmem_U17341 ( .A1(MEM_stage_inst_dmem_n18596), .A2(MEM_stage_inst_dmem_n18595), .ZN(MEM_stage_inst_dmem_n10099) );
NAND2_X1 MEM_stage_inst_dmem_U17340 ( .A1(MEM_stage_inst_dmem_n111), .A2(MEM_stage_inst_dmem_n18612), .ZN(MEM_stage_inst_dmem_n18595) );
NAND2_X1 MEM_stage_inst_dmem_U17339 ( .A1(MEM_stage_inst_dmem_ram_2872), .A2(MEM_stage_inst_dmem_n18611), .ZN(MEM_stage_inst_dmem_n18596) );
NAND2_X1 MEM_stage_inst_dmem_U17338 ( .A1(MEM_stage_inst_dmem_n18594), .A2(MEM_stage_inst_dmem_n18593), .ZN(MEM_stage_inst_dmem_n10100) );
NAND2_X1 MEM_stage_inst_dmem_U17337 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n18612), .ZN(MEM_stage_inst_dmem_n18593) );
NAND2_X1 MEM_stage_inst_dmem_U17336 ( .A1(MEM_stage_inst_dmem_ram_2873), .A2(MEM_stage_inst_dmem_n18611), .ZN(MEM_stage_inst_dmem_n18594) );
NAND2_X1 MEM_stage_inst_dmem_U17335 ( .A1(MEM_stage_inst_dmem_n18592), .A2(MEM_stage_inst_dmem_n18591), .ZN(MEM_stage_inst_dmem_n10101) );
NAND2_X1 MEM_stage_inst_dmem_U17334 ( .A1(MEM_stage_inst_dmem_n18867), .A2(MEM_stage_inst_dmem_n18612), .ZN(MEM_stage_inst_dmem_n18591) );
NAND2_X1 MEM_stage_inst_dmem_U17333 ( .A1(MEM_stage_inst_dmem_ram_2874), .A2(MEM_stage_inst_dmem_n18611), .ZN(MEM_stage_inst_dmem_n18592) );
NAND2_X1 MEM_stage_inst_dmem_U17332 ( .A1(MEM_stage_inst_dmem_n18590), .A2(MEM_stage_inst_dmem_n18589), .ZN(MEM_stage_inst_dmem_n10102) );
NAND2_X1 MEM_stage_inst_dmem_U17331 ( .A1(MEM_stage_inst_dmem_n18864), .A2(MEM_stage_inst_dmem_n18612), .ZN(MEM_stage_inst_dmem_n18589) );
NAND2_X1 MEM_stage_inst_dmem_U17330 ( .A1(MEM_stage_inst_dmem_ram_2875), .A2(MEM_stage_inst_dmem_n18611), .ZN(MEM_stage_inst_dmem_n18590) );
NAND2_X1 MEM_stage_inst_dmem_U17329 ( .A1(MEM_stage_inst_dmem_n18588), .A2(MEM_stage_inst_dmem_n18587), .ZN(MEM_stage_inst_dmem_n10103) );
NAND2_X1 MEM_stage_inst_dmem_U17328 ( .A1(MEM_stage_inst_dmem_n18861), .A2(MEM_stage_inst_dmem_n18612), .ZN(MEM_stage_inst_dmem_n18587) );
NAND2_X1 MEM_stage_inst_dmem_U17327 ( .A1(MEM_stage_inst_dmem_ram_2876), .A2(MEM_stage_inst_dmem_n18611), .ZN(MEM_stage_inst_dmem_n18588) );
NAND2_X1 MEM_stage_inst_dmem_U17326 ( .A1(MEM_stage_inst_dmem_n18586), .A2(MEM_stage_inst_dmem_n18585), .ZN(MEM_stage_inst_dmem_n10104) );
NAND2_X1 MEM_stage_inst_dmem_U17325 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n18612), .ZN(MEM_stage_inst_dmem_n18585) );
NAND2_X1 MEM_stage_inst_dmem_U17324 ( .A1(MEM_stage_inst_dmem_ram_2877), .A2(MEM_stage_inst_dmem_n18611), .ZN(MEM_stage_inst_dmem_n18586) );
NAND2_X1 MEM_stage_inst_dmem_U17323 ( .A1(MEM_stage_inst_dmem_n18584), .A2(MEM_stage_inst_dmem_n18583), .ZN(MEM_stage_inst_dmem_n10105) );
NAND2_X1 MEM_stage_inst_dmem_U17322 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n18612), .ZN(MEM_stage_inst_dmem_n18583) );
NAND2_X1 MEM_stage_inst_dmem_U17321 ( .A1(MEM_stage_inst_dmem_ram_2878), .A2(MEM_stage_inst_dmem_n18611), .ZN(MEM_stage_inst_dmem_n18584) );
NAND2_X1 MEM_stage_inst_dmem_U17320 ( .A1(MEM_stage_inst_dmem_n18582), .A2(MEM_stage_inst_dmem_n18581), .ZN(MEM_stage_inst_dmem_n10106) );
NAND2_X1 MEM_stage_inst_dmem_U17319 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n18612), .ZN(MEM_stage_inst_dmem_n18581) );
NAND2_X1 MEM_stage_inst_dmem_U17318 ( .A1(MEM_stage_inst_dmem_ram_2879), .A2(MEM_stage_inst_dmem_n18611), .ZN(MEM_stage_inst_dmem_n18582) );
NAND2_X1 MEM_stage_inst_dmem_U17317 ( .A1(MEM_stage_inst_dmem_n21359), .A2(MEM_stage_inst_dmem_n18683), .ZN(MEM_stage_inst_dmem_n18611) );
NAND2_X1 MEM_stage_inst_dmem_U17316 ( .A1(MEM_stage_inst_dmem_n18580), .A2(MEM_stage_inst_dmem_n18579), .ZN(MEM_stage_inst_dmem_n10107) );
NAND2_X1 MEM_stage_inst_dmem_U17315 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n18578), .ZN(MEM_stage_inst_dmem_n18579) );
NAND2_X1 MEM_stage_inst_dmem_U17314 ( .A1(MEM_stage_inst_dmem_ram_2880), .A2(MEM_stage_inst_dmem_n18577), .ZN(MEM_stage_inst_dmem_n18580) );
NAND2_X1 MEM_stage_inst_dmem_U17313 ( .A1(MEM_stage_inst_dmem_n18576), .A2(MEM_stage_inst_dmem_n18575), .ZN(MEM_stage_inst_dmem_n10108) );
NAND2_X1 MEM_stage_inst_dmem_U17312 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n18578), .ZN(MEM_stage_inst_dmem_n18575) );
NAND2_X1 MEM_stage_inst_dmem_U17311 ( .A1(MEM_stage_inst_dmem_ram_2881), .A2(MEM_stage_inst_dmem_n18577), .ZN(MEM_stage_inst_dmem_n18576) );
NAND2_X1 MEM_stage_inst_dmem_U17310 ( .A1(MEM_stage_inst_dmem_n18574), .A2(MEM_stage_inst_dmem_n18573), .ZN(MEM_stage_inst_dmem_n10109) );
NAND2_X1 MEM_stage_inst_dmem_U17309 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n18578), .ZN(MEM_stage_inst_dmem_n18573) );
NAND2_X1 MEM_stage_inst_dmem_U17308 ( .A1(MEM_stage_inst_dmem_ram_2882), .A2(MEM_stage_inst_dmem_n18577), .ZN(MEM_stage_inst_dmem_n18574) );
NAND2_X1 MEM_stage_inst_dmem_U17307 ( .A1(MEM_stage_inst_dmem_n18572), .A2(MEM_stage_inst_dmem_n18571), .ZN(MEM_stage_inst_dmem_n10110) );
NAND2_X1 MEM_stage_inst_dmem_U17306 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n18578), .ZN(MEM_stage_inst_dmem_n18571) );
NAND2_X1 MEM_stage_inst_dmem_U17305 ( .A1(MEM_stage_inst_dmem_ram_2883), .A2(MEM_stage_inst_dmem_n18577), .ZN(MEM_stage_inst_dmem_n18572) );
NAND2_X1 MEM_stage_inst_dmem_U17304 ( .A1(MEM_stage_inst_dmem_n18570), .A2(MEM_stage_inst_dmem_n18569), .ZN(MEM_stage_inst_dmem_n10111) );
NAND2_X1 MEM_stage_inst_dmem_U17303 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n18578), .ZN(MEM_stage_inst_dmem_n18569) );
NAND2_X1 MEM_stage_inst_dmem_U17302 ( .A1(MEM_stage_inst_dmem_ram_2884), .A2(MEM_stage_inst_dmem_n18577), .ZN(MEM_stage_inst_dmem_n18570) );
NAND2_X1 MEM_stage_inst_dmem_U17301 ( .A1(MEM_stage_inst_dmem_n18568), .A2(MEM_stage_inst_dmem_n18567), .ZN(MEM_stage_inst_dmem_n10112) );
NAND2_X1 MEM_stage_inst_dmem_U17300 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n18578), .ZN(MEM_stage_inst_dmem_n18567) );
NAND2_X1 MEM_stage_inst_dmem_U17299 ( .A1(MEM_stage_inst_dmem_ram_2885), .A2(MEM_stage_inst_dmem_n18577), .ZN(MEM_stage_inst_dmem_n18568) );
NAND2_X1 MEM_stage_inst_dmem_U17298 ( .A1(MEM_stage_inst_dmem_n18566), .A2(MEM_stage_inst_dmem_n18565), .ZN(MEM_stage_inst_dmem_n10113) );
NAND2_X1 MEM_stage_inst_dmem_U17297 ( .A1(MEM_stage_inst_dmem_n21340), .A2(MEM_stage_inst_dmem_n18578), .ZN(MEM_stage_inst_dmem_n18565) );
NAND2_X1 MEM_stage_inst_dmem_U17296 ( .A1(MEM_stage_inst_dmem_ram_2886), .A2(MEM_stage_inst_dmem_n18577), .ZN(MEM_stage_inst_dmem_n18566) );
NAND2_X1 MEM_stage_inst_dmem_U17295 ( .A1(MEM_stage_inst_dmem_n18564), .A2(MEM_stage_inst_dmem_n18563), .ZN(MEM_stage_inst_dmem_n10114) );
NAND2_X1 MEM_stage_inst_dmem_U17294 ( .A1(MEM_stage_inst_dmem_n18), .A2(MEM_stage_inst_dmem_n18578), .ZN(MEM_stage_inst_dmem_n18563) );
NAND2_X1 MEM_stage_inst_dmem_U17293 ( .A1(MEM_stage_inst_dmem_ram_2887), .A2(MEM_stage_inst_dmem_n18577), .ZN(MEM_stage_inst_dmem_n18564) );
NAND2_X1 MEM_stage_inst_dmem_U17292 ( .A1(MEM_stage_inst_dmem_n18562), .A2(MEM_stage_inst_dmem_n18561), .ZN(MEM_stage_inst_dmem_n10115) );
NAND2_X1 MEM_stage_inst_dmem_U17291 ( .A1(MEM_stage_inst_dmem_n21335), .A2(MEM_stage_inst_dmem_n18578), .ZN(MEM_stage_inst_dmem_n18561) );
NAND2_X1 MEM_stage_inst_dmem_U17290 ( .A1(MEM_stage_inst_dmem_ram_2888), .A2(MEM_stage_inst_dmem_n18577), .ZN(MEM_stage_inst_dmem_n18562) );
NAND2_X1 MEM_stage_inst_dmem_U17289 ( .A1(MEM_stage_inst_dmem_n18560), .A2(MEM_stage_inst_dmem_n18559), .ZN(MEM_stage_inst_dmem_n10116) );
NAND2_X1 MEM_stage_inst_dmem_U17288 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n18578), .ZN(MEM_stage_inst_dmem_n18559) );
NAND2_X1 MEM_stage_inst_dmem_U17287 ( .A1(MEM_stage_inst_dmem_ram_2889), .A2(MEM_stage_inst_dmem_n18577), .ZN(MEM_stage_inst_dmem_n18560) );
NAND2_X1 MEM_stage_inst_dmem_U17286 ( .A1(MEM_stage_inst_dmem_n18558), .A2(MEM_stage_inst_dmem_n18557), .ZN(MEM_stage_inst_dmem_n10117) );
NAND2_X1 MEM_stage_inst_dmem_U17285 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n18578), .ZN(MEM_stage_inst_dmem_n18557) );
NAND2_X1 MEM_stage_inst_dmem_U17284 ( .A1(MEM_stage_inst_dmem_ram_2890), .A2(MEM_stage_inst_dmem_n18577), .ZN(MEM_stage_inst_dmem_n18558) );
NAND2_X1 MEM_stage_inst_dmem_U17283 ( .A1(MEM_stage_inst_dmem_n18556), .A2(MEM_stage_inst_dmem_n18555), .ZN(MEM_stage_inst_dmem_n10118) );
NAND2_X1 MEM_stage_inst_dmem_U17282 ( .A1(MEM_stage_inst_dmem_n20904), .A2(MEM_stage_inst_dmem_n18578), .ZN(MEM_stage_inst_dmem_n18555) );
NAND2_X1 MEM_stage_inst_dmem_U17281 ( .A1(MEM_stage_inst_dmem_ram_2891), .A2(MEM_stage_inst_dmem_n18577), .ZN(MEM_stage_inst_dmem_n18556) );
NAND2_X1 MEM_stage_inst_dmem_U17280 ( .A1(MEM_stage_inst_dmem_n18554), .A2(MEM_stage_inst_dmem_n18553), .ZN(MEM_stage_inst_dmem_n10119) );
NAND2_X1 MEM_stage_inst_dmem_U17279 ( .A1(MEM_stage_inst_dmem_n21474), .A2(MEM_stage_inst_dmem_n18578), .ZN(MEM_stage_inst_dmem_n18553) );
NAND2_X1 MEM_stage_inst_dmem_U17278 ( .A1(MEM_stage_inst_dmem_ram_2892), .A2(MEM_stage_inst_dmem_n18577), .ZN(MEM_stage_inst_dmem_n18554) );
NAND2_X1 MEM_stage_inst_dmem_U17277 ( .A1(MEM_stage_inst_dmem_n18552), .A2(MEM_stage_inst_dmem_n18551), .ZN(MEM_stage_inst_dmem_n10120) );
NAND2_X1 MEM_stage_inst_dmem_U17276 ( .A1(EX_pipeline_reg_out_18), .A2(MEM_stage_inst_dmem_n18578), .ZN(MEM_stage_inst_dmem_n18551) );
NAND2_X1 MEM_stage_inst_dmem_U17275 ( .A1(MEM_stage_inst_dmem_ram_2893), .A2(MEM_stage_inst_dmem_n18577), .ZN(MEM_stage_inst_dmem_n18552) );
NAND2_X1 MEM_stage_inst_dmem_U17274 ( .A1(MEM_stage_inst_dmem_n18550), .A2(MEM_stage_inst_dmem_n18549), .ZN(MEM_stage_inst_dmem_n10121) );
NAND2_X1 MEM_stage_inst_dmem_U17273 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n18578), .ZN(MEM_stage_inst_dmem_n18549) );
NAND2_X1 MEM_stage_inst_dmem_U17272 ( .A1(MEM_stage_inst_dmem_ram_2894), .A2(MEM_stage_inst_dmem_n18577), .ZN(MEM_stage_inst_dmem_n18550) );
NAND2_X1 MEM_stage_inst_dmem_U17271 ( .A1(MEM_stage_inst_dmem_n18548), .A2(MEM_stage_inst_dmem_n18547), .ZN(MEM_stage_inst_dmem_n10122) );
NAND2_X1 MEM_stage_inst_dmem_U17270 ( .A1(MEM_stage_inst_dmem_n21320), .A2(MEM_stage_inst_dmem_n18578), .ZN(MEM_stage_inst_dmem_n18547) );
INV_X1 MEM_stage_inst_dmem_U17269 ( .A(MEM_stage_inst_dmem_n18577), .ZN(MEM_stage_inst_dmem_n18578) );
NAND2_X1 MEM_stage_inst_dmem_U17268 ( .A1(MEM_stage_inst_dmem_ram_2895), .A2(MEM_stage_inst_dmem_n18577), .ZN(MEM_stage_inst_dmem_n18548) );
NAND2_X1 MEM_stage_inst_dmem_U17267 ( .A1(MEM_stage_inst_dmem_n21319), .A2(MEM_stage_inst_dmem_n18683), .ZN(MEM_stage_inst_dmem_n18577) );
NAND2_X1 MEM_stage_inst_dmem_U17266 ( .A1(MEM_stage_inst_dmem_n18546), .A2(MEM_stage_inst_dmem_n18545), .ZN(MEM_stage_inst_dmem_n10123) );
NAND2_X1 MEM_stage_inst_dmem_U17265 ( .A1(MEM_stage_inst_dmem_n19275), .A2(MEM_stage_inst_dmem_n18544), .ZN(MEM_stage_inst_dmem_n18545) );
NAND2_X1 MEM_stage_inst_dmem_U17264 ( .A1(MEM_stage_inst_dmem_ram_2896), .A2(MEM_stage_inst_dmem_n18543), .ZN(MEM_stage_inst_dmem_n18546) );
NAND2_X1 MEM_stage_inst_dmem_U17263 ( .A1(MEM_stage_inst_dmem_n18542), .A2(MEM_stage_inst_dmem_n18541), .ZN(MEM_stage_inst_dmem_n10124) );
NAND2_X1 MEM_stage_inst_dmem_U17262 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n18544), .ZN(MEM_stage_inst_dmem_n18541) );
NAND2_X1 MEM_stage_inst_dmem_U17261 ( .A1(MEM_stage_inst_dmem_ram_2897), .A2(MEM_stage_inst_dmem_n18543), .ZN(MEM_stage_inst_dmem_n18542) );
NAND2_X1 MEM_stage_inst_dmem_U17260 ( .A1(MEM_stage_inst_dmem_n18540), .A2(MEM_stage_inst_dmem_n18539), .ZN(MEM_stage_inst_dmem_n10125) );
NAND2_X1 MEM_stage_inst_dmem_U17259 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n18544), .ZN(MEM_stage_inst_dmem_n18539) );
NAND2_X1 MEM_stage_inst_dmem_U17258 ( .A1(MEM_stage_inst_dmem_ram_2898), .A2(MEM_stage_inst_dmem_n18543), .ZN(MEM_stage_inst_dmem_n18540) );
NAND2_X1 MEM_stage_inst_dmem_U17257 ( .A1(MEM_stage_inst_dmem_n18538), .A2(MEM_stage_inst_dmem_n18537), .ZN(MEM_stage_inst_dmem_n10126) );
NAND2_X1 MEM_stage_inst_dmem_U17256 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n18544), .ZN(MEM_stage_inst_dmem_n18537) );
NAND2_X1 MEM_stage_inst_dmem_U17255 ( .A1(MEM_stage_inst_dmem_ram_2899), .A2(MEM_stage_inst_dmem_n18543), .ZN(MEM_stage_inst_dmem_n18538) );
NAND2_X1 MEM_stage_inst_dmem_U17254 ( .A1(MEM_stage_inst_dmem_n18536), .A2(MEM_stage_inst_dmem_n18535), .ZN(MEM_stage_inst_dmem_n10127) );
NAND2_X1 MEM_stage_inst_dmem_U17253 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n18544), .ZN(MEM_stage_inst_dmem_n18535) );
NAND2_X1 MEM_stage_inst_dmem_U17252 ( .A1(MEM_stage_inst_dmem_ram_2900), .A2(MEM_stage_inst_dmem_n18543), .ZN(MEM_stage_inst_dmem_n18536) );
NAND2_X1 MEM_stage_inst_dmem_U17251 ( .A1(MEM_stage_inst_dmem_n18534), .A2(MEM_stage_inst_dmem_n18533), .ZN(MEM_stage_inst_dmem_n10128) );
NAND2_X1 MEM_stage_inst_dmem_U17250 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n18544), .ZN(MEM_stage_inst_dmem_n18533) );
NAND2_X1 MEM_stage_inst_dmem_U17249 ( .A1(MEM_stage_inst_dmem_ram_2901), .A2(MEM_stage_inst_dmem_n18543), .ZN(MEM_stage_inst_dmem_n18534) );
NAND2_X1 MEM_stage_inst_dmem_U17248 ( .A1(MEM_stage_inst_dmem_n18532), .A2(MEM_stage_inst_dmem_n18531), .ZN(MEM_stage_inst_dmem_n10129) );
NAND2_X1 MEM_stage_inst_dmem_U17247 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n18544), .ZN(MEM_stage_inst_dmem_n18531) );
NAND2_X1 MEM_stage_inst_dmem_U17246 ( .A1(MEM_stage_inst_dmem_ram_2902), .A2(MEM_stage_inst_dmem_n18543), .ZN(MEM_stage_inst_dmem_n18532) );
NAND2_X1 MEM_stage_inst_dmem_U17245 ( .A1(MEM_stage_inst_dmem_n18530), .A2(MEM_stage_inst_dmem_n18529), .ZN(MEM_stage_inst_dmem_n10130) );
NAND2_X1 MEM_stage_inst_dmem_U17244 ( .A1(MEM_stage_inst_dmem_n13886), .A2(MEM_stage_inst_dmem_n18544), .ZN(MEM_stage_inst_dmem_n18529) );
NAND2_X1 MEM_stage_inst_dmem_U17243 ( .A1(MEM_stage_inst_dmem_ram_2903), .A2(MEM_stage_inst_dmem_n18543), .ZN(MEM_stage_inst_dmem_n18530) );
NAND2_X1 MEM_stage_inst_dmem_U17242 ( .A1(MEM_stage_inst_dmem_n18528), .A2(MEM_stage_inst_dmem_n18527), .ZN(MEM_stage_inst_dmem_n10131) );
NAND2_X1 MEM_stage_inst_dmem_U17241 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n18544), .ZN(MEM_stage_inst_dmem_n18527) );
NAND2_X1 MEM_stage_inst_dmem_U17240 ( .A1(MEM_stage_inst_dmem_ram_2904), .A2(MEM_stage_inst_dmem_n18543), .ZN(MEM_stage_inst_dmem_n18528) );
NAND2_X1 MEM_stage_inst_dmem_U17239 ( .A1(MEM_stage_inst_dmem_n18526), .A2(MEM_stage_inst_dmem_n18525), .ZN(MEM_stage_inst_dmem_n10132) );
NAND2_X1 MEM_stage_inst_dmem_U17238 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n18544), .ZN(MEM_stage_inst_dmem_n18525) );
NAND2_X1 MEM_stage_inst_dmem_U17237 ( .A1(MEM_stage_inst_dmem_ram_2905), .A2(MEM_stage_inst_dmem_n18543), .ZN(MEM_stage_inst_dmem_n18526) );
NAND2_X1 MEM_stage_inst_dmem_U17236 ( .A1(MEM_stage_inst_dmem_n18524), .A2(MEM_stage_inst_dmem_n18523), .ZN(MEM_stage_inst_dmem_n10133) );
NAND2_X1 MEM_stage_inst_dmem_U17235 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n18544), .ZN(MEM_stage_inst_dmem_n18523) );
NAND2_X1 MEM_stage_inst_dmem_U17234 ( .A1(MEM_stage_inst_dmem_ram_2906), .A2(MEM_stage_inst_dmem_n18543), .ZN(MEM_stage_inst_dmem_n18524) );
NAND2_X1 MEM_stage_inst_dmem_U17233 ( .A1(MEM_stage_inst_dmem_n18522), .A2(MEM_stage_inst_dmem_n18521), .ZN(MEM_stage_inst_dmem_n10134) );
NAND2_X1 MEM_stage_inst_dmem_U17232 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n18544), .ZN(MEM_stage_inst_dmem_n18521) );
NAND2_X1 MEM_stage_inst_dmem_U17231 ( .A1(MEM_stage_inst_dmem_ram_2907), .A2(MEM_stage_inst_dmem_n18543), .ZN(MEM_stage_inst_dmem_n18522) );
NAND2_X1 MEM_stage_inst_dmem_U17230 ( .A1(MEM_stage_inst_dmem_n18520), .A2(MEM_stage_inst_dmem_n18519), .ZN(MEM_stage_inst_dmem_n10135) );
NAND2_X1 MEM_stage_inst_dmem_U17229 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n18544), .ZN(MEM_stage_inst_dmem_n18519) );
NAND2_X1 MEM_stage_inst_dmem_U17228 ( .A1(MEM_stage_inst_dmem_ram_2908), .A2(MEM_stage_inst_dmem_n18543), .ZN(MEM_stage_inst_dmem_n18520) );
NAND2_X1 MEM_stage_inst_dmem_U17227 ( .A1(MEM_stage_inst_dmem_n18518), .A2(MEM_stage_inst_dmem_n18517), .ZN(MEM_stage_inst_dmem_n10136) );
NAND2_X1 MEM_stage_inst_dmem_U17226 ( .A1(MEM_stage_inst_dmem_n19242), .A2(MEM_stage_inst_dmem_n18544), .ZN(MEM_stage_inst_dmem_n18517) );
NAND2_X1 MEM_stage_inst_dmem_U17225 ( .A1(MEM_stage_inst_dmem_ram_2909), .A2(MEM_stage_inst_dmem_n18543), .ZN(MEM_stage_inst_dmem_n18518) );
NAND2_X1 MEM_stage_inst_dmem_U17224 ( .A1(MEM_stage_inst_dmem_n18516), .A2(MEM_stage_inst_dmem_n18515), .ZN(MEM_stage_inst_dmem_n10137) );
NAND2_X1 MEM_stage_inst_dmem_U17223 ( .A1(MEM_stage_inst_dmem_n115), .A2(MEM_stage_inst_dmem_n18544), .ZN(MEM_stage_inst_dmem_n18515) );
NAND2_X1 MEM_stage_inst_dmem_U17222 ( .A1(MEM_stage_inst_dmem_ram_2910), .A2(MEM_stage_inst_dmem_n18543), .ZN(MEM_stage_inst_dmem_n18516) );
NAND2_X1 MEM_stage_inst_dmem_U17221 ( .A1(MEM_stage_inst_dmem_n18514), .A2(MEM_stage_inst_dmem_n18513), .ZN(MEM_stage_inst_dmem_n10138) );
NAND2_X1 MEM_stage_inst_dmem_U17220 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n18544), .ZN(MEM_stage_inst_dmem_n18513) );
INV_X1 MEM_stage_inst_dmem_U17219 ( .A(MEM_stage_inst_dmem_n18543), .ZN(MEM_stage_inst_dmem_n18544) );
NAND2_X1 MEM_stage_inst_dmem_U17218 ( .A1(MEM_stage_inst_dmem_ram_2911), .A2(MEM_stage_inst_dmem_n18543), .ZN(MEM_stage_inst_dmem_n18514) );
NAND2_X1 MEM_stage_inst_dmem_U17217 ( .A1(MEM_stage_inst_dmem_n21284), .A2(MEM_stage_inst_dmem_n18683), .ZN(MEM_stage_inst_dmem_n18543) );
NAND2_X1 MEM_stage_inst_dmem_U17216 ( .A1(MEM_stage_inst_dmem_n18512), .A2(MEM_stage_inst_dmem_n18511), .ZN(MEM_stage_inst_dmem_n10139) );
NAND2_X1 MEM_stage_inst_dmem_U17215 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n18510), .ZN(MEM_stage_inst_dmem_n18511) );
NAND2_X1 MEM_stage_inst_dmem_U17214 ( .A1(MEM_stage_inst_dmem_ram_2912), .A2(MEM_stage_inst_dmem_n18509), .ZN(MEM_stage_inst_dmem_n18512) );
NAND2_X1 MEM_stage_inst_dmem_U17213 ( .A1(MEM_stage_inst_dmem_n18508), .A2(MEM_stage_inst_dmem_n18507), .ZN(MEM_stage_inst_dmem_n10140) );
NAND2_X1 MEM_stage_inst_dmem_U17212 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n18510), .ZN(MEM_stage_inst_dmem_n18507) );
NAND2_X1 MEM_stage_inst_dmem_U17211 ( .A1(MEM_stage_inst_dmem_ram_2913), .A2(MEM_stage_inst_dmem_n18509), .ZN(MEM_stage_inst_dmem_n18508) );
NAND2_X1 MEM_stage_inst_dmem_U17210 ( .A1(MEM_stage_inst_dmem_n18506), .A2(MEM_stage_inst_dmem_n18505), .ZN(MEM_stage_inst_dmem_n10141) );
NAND2_X1 MEM_stage_inst_dmem_U17209 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n18510), .ZN(MEM_stage_inst_dmem_n18505) );
NAND2_X1 MEM_stage_inst_dmem_U17208 ( .A1(MEM_stage_inst_dmem_ram_2914), .A2(MEM_stage_inst_dmem_n18509), .ZN(MEM_stage_inst_dmem_n18506) );
NAND2_X1 MEM_stage_inst_dmem_U17207 ( .A1(MEM_stage_inst_dmem_n18504), .A2(MEM_stage_inst_dmem_n18503), .ZN(MEM_stage_inst_dmem_n10142) );
NAND2_X1 MEM_stage_inst_dmem_U17206 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n18510), .ZN(MEM_stage_inst_dmem_n18503) );
NAND2_X1 MEM_stage_inst_dmem_U17205 ( .A1(MEM_stage_inst_dmem_ram_2915), .A2(MEM_stage_inst_dmem_n18509), .ZN(MEM_stage_inst_dmem_n18504) );
NAND2_X1 MEM_stage_inst_dmem_U17204 ( .A1(MEM_stage_inst_dmem_n18502), .A2(MEM_stage_inst_dmem_n18501), .ZN(MEM_stage_inst_dmem_n10143) );
NAND2_X1 MEM_stage_inst_dmem_U17203 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n18510), .ZN(MEM_stage_inst_dmem_n18501) );
NAND2_X1 MEM_stage_inst_dmem_U17202 ( .A1(MEM_stage_inst_dmem_ram_2916), .A2(MEM_stage_inst_dmem_n18509), .ZN(MEM_stage_inst_dmem_n18502) );
NAND2_X1 MEM_stage_inst_dmem_U17201 ( .A1(MEM_stage_inst_dmem_n18500), .A2(MEM_stage_inst_dmem_n18499), .ZN(MEM_stage_inst_dmem_n10144) );
NAND2_X1 MEM_stage_inst_dmem_U17200 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n18510), .ZN(MEM_stage_inst_dmem_n18499) );
NAND2_X1 MEM_stage_inst_dmem_U17199 ( .A1(MEM_stage_inst_dmem_ram_2917), .A2(MEM_stage_inst_dmem_n18509), .ZN(MEM_stage_inst_dmem_n18500) );
NAND2_X1 MEM_stage_inst_dmem_U17198 ( .A1(MEM_stage_inst_dmem_n18498), .A2(MEM_stage_inst_dmem_n18497), .ZN(MEM_stage_inst_dmem_n10145) );
NAND2_X1 MEM_stage_inst_dmem_U17197 ( .A1(MEM_stage_inst_dmem_n21340), .A2(MEM_stage_inst_dmem_n18510), .ZN(MEM_stage_inst_dmem_n18497) );
NAND2_X1 MEM_stage_inst_dmem_U17196 ( .A1(MEM_stage_inst_dmem_ram_2918), .A2(MEM_stage_inst_dmem_n18509), .ZN(MEM_stage_inst_dmem_n18498) );
NAND2_X1 MEM_stage_inst_dmem_U17195 ( .A1(MEM_stage_inst_dmem_n18496), .A2(MEM_stage_inst_dmem_n18495), .ZN(MEM_stage_inst_dmem_n10146) );
NAND2_X1 MEM_stage_inst_dmem_U17194 ( .A1(MEM_stage_inst_dmem_n17), .A2(MEM_stage_inst_dmem_n18510), .ZN(MEM_stage_inst_dmem_n18495) );
NAND2_X1 MEM_stage_inst_dmem_U17193 ( .A1(MEM_stage_inst_dmem_ram_2919), .A2(MEM_stage_inst_dmem_n18509), .ZN(MEM_stage_inst_dmem_n18496) );
NAND2_X1 MEM_stage_inst_dmem_U17192 ( .A1(MEM_stage_inst_dmem_n18494), .A2(MEM_stage_inst_dmem_n18493), .ZN(MEM_stage_inst_dmem_n10147) );
NAND2_X1 MEM_stage_inst_dmem_U17191 ( .A1(MEM_stage_inst_dmem_n21335), .A2(MEM_stage_inst_dmem_n18510), .ZN(MEM_stage_inst_dmem_n18493) );
NAND2_X1 MEM_stage_inst_dmem_U17190 ( .A1(MEM_stage_inst_dmem_ram_2920), .A2(MEM_stage_inst_dmem_n18509), .ZN(MEM_stage_inst_dmem_n18494) );
NAND2_X1 MEM_stage_inst_dmem_U17189 ( .A1(MEM_stage_inst_dmem_n18492), .A2(MEM_stage_inst_dmem_n18491), .ZN(MEM_stage_inst_dmem_n10148) );
NAND2_X1 MEM_stage_inst_dmem_U17188 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n18510), .ZN(MEM_stage_inst_dmem_n18491) );
NAND2_X1 MEM_stage_inst_dmem_U17187 ( .A1(MEM_stage_inst_dmem_ram_2921), .A2(MEM_stage_inst_dmem_n18509), .ZN(MEM_stage_inst_dmem_n18492) );
NAND2_X1 MEM_stage_inst_dmem_U17186 ( .A1(MEM_stage_inst_dmem_n18490), .A2(MEM_stage_inst_dmem_n18489), .ZN(MEM_stage_inst_dmem_n10149) );
NAND2_X1 MEM_stage_inst_dmem_U17185 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n18510), .ZN(MEM_stage_inst_dmem_n18489) );
NAND2_X1 MEM_stage_inst_dmem_U17184 ( .A1(MEM_stage_inst_dmem_ram_2922), .A2(MEM_stage_inst_dmem_n18509), .ZN(MEM_stage_inst_dmem_n18490) );
NAND2_X1 MEM_stage_inst_dmem_U17183 ( .A1(MEM_stage_inst_dmem_n18488), .A2(MEM_stage_inst_dmem_n18487), .ZN(MEM_stage_inst_dmem_n10150) );
NAND2_X1 MEM_stage_inst_dmem_U17182 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n18510), .ZN(MEM_stage_inst_dmem_n18487) );
NAND2_X1 MEM_stage_inst_dmem_U17181 ( .A1(MEM_stage_inst_dmem_ram_2923), .A2(MEM_stage_inst_dmem_n18509), .ZN(MEM_stage_inst_dmem_n18488) );
NAND2_X1 MEM_stage_inst_dmem_U17180 ( .A1(MEM_stage_inst_dmem_n18486), .A2(MEM_stage_inst_dmem_n18485), .ZN(MEM_stage_inst_dmem_n10151) );
NAND2_X1 MEM_stage_inst_dmem_U17179 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n18510), .ZN(MEM_stage_inst_dmem_n18485) );
NAND2_X1 MEM_stage_inst_dmem_U17178 ( .A1(MEM_stage_inst_dmem_ram_2924), .A2(MEM_stage_inst_dmem_n18509), .ZN(MEM_stage_inst_dmem_n18486) );
NAND2_X1 MEM_stage_inst_dmem_U17177 ( .A1(MEM_stage_inst_dmem_n18484), .A2(MEM_stage_inst_dmem_n18483), .ZN(MEM_stage_inst_dmem_n10152) );
NAND2_X1 MEM_stage_inst_dmem_U17176 ( .A1(MEM_stage_inst_dmem_n20512), .A2(MEM_stage_inst_dmem_n18510), .ZN(MEM_stage_inst_dmem_n18483) );
NAND2_X1 MEM_stage_inst_dmem_U17175 ( .A1(MEM_stage_inst_dmem_ram_2925), .A2(MEM_stage_inst_dmem_n18509), .ZN(MEM_stage_inst_dmem_n18484) );
NAND2_X1 MEM_stage_inst_dmem_U17174 ( .A1(MEM_stage_inst_dmem_n18482), .A2(MEM_stage_inst_dmem_n18481), .ZN(MEM_stage_inst_dmem_n10153) );
NAND2_X1 MEM_stage_inst_dmem_U17173 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n18510), .ZN(MEM_stage_inst_dmem_n18481) );
NAND2_X1 MEM_stage_inst_dmem_U17172 ( .A1(MEM_stage_inst_dmem_ram_2926), .A2(MEM_stage_inst_dmem_n18509), .ZN(MEM_stage_inst_dmem_n18482) );
NAND2_X1 MEM_stage_inst_dmem_U17171 ( .A1(MEM_stage_inst_dmem_n18480), .A2(MEM_stage_inst_dmem_n18479), .ZN(MEM_stage_inst_dmem_n10154) );
NAND2_X1 MEM_stage_inst_dmem_U17170 ( .A1(MEM_stage_inst_dmem_n21320), .A2(MEM_stage_inst_dmem_n18510), .ZN(MEM_stage_inst_dmem_n18479) );
INV_X1 MEM_stage_inst_dmem_U17169 ( .A(MEM_stage_inst_dmem_n18509), .ZN(MEM_stage_inst_dmem_n18510) );
NAND2_X1 MEM_stage_inst_dmem_U17168 ( .A1(MEM_stage_inst_dmem_ram_2927), .A2(MEM_stage_inst_dmem_n18509), .ZN(MEM_stage_inst_dmem_n18480) );
NAND2_X1 MEM_stage_inst_dmem_U17167 ( .A1(MEM_stage_inst_dmem_n21249), .A2(MEM_stage_inst_dmem_n18683), .ZN(MEM_stage_inst_dmem_n18509) );
NAND2_X1 MEM_stage_inst_dmem_U17166 ( .A1(MEM_stage_inst_dmem_n18478), .A2(MEM_stage_inst_dmem_n18477), .ZN(MEM_stage_inst_dmem_n10155) );
NAND2_X1 MEM_stage_inst_dmem_U17165 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n18476), .ZN(MEM_stage_inst_dmem_n18477) );
NAND2_X1 MEM_stage_inst_dmem_U17164 ( .A1(MEM_stage_inst_dmem_ram_2928), .A2(MEM_stage_inst_dmem_n18475), .ZN(MEM_stage_inst_dmem_n18478) );
NAND2_X1 MEM_stage_inst_dmem_U17163 ( .A1(MEM_stage_inst_dmem_n18474), .A2(MEM_stage_inst_dmem_n18473), .ZN(MEM_stage_inst_dmem_n10156) );
NAND2_X1 MEM_stage_inst_dmem_U17162 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n18476), .ZN(MEM_stage_inst_dmem_n18473) );
NAND2_X1 MEM_stage_inst_dmem_U17161 ( .A1(MEM_stage_inst_dmem_ram_2929), .A2(MEM_stage_inst_dmem_n18475), .ZN(MEM_stage_inst_dmem_n18474) );
NAND2_X1 MEM_stage_inst_dmem_U17160 ( .A1(MEM_stage_inst_dmem_n18472), .A2(MEM_stage_inst_dmem_n18471), .ZN(MEM_stage_inst_dmem_n10157) );
NAND2_X1 MEM_stage_inst_dmem_U17159 ( .A1(MEM_stage_inst_dmem_n18887), .A2(MEM_stage_inst_dmem_n18476), .ZN(MEM_stage_inst_dmem_n18471) );
NAND2_X1 MEM_stage_inst_dmem_U17158 ( .A1(MEM_stage_inst_dmem_ram_2930), .A2(MEM_stage_inst_dmem_n18475), .ZN(MEM_stage_inst_dmem_n18472) );
NAND2_X1 MEM_stage_inst_dmem_U17157 ( .A1(MEM_stage_inst_dmem_n18470), .A2(MEM_stage_inst_dmem_n18469), .ZN(MEM_stage_inst_dmem_n10158) );
NAND2_X1 MEM_stage_inst_dmem_U17156 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n18476), .ZN(MEM_stage_inst_dmem_n18469) );
NAND2_X1 MEM_stage_inst_dmem_U17155 ( .A1(MEM_stage_inst_dmem_ram_2931), .A2(MEM_stage_inst_dmem_n18475), .ZN(MEM_stage_inst_dmem_n18470) );
NAND2_X1 MEM_stage_inst_dmem_U17154 ( .A1(MEM_stage_inst_dmem_n18468), .A2(MEM_stage_inst_dmem_n18467), .ZN(MEM_stage_inst_dmem_n10159) );
NAND2_X1 MEM_stage_inst_dmem_U17153 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n18476), .ZN(MEM_stage_inst_dmem_n18467) );
NAND2_X1 MEM_stage_inst_dmem_U17152 ( .A1(MEM_stage_inst_dmem_ram_2932), .A2(MEM_stage_inst_dmem_n18475), .ZN(MEM_stage_inst_dmem_n18468) );
NAND2_X1 MEM_stage_inst_dmem_U17151 ( .A1(MEM_stage_inst_dmem_n18466), .A2(MEM_stage_inst_dmem_n18465), .ZN(MEM_stage_inst_dmem_n10160) );
NAND2_X1 MEM_stage_inst_dmem_U17150 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n18476), .ZN(MEM_stage_inst_dmem_n18465) );
NAND2_X1 MEM_stage_inst_dmem_U17149 ( .A1(MEM_stage_inst_dmem_ram_2933), .A2(MEM_stage_inst_dmem_n18475), .ZN(MEM_stage_inst_dmem_n18466) );
NAND2_X1 MEM_stage_inst_dmem_U17148 ( .A1(MEM_stage_inst_dmem_n18464), .A2(MEM_stage_inst_dmem_n18463), .ZN(MEM_stage_inst_dmem_n10161) );
NAND2_X1 MEM_stage_inst_dmem_U17147 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n18476), .ZN(MEM_stage_inst_dmem_n18463) );
NAND2_X1 MEM_stage_inst_dmem_U17146 ( .A1(MEM_stage_inst_dmem_ram_2934), .A2(MEM_stage_inst_dmem_n18475), .ZN(MEM_stage_inst_dmem_n18464) );
NAND2_X1 MEM_stage_inst_dmem_U17145 ( .A1(MEM_stage_inst_dmem_n18462), .A2(MEM_stage_inst_dmem_n18461), .ZN(MEM_stage_inst_dmem_n10162) );
NAND2_X1 MEM_stage_inst_dmem_U17144 ( .A1(MEM_stage_inst_dmem_n18875), .A2(MEM_stage_inst_dmem_n18476), .ZN(MEM_stage_inst_dmem_n18461) );
NAND2_X1 MEM_stage_inst_dmem_U17143 ( .A1(MEM_stage_inst_dmem_ram_2935), .A2(MEM_stage_inst_dmem_n18475), .ZN(MEM_stage_inst_dmem_n18462) );
NAND2_X1 MEM_stage_inst_dmem_U17142 ( .A1(MEM_stage_inst_dmem_n18460), .A2(MEM_stage_inst_dmem_n18459), .ZN(MEM_stage_inst_dmem_n10163) );
NAND2_X1 MEM_stage_inst_dmem_U17141 ( .A1(MEM_stage_inst_dmem_n111), .A2(MEM_stage_inst_dmem_n18476), .ZN(MEM_stage_inst_dmem_n18459) );
NAND2_X1 MEM_stage_inst_dmem_U17140 ( .A1(MEM_stage_inst_dmem_ram_2936), .A2(MEM_stage_inst_dmem_n18475), .ZN(MEM_stage_inst_dmem_n18460) );
NAND2_X1 MEM_stage_inst_dmem_U17139 ( .A1(MEM_stage_inst_dmem_n18458), .A2(MEM_stage_inst_dmem_n18457), .ZN(MEM_stage_inst_dmem_n10164) );
NAND2_X1 MEM_stage_inst_dmem_U17138 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n18476), .ZN(MEM_stage_inst_dmem_n18457) );
NAND2_X1 MEM_stage_inst_dmem_U17137 ( .A1(MEM_stage_inst_dmem_ram_2937), .A2(MEM_stage_inst_dmem_n18475), .ZN(MEM_stage_inst_dmem_n18458) );
NAND2_X1 MEM_stage_inst_dmem_U17136 ( .A1(MEM_stage_inst_dmem_n18456), .A2(MEM_stage_inst_dmem_n18455), .ZN(MEM_stage_inst_dmem_n10165) );
NAND2_X1 MEM_stage_inst_dmem_U17135 ( .A1(MEM_stage_inst_dmem_n18867), .A2(MEM_stage_inst_dmem_n18476), .ZN(MEM_stage_inst_dmem_n18455) );
NAND2_X1 MEM_stage_inst_dmem_U17134 ( .A1(MEM_stage_inst_dmem_ram_2938), .A2(MEM_stage_inst_dmem_n18475), .ZN(MEM_stage_inst_dmem_n18456) );
NAND2_X1 MEM_stage_inst_dmem_U17133 ( .A1(MEM_stage_inst_dmem_n18454), .A2(MEM_stage_inst_dmem_n18453), .ZN(MEM_stage_inst_dmem_n10166) );
NAND2_X1 MEM_stage_inst_dmem_U17132 ( .A1(MEM_stage_inst_dmem_n18864), .A2(MEM_stage_inst_dmem_n18476), .ZN(MEM_stage_inst_dmem_n18453) );
NAND2_X1 MEM_stage_inst_dmem_U17131 ( .A1(MEM_stage_inst_dmem_ram_2939), .A2(MEM_stage_inst_dmem_n18475), .ZN(MEM_stage_inst_dmem_n18454) );
NAND2_X1 MEM_stage_inst_dmem_U17130 ( .A1(MEM_stage_inst_dmem_n18452), .A2(MEM_stage_inst_dmem_n18451), .ZN(MEM_stage_inst_dmem_n10167) );
NAND2_X1 MEM_stage_inst_dmem_U17129 ( .A1(MEM_stage_inst_dmem_n18861), .A2(MEM_stage_inst_dmem_n18476), .ZN(MEM_stage_inst_dmem_n18451) );
NAND2_X1 MEM_stage_inst_dmem_U17128 ( .A1(MEM_stage_inst_dmem_ram_2940), .A2(MEM_stage_inst_dmem_n18475), .ZN(MEM_stage_inst_dmem_n18452) );
NAND2_X1 MEM_stage_inst_dmem_U17127 ( .A1(MEM_stage_inst_dmem_n18450), .A2(MEM_stage_inst_dmem_n18449), .ZN(MEM_stage_inst_dmem_n10168) );
NAND2_X1 MEM_stage_inst_dmem_U17126 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n18476), .ZN(MEM_stage_inst_dmem_n18449) );
NAND2_X1 MEM_stage_inst_dmem_U17125 ( .A1(MEM_stage_inst_dmem_ram_2941), .A2(MEM_stage_inst_dmem_n18475), .ZN(MEM_stage_inst_dmem_n18450) );
NAND2_X1 MEM_stage_inst_dmem_U17124 ( .A1(MEM_stage_inst_dmem_n18448), .A2(MEM_stage_inst_dmem_n18447), .ZN(MEM_stage_inst_dmem_n10169) );
NAND2_X1 MEM_stage_inst_dmem_U17123 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n18476), .ZN(MEM_stage_inst_dmem_n18447) );
NAND2_X1 MEM_stage_inst_dmem_U17122 ( .A1(MEM_stage_inst_dmem_ram_2942), .A2(MEM_stage_inst_dmem_n18475), .ZN(MEM_stage_inst_dmem_n18448) );
NAND2_X1 MEM_stage_inst_dmem_U17121 ( .A1(MEM_stage_inst_dmem_n18446), .A2(MEM_stage_inst_dmem_n18445), .ZN(MEM_stage_inst_dmem_n10170) );
NAND2_X1 MEM_stage_inst_dmem_U17120 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n18476), .ZN(MEM_stage_inst_dmem_n18445) );
INV_X1 MEM_stage_inst_dmem_U17119 ( .A(MEM_stage_inst_dmem_n18475), .ZN(MEM_stage_inst_dmem_n18476) );
NAND2_X1 MEM_stage_inst_dmem_U17118 ( .A1(MEM_stage_inst_dmem_ram_2943), .A2(MEM_stage_inst_dmem_n18475), .ZN(MEM_stage_inst_dmem_n18446) );
NAND2_X1 MEM_stage_inst_dmem_U17117 ( .A1(MEM_stage_inst_dmem_n21214), .A2(MEM_stage_inst_dmem_n18683), .ZN(MEM_stage_inst_dmem_n18475) );
NAND2_X1 MEM_stage_inst_dmem_U17116 ( .A1(MEM_stage_inst_dmem_n18444), .A2(MEM_stage_inst_dmem_n18443), .ZN(MEM_stage_inst_dmem_n10171) );
NAND2_X1 MEM_stage_inst_dmem_U17115 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n18442), .ZN(MEM_stage_inst_dmem_n18443) );
NAND2_X1 MEM_stage_inst_dmem_U17114 ( .A1(MEM_stage_inst_dmem_ram_2944), .A2(MEM_stage_inst_dmem_n18441), .ZN(MEM_stage_inst_dmem_n18444) );
NAND2_X1 MEM_stage_inst_dmem_U17113 ( .A1(MEM_stage_inst_dmem_n18440), .A2(MEM_stage_inst_dmem_n18439), .ZN(MEM_stage_inst_dmem_n10172) );
NAND2_X1 MEM_stage_inst_dmem_U17112 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n18442), .ZN(MEM_stage_inst_dmem_n18439) );
NAND2_X1 MEM_stage_inst_dmem_U17111 ( .A1(MEM_stage_inst_dmem_ram_2945), .A2(MEM_stage_inst_dmem_n18441), .ZN(MEM_stage_inst_dmem_n18440) );
NAND2_X1 MEM_stage_inst_dmem_U17110 ( .A1(MEM_stage_inst_dmem_n18438), .A2(MEM_stage_inst_dmem_n18437), .ZN(MEM_stage_inst_dmem_n10173) );
NAND2_X1 MEM_stage_inst_dmem_U17109 ( .A1(MEM_stage_inst_dmem_n18887), .A2(MEM_stage_inst_dmem_n18442), .ZN(MEM_stage_inst_dmem_n18437) );
NAND2_X1 MEM_stage_inst_dmem_U17108 ( .A1(MEM_stage_inst_dmem_ram_2946), .A2(MEM_stage_inst_dmem_n18441), .ZN(MEM_stage_inst_dmem_n18438) );
NAND2_X1 MEM_stage_inst_dmem_U17107 ( .A1(MEM_stage_inst_dmem_n18436), .A2(MEM_stage_inst_dmem_n18435), .ZN(MEM_stage_inst_dmem_n10174) );
NAND2_X1 MEM_stage_inst_dmem_U17106 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n18442), .ZN(MEM_stage_inst_dmem_n18435) );
NAND2_X1 MEM_stage_inst_dmem_U17105 ( .A1(MEM_stage_inst_dmem_ram_2947), .A2(MEM_stage_inst_dmem_n18441), .ZN(MEM_stage_inst_dmem_n18436) );
NAND2_X1 MEM_stage_inst_dmem_U17104 ( .A1(MEM_stage_inst_dmem_n18434), .A2(MEM_stage_inst_dmem_n18433), .ZN(MEM_stage_inst_dmem_n10175) );
NAND2_X1 MEM_stage_inst_dmem_U17103 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n18442), .ZN(MEM_stage_inst_dmem_n18433) );
NAND2_X1 MEM_stage_inst_dmem_U17102 ( .A1(MEM_stage_inst_dmem_ram_2948), .A2(MEM_stage_inst_dmem_n18441), .ZN(MEM_stage_inst_dmem_n18434) );
NAND2_X1 MEM_stage_inst_dmem_U17101 ( .A1(MEM_stage_inst_dmem_n18432), .A2(MEM_stage_inst_dmem_n18431), .ZN(MEM_stage_inst_dmem_n10176) );
NAND2_X1 MEM_stage_inst_dmem_U17100 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n18442), .ZN(MEM_stage_inst_dmem_n18431) );
NAND2_X1 MEM_stage_inst_dmem_U17099 ( .A1(MEM_stage_inst_dmem_ram_2949), .A2(MEM_stage_inst_dmem_n18441), .ZN(MEM_stage_inst_dmem_n18432) );
NAND2_X1 MEM_stage_inst_dmem_U17098 ( .A1(MEM_stage_inst_dmem_n18430), .A2(MEM_stage_inst_dmem_n18429), .ZN(MEM_stage_inst_dmem_n10177) );
NAND2_X1 MEM_stage_inst_dmem_U17097 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n18442), .ZN(MEM_stage_inst_dmem_n18429) );
NAND2_X1 MEM_stage_inst_dmem_U17096 ( .A1(MEM_stage_inst_dmem_ram_2950), .A2(MEM_stage_inst_dmem_n18441), .ZN(MEM_stage_inst_dmem_n18430) );
NAND2_X1 MEM_stage_inst_dmem_U17095 ( .A1(MEM_stage_inst_dmem_n18428), .A2(MEM_stage_inst_dmem_n18427), .ZN(MEM_stage_inst_dmem_n10178) );
NAND2_X1 MEM_stage_inst_dmem_U17094 ( .A1(MEM_stage_inst_dmem_n18875), .A2(MEM_stage_inst_dmem_n18442), .ZN(MEM_stage_inst_dmem_n18427) );
NAND2_X1 MEM_stage_inst_dmem_U17093 ( .A1(MEM_stage_inst_dmem_ram_2951), .A2(MEM_stage_inst_dmem_n18441), .ZN(MEM_stage_inst_dmem_n18428) );
NAND2_X1 MEM_stage_inst_dmem_U17092 ( .A1(MEM_stage_inst_dmem_n18426), .A2(MEM_stage_inst_dmem_n18425), .ZN(MEM_stage_inst_dmem_n10179) );
NAND2_X1 MEM_stage_inst_dmem_U17091 ( .A1(MEM_stage_inst_dmem_n111), .A2(MEM_stage_inst_dmem_n18442), .ZN(MEM_stage_inst_dmem_n18425) );
NAND2_X1 MEM_stage_inst_dmem_U17090 ( .A1(MEM_stage_inst_dmem_ram_2952), .A2(MEM_stage_inst_dmem_n18441), .ZN(MEM_stage_inst_dmem_n18426) );
NAND2_X1 MEM_stage_inst_dmem_U17089 ( .A1(MEM_stage_inst_dmem_n18424), .A2(MEM_stage_inst_dmem_n18423), .ZN(MEM_stage_inst_dmem_n10180) );
NAND2_X1 MEM_stage_inst_dmem_U17088 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n18442), .ZN(MEM_stage_inst_dmem_n18423) );
NAND2_X1 MEM_stage_inst_dmem_U17087 ( .A1(MEM_stage_inst_dmem_ram_2953), .A2(MEM_stage_inst_dmem_n18441), .ZN(MEM_stage_inst_dmem_n18424) );
NAND2_X1 MEM_stage_inst_dmem_U17086 ( .A1(MEM_stage_inst_dmem_n18422), .A2(MEM_stage_inst_dmem_n18421), .ZN(MEM_stage_inst_dmem_n10181) );
NAND2_X1 MEM_stage_inst_dmem_U17085 ( .A1(MEM_stage_inst_dmem_n18867), .A2(MEM_stage_inst_dmem_n18442), .ZN(MEM_stage_inst_dmem_n18421) );
NAND2_X1 MEM_stage_inst_dmem_U17084 ( .A1(MEM_stage_inst_dmem_ram_2954), .A2(MEM_stage_inst_dmem_n18441), .ZN(MEM_stage_inst_dmem_n18422) );
NAND2_X1 MEM_stage_inst_dmem_U17083 ( .A1(MEM_stage_inst_dmem_n18420), .A2(MEM_stage_inst_dmem_n18419), .ZN(MEM_stage_inst_dmem_n10182) );
NAND2_X1 MEM_stage_inst_dmem_U17082 ( .A1(MEM_stage_inst_dmem_n18864), .A2(MEM_stage_inst_dmem_n18442), .ZN(MEM_stage_inst_dmem_n18419) );
NAND2_X1 MEM_stage_inst_dmem_U17081 ( .A1(MEM_stage_inst_dmem_ram_2955), .A2(MEM_stage_inst_dmem_n18441), .ZN(MEM_stage_inst_dmem_n18420) );
NAND2_X1 MEM_stage_inst_dmem_U17080 ( .A1(MEM_stage_inst_dmem_n18418), .A2(MEM_stage_inst_dmem_n18417), .ZN(MEM_stage_inst_dmem_n10183) );
NAND2_X1 MEM_stage_inst_dmem_U17079 ( .A1(MEM_stage_inst_dmem_n18861), .A2(MEM_stage_inst_dmem_n18442), .ZN(MEM_stage_inst_dmem_n18417) );
NAND2_X1 MEM_stage_inst_dmem_U17078 ( .A1(MEM_stage_inst_dmem_ram_2956), .A2(MEM_stage_inst_dmem_n18441), .ZN(MEM_stage_inst_dmem_n18418) );
NAND2_X1 MEM_stage_inst_dmem_U17077 ( .A1(MEM_stage_inst_dmem_n18416), .A2(MEM_stage_inst_dmem_n18415), .ZN(MEM_stage_inst_dmem_n10184) );
NAND2_X1 MEM_stage_inst_dmem_U17076 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n18442), .ZN(MEM_stage_inst_dmem_n18415) );
NAND2_X1 MEM_stage_inst_dmem_U17075 ( .A1(MEM_stage_inst_dmem_ram_2957), .A2(MEM_stage_inst_dmem_n18441), .ZN(MEM_stage_inst_dmem_n18416) );
NAND2_X1 MEM_stage_inst_dmem_U17074 ( .A1(MEM_stage_inst_dmem_n18414), .A2(MEM_stage_inst_dmem_n18413), .ZN(MEM_stage_inst_dmem_n10185) );
NAND2_X1 MEM_stage_inst_dmem_U17073 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n18442), .ZN(MEM_stage_inst_dmem_n18413) );
NAND2_X1 MEM_stage_inst_dmem_U17072 ( .A1(MEM_stage_inst_dmem_ram_2958), .A2(MEM_stage_inst_dmem_n18441), .ZN(MEM_stage_inst_dmem_n18414) );
NAND2_X1 MEM_stage_inst_dmem_U17071 ( .A1(MEM_stage_inst_dmem_n18412), .A2(MEM_stage_inst_dmem_n18411), .ZN(MEM_stage_inst_dmem_n10186) );
NAND2_X1 MEM_stage_inst_dmem_U17070 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n18442), .ZN(MEM_stage_inst_dmem_n18411) );
INV_X1 MEM_stage_inst_dmem_U17069 ( .A(MEM_stage_inst_dmem_n18441), .ZN(MEM_stage_inst_dmem_n18442) );
NAND2_X1 MEM_stage_inst_dmem_U17068 ( .A1(MEM_stage_inst_dmem_ram_2959), .A2(MEM_stage_inst_dmem_n18441), .ZN(MEM_stage_inst_dmem_n18412) );
NAND2_X1 MEM_stage_inst_dmem_U17067 ( .A1(MEM_stage_inst_dmem_n21179), .A2(MEM_stage_inst_dmem_n18683), .ZN(MEM_stage_inst_dmem_n18441) );
NAND2_X1 MEM_stage_inst_dmem_U17066 ( .A1(MEM_stage_inst_dmem_n18410), .A2(MEM_stage_inst_dmem_n18409), .ZN(MEM_stage_inst_dmem_n10187) );
NAND2_X1 MEM_stage_inst_dmem_U17065 ( .A1(MEM_stage_inst_dmem_n19275), .A2(MEM_stage_inst_dmem_n18408), .ZN(MEM_stage_inst_dmem_n18409) );
NAND2_X1 MEM_stage_inst_dmem_U17064 ( .A1(MEM_stage_inst_dmem_ram_2960), .A2(MEM_stage_inst_dmem_n18407), .ZN(MEM_stage_inst_dmem_n18410) );
NAND2_X1 MEM_stage_inst_dmem_U17063 ( .A1(MEM_stage_inst_dmem_n18406), .A2(MEM_stage_inst_dmem_n18405), .ZN(MEM_stage_inst_dmem_n10188) );
NAND2_X1 MEM_stage_inst_dmem_U17062 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n18408), .ZN(MEM_stage_inst_dmem_n18405) );
NAND2_X1 MEM_stage_inst_dmem_U17061 ( .A1(MEM_stage_inst_dmem_ram_2961), .A2(MEM_stage_inst_dmem_n18407), .ZN(MEM_stage_inst_dmem_n18406) );
NAND2_X1 MEM_stage_inst_dmem_U17060 ( .A1(MEM_stage_inst_dmem_n18404), .A2(MEM_stage_inst_dmem_n18403), .ZN(MEM_stage_inst_dmem_n10189) );
NAND2_X1 MEM_stage_inst_dmem_U17059 ( .A1(MEM_stage_inst_dmem_n16789), .A2(MEM_stage_inst_dmem_n18408), .ZN(MEM_stage_inst_dmem_n18403) );
NAND2_X1 MEM_stage_inst_dmem_U17058 ( .A1(MEM_stage_inst_dmem_ram_2962), .A2(MEM_stage_inst_dmem_n18407), .ZN(MEM_stage_inst_dmem_n18404) );
NAND2_X1 MEM_stage_inst_dmem_U17057 ( .A1(MEM_stage_inst_dmem_n18402), .A2(MEM_stage_inst_dmem_n18401), .ZN(MEM_stage_inst_dmem_n10190) );
NAND2_X1 MEM_stage_inst_dmem_U17056 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n18408), .ZN(MEM_stage_inst_dmem_n18401) );
NAND2_X1 MEM_stage_inst_dmem_U17055 ( .A1(MEM_stage_inst_dmem_ram_2963), .A2(MEM_stage_inst_dmem_n18407), .ZN(MEM_stage_inst_dmem_n18402) );
NAND2_X1 MEM_stage_inst_dmem_U17054 ( .A1(MEM_stage_inst_dmem_n18400), .A2(MEM_stage_inst_dmem_n18399), .ZN(MEM_stage_inst_dmem_n10191) );
NAND2_X1 MEM_stage_inst_dmem_U17053 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n18408), .ZN(MEM_stage_inst_dmem_n18399) );
NAND2_X1 MEM_stage_inst_dmem_U17052 ( .A1(MEM_stage_inst_dmem_ram_2964), .A2(MEM_stage_inst_dmem_n18407), .ZN(MEM_stage_inst_dmem_n18400) );
NAND2_X1 MEM_stage_inst_dmem_U17051 ( .A1(MEM_stage_inst_dmem_n18398), .A2(MEM_stage_inst_dmem_n18397), .ZN(MEM_stage_inst_dmem_n10192) );
NAND2_X1 MEM_stage_inst_dmem_U17050 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n18408), .ZN(MEM_stage_inst_dmem_n18397) );
NAND2_X1 MEM_stage_inst_dmem_U17049 ( .A1(MEM_stage_inst_dmem_ram_2965), .A2(MEM_stage_inst_dmem_n18407), .ZN(MEM_stage_inst_dmem_n18398) );
NAND2_X1 MEM_stage_inst_dmem_U17048 ( .A1(MEM_stage_inst_dmem_n18396), .A2(MEM_stage_inst_dmem_n18395), .ZN(MEM_stage_inst_dmem_n10193) );
NAND2_X1 MEM_stage_inst_dmem_U17047 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n18408), .ZN(MEM_stage_inst_dmem_n18395) );
NAND2_X1 MEM_stage_inst_dmem_U17046 ( .A1(MEM_stage_inst_dmem_ram_2966), .A2(MEM_stage_inst_dmem_n18407), .ZN(MEM_stage_inst_dmem_n18396) );
NAND2_X1 MEM_stage_inst_dmem_U17045 ( .A1(MEM_stage_inst_dmem_n18394), .A2(MEM_stage_inst_dmem_n18393), .ZN(MEM_stage_inst_dmem_n10194) );
NAND2_X1 MEM_stage_inst_dmem_U17044 ( .A1(MEM_stage_inst_dmem_n18875), .A2(MEM_stage_inst_dmem_n18408), .ZN(MEM_stage_inst_dmem_n18393) );
NAND2_X1 MEM_stage_inst_dmem_U17043 ( .A1(MEM_stage_inst_dmem_ram_2967), .A2(MEM_stage_inst_dmem_n18407), .ZN(MEM_stage_inst_dmem_n18394) );
NAND2_X1 MEM_stage_inst_dmem_U17042 ( .A1(MEM_stage_inst_dmem_n18392), .A2(MEM_stage_inst_dmem_n18391), .ZN(MEM_stage_inst_dmem_n10195) );
NAND2_X1 MEM_stage_inst_dmem_U17041 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n18408), .ZN(MEM_stage_inst_dmem_n18391) );
NAND2_X1 MEM_stage_inst_dmem_U17040 ( .A1(MEM_stage_inst_dmem_ram_2968), .A2(MEM_stage_inst_dmem_n18407), .ZN(MEM_stage_inst_dmem_n18392) );
NAND2_X1 MEM_stage_inst_dmem_U17039 ( .A1(MEM_stage_inst_dmem_n18390), .A2(MEM_stage_inst_dmem_n18389), .ZN(MEM_stage_inst_dmem_n10196) );
NAND2_X1 MEM_stage_inst_dmem_U17038 ( .A1(MEM_stage_inst_dmem_n19251), .A2(MEM_stage_inst_dmem_n18408), .ZN(MEM_stage_inst_dmem_n18389) );
NAND2_X1 MEM_stage_inst_dmem_U17037 ( .A1(MEM_stage_inst_dmem_ram_2969), .A2(MEM_stage_inst_dmem_n18407), .ZN(MEM_stage_inst_dmem_n18390) );
NAND2_X1 MEM_stage_inst_dmem_U17036 ( .A1(MEM_stage_inst_dmem_n18388), .A2(MEM_stage_inst_dmem_n18387), .ZN(MEM_stage_inst_dmem_n10197) );
NAND2_X1 MEM_stage_inst_dmem_U17035 ( .A1(MEM_stage_inst_dmem_n16769), .A2(MEM_stage_inst_dmem_n18408), .ZN(MEM_stage_inst_dmem_n18387) );
NAND2_X1 MEM_stage_inst_dmem_U17034 ( .A1(MEM_stage_inst_dmem_ram_2970), .A2(MEM_stage_inst_dmem_n18407), .ZN(MEM_stage_inst_dmem_n18388) );
NAND2_X1 MEM_stage_inst_dmem_U17033 ( .A1(MEM_stage_inst_dmem_n18386), .A2(MEM_stage_inst_dmem_n18385), .ZN(MEM_stage_inst_dmem_n10198) );
NAND2_X1 MEM_stage_inst_dmem_U17032 ( .A1(MEM_stage_inst_dmem_n20904), .A2(MEM_stage_inst_dmem_n18408), .ZN(MEM_stage_inst_dmem_n18385) );
NAND2_X1 MEM_stage_inst_dmem_U17031 ( .A1(MEM_stage_inst_dmem_ram_2971), .A2(MEM_stage_inst_dmem_n18407), .ZN(MEM_stage_inst_dmem_n18386) );
NAND2_X1 MEM_stage_inst_dmem_U17030 ( .A1(MEM_stage_inst_dmem_n18384), .A2(MEM_stage_inst_dmem_n18383), .ZN(MEM_stage_inst_dmem_n10199) );
NAND2_X1 MEM_stage_inst_dmem_U17029 ( .A1(MEM_stage_inst_dmem_n21474), .A2(MEM_stage_inst_dmem_n18408), .ZN(MEM_stage_inst_dmem_n18383) );
NAND2_X1 MEM_stage_inst_dmem_U17028 ( .A1(MEM_stage_inst_dmem_ram_2972), .A2(MEM_stage_inst_dmem_n18407), .ZN(MEM_stage_inst_dmem_n18384) );
NAND2_X1 MEM_stage_inst_dmem_U17027 ( .A1(MEM_stage_inst_dmem_n18382), .A2(MEM_stage_inst_dmem_n18381), .ZN(MEM_stage_inst_dmem_n10200) );
NAND2_X1 MEM_stage_inst_dmem_U17026 ( .A1(MEM_stage_inst_dmem_n19242), .A2(MEM_stage_inst_dmem_n18408), .ZN(MEM_stage_inst_dmem_n18381) );
NAND2_X1 MEM_stage_inst_dmem_U17025 ( .A1(MEM_stage_inst_dmem_ram_2973), .A2(MEM_stage_inst_dmem_n18407), .ZN(MEM_stage_inst_dmem_n18382) );
NAND2_X1 MEM_stage_inst_dmem_U17024 ( .A1(MEM_stage_inst_dmem_n18380), .A2(MEM_stage_inst_dmem_n18379), .ZN(MEM_stage_inst_dmem_n10201) );
NAND2_X1 MEM_stage_inst_dmem_U17023 ( .A1(MEM_stage_inst_dmem_n115), .A2(MEM_stage_inst_dmem_n18408), .ZN(MEM_stage_inst_dmem_n18379) );
NAND2_X1 MEM_stage_inst_dmem_U17022 ( .A1(MEM_stage_inst_dmem_ram_2974), .A2(MEM_stage_inst_dmem_n18407), .ZN(MEM_stage_inst_dmem_n18380) );
NAND2_X1 MEM_stage_inst_dmem_U17021 ( .A1(MEM_stage_inst_dmem_n18378), .A2(MEM_stage_inst_dmem_n18377), .ZN(MEM_stage_inst_dmem_n10202) );
NAND2_X1 MEM_stage_inst_dmem_U17020 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n18408), .ZN(MEM_stage_inst_dmem_n18377) );
INV_X1 MEM_stage_inst_dmem_U17019 ( .A(MEM_stage_inst_dmem_n18407), .ZN(MEM_stage_inst_dmem_n18408) );
NAND2_X1 MEM_stage_inst_dmem_U17018 ( .A1(MEM_stage_inst_dmem_ram_2975), .A2(MEM_stage_inst_dmem_n18407), .ZN(MEM_stage_inst_dmem_n18378) );
NAND2_X1 MEM_stage_inst_dmem_U17017 ( .A1(MEM_stage_inst_dmem_n21144), .A2(MEM_stage_inst_dmem_n18683), .ZN(MEM_stage_inst_dmem_n18407) );
NAND2_X1 MEM_stage_inst_dmem_U17016 ( .A1(MEM_stage_inst_dmem_n18376), .A2(MEM_stage_inst_dmem_n18375), .ZN(MEM_stage_inst_dmem_n10203) );
NAND2_X1 MEM_stage_inst_dmem_U17015 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n18374), .ZN(MEM_stage_inst_dmem_n18375) );
NAND2_X1 MEM_stage_inst_dmem_U17014 ( .A1(MEM_stage_inst_dmem_ram_2976), .A2(MEM_stage_inst_dmem_n18373), .ZN(MEM_stage_inst_dmem_n18376) );
NAND2_X1 MEM_stage_inst_dmem_U17013 ( .A1(MEM_stage_inst_dmem_n18372), .A2(MEM_stage_inst_dmem_n18371), .ZN(MEM_stage_inst_dmem_n10204) );
NAND2_X1 MEM_stage_inst_dmem_U17012 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n18374), .ZN(MEM_stage_inst_dmem_n18371) );
NAND2_X1 MEM_stage_inst_dmem_U17011 ( .A1(MEM_stage_inst_dmem_ram_2977), .A2(MEM_stage_inst_dmem_n18373), .ZN(MEM_stage_inst_dmem_n18372) );
NAND2_X1 MEM_stage_inst_dmem_U17010 ( .A1(MEM_stage_inst_dmem_n18370), .A2(MEM_stage_inst_dmem_n18369), .ZN(MEM_stage_inst_dmem_n10205) );
NAND2_X1 MEM_stage_inst_dmem_U17009 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n18374), .ZN(MEM_stage_inst_dmem_n18369) );
NAND2_X1 MEM_stage_inst_dmem_U17008 ( .A1(MEM_stage_inst_dmem_ram_2978), .A2(MEM_stage_inst_dmem_n18373), .ZN(MEM_stage_inst_dmem_n18370) );
NAND2_X1 MEM_stage_inst_dmem_U17007 ( .A1(MEM_stage_inst_dmem_n18368), .A2(MEM_stage_inst_dmem_n18367), .ZN(MEM_stage_inst_dmem_n10206) );
NAND2_X1 MEM_stage_inst_dmem_U17006 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n18374), .ZN(MEM_stage_inst_dmem_n18367) );
NAND2_X1 MEM_stage_inst_dmem_U17005 ( .A1(MEM_stage_inst_dmem_ram_2979), .A2(MEM_stage_inst_dmem_n18373), .ZN(MEM_stage_inst_dmem_n18368) );
NAND2_X1 MEM_stage_inst_dmem_U17004 ( .A1(MEM_stage_inst_dmem_n18366), .A2(MEM_stage_inst_dmem_n18365), .ZN(MEM_stage_inst_dmem_n10207) );
NAND2_X1 MEM_stage_inst_dmem_U17003 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n18374), .ZN(MEM_stage_inst_dmem_n18365) );
NAND2_X1 MEM_stage_inst_dmem_U17002 ( .A1(MEM_stage_inst_dmem_ram_2980), .A2(MEM_stage_inst_dmem_n18373), .ZN(MEM_stage_inst_dmem_n18366) );
NAND2_X1 MEM_stage_inst_dmem_U17001 ( .A1(MEM_stage_inst_dmem_n18364), .A2(MEM_stage_inst_dmem_n18363), .ZN(MEM_stage_inst_dmem_n10208) );
NAND2_X1 MEM_stage_inst_dmem_U17000 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n18374), .ZN(MEM_stage_inst_dmem_n18363) );
NAND2_X1 MEM_stage_inst_dmem_U16999 ( .A1(MEM_stage_inst_dmem_ram_2981), .A2(MEM_stage_inst_dmem_n18373), .ZN(MEM_stage_inst_dmem_n18364) );
NAND2_X1 MEM_stage_inst_dmem_U16998 ( .A1(MEM_stage_inst_dmem_n18362), .A2(MEM_stage_inst_dmem_n18361), .ZN(MEM_stage_inst_dmem_n10209) );
NAND2_X1 MEM_stage_inst_dmem_U16997 ( .A1(MEM_stage_inst_dmem_n21340), .A2(MEM_stage_inst_dmem_n18374), .ZN(MEM_stage_inst_dmem_n18361) );
NAND2_X1 MEM_stage_inst_dmem_U16996 ( .A1(MEM_stage_inst_dmem_ram_2982), .A2(MEM_stage_inst_dmem_n18373), .ZN(MEM_stage_inst_dmem_n18362) );
NAND2_X1 MEM_stage_inst_dmem_U16995 ( .A1(MEM_stage_inst_dmem_n18360), .A2(MEM_stage_inst_dmem_n18359), .ZN(MEM_stage_inst_dmem_n10210) );
NAND2_X1 MEM_stage_inst_dmem_U16994 ( .A1(MEM_stage_inst_dmem_n18), .A2(MEM_stage_inst_dmem_n18374), .ZN(MEM_stage_inst_dmem_n18359) );
NAND2_X1 MEM_stage_inst_dmem_U16993 ( .A1(MEM_stage_inst_dmem_ram_2983), .A2(MEM_stage_inst_dmem_n18373), .ZN(MEM_stage_inst_dmem_n18360) );
NAND2_X1 MEM_stage_inst_dmem_U16992 ( .A1(MEM_stage_inst_dmem_n18358), .A2(MEM_stage_inst_dmem_n18357), .ZN(MEM_stage_inst_dmem_n10211) );
NAND2_X1 MEM_stage_inst_dmem_U16991 ( .A1(MEM_stage_inst_dmem_n21335), .A2(MEM_stage_inst_dmem_n18374), .ZN(MEM_stage_inst_dmem_n18357) );
NAND2_X1 MEM_stage_inst_dmem_U16990 ( .A1(MEM_stage_inst_dmem_ram_2984), .A2(MEM_stage_inst_dmem_n18373), .ZN(MEM_stage_inst_dmem_n18358) );
NAND2_X1 MEM_stage_inst_dmem_U16989 ( .A1(MEM_stage_inst_dmem_n18356), .A2(MEM_stage_inst_dmem_n18355), .ZN(MEM_stage_inst_dmem_n10212) );
NAND2_X1 MEM_stage_inst_dmem_U16988 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n18374), .ZN(MEM_stage_inst_dmem_n18355) );
NAND2_X1 MEM_stage_inst_dmem_U16987 ( .A1(MEM_stage_inst_dmem_ram_2985), .A2(MEM_stage_inst_dmem_n18373), .ZN(MEM_stage_inst_dmem_n18356) );
NAND2_X1 MEM_stage_inst_dmem_U16986 ( .A1(MEM_stage_inst_dmem_n18354), .A2(MEM_stage_inst_dmem_n18353), .ZN(MEM_stage_inst_dmem_n10213) );
NAND2_X1 MEM_stage_inst_dmem_U16985 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n18374), .ZN(MEM_stage_inst_dmem_n18353) );
NAND2_X1 MEM_stage_inst_dmem_U16984 ( .A1(MEM_stage_inst_dmem_ram_2986), .A2(MEM_stage_inst_dmem_n18373), .ZN(MEM_stage_inst_dmem_n18354) );
NAND2_X1 MEM_stage_inst_dmem_U16983 ( .A1(MEM_stage_inst_dmem_n18352), .A2(MEM_stage_inst_dmem_n18351), .ZN(MEM_stage_inst_dmem_n10214) );
NAND2_X1 MEM_stage_inst_dmem_U16982 ( .A1(MEM_stage_inst_dmem_n14705), .A2(MEM_stage_inst_dmem_n18374), .ZN(MEM_stage_inst_dmem_n18351) );
NAND2_X1 MEM_stage_inst_dmem_U16981 ( .A1(MEM_stage_inst_dmem_ram_2987), .A2(MEM_stage_inst_dmem_n18373), .ZN(MEM_stage_inst_dmem_n18352) );
NAND2_X1 MEM_stage_inst_dmem_U16980 ( .A1(MEM_stage_inst_dmem_n18350), .A2(MEM_stage_inst_dmem_n18349), .ZN(MEM_stage_inst_dmem_n10215) );
NAND2_X1 MEM_stage_inst_dmem_U16979 ( .A1(MEM_stage_inst_dmem_n14702), .A2(MEM_stage_inst_dmem_n18374), .ZN(MEM_stage_inst_dmem_n18349) );
NAND2_X1 MEM_stage_inst_dmem_U16978 ( .A1(MEM_stage_inst_dmem_ram_2988), .A2(MEM_stage_inst_dmem_n18373), .ZN(MEM_stage_inst_dmem_n18350) );
NAND2_X1 MEM_stage_inst_dmem_U16977 ( .A1(MEM_stage_inst_dmem_n18348), .A2(MEM_stage_inst_dmem_n18347), .ZN(MEM_stage_inst_dmem_n10216) );
NAND2_X1 MEM_stage_inst_dmem_U16976 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n18374), .ZN(MEM_stage_inst_dmem_n18347) );
NAND2_X1 MEM_stage_inst_dmem_U16975 ( .A1(MEM_stage_inst_dmem_ram_2989), .A2(MEM_stage_inst_dmem_n18373), .ZN(MEM_stage_inst_dmem_n18348) );
NAND2_X1 MEM_stage_inst_dmem_U16974 ( .A1(MEM_stage_inst_dmem_n18346), .A2(MEM_stage_inst_dmem_n18345), .ZN(MEM_stage_inst_dmem_n10217) );
NAND2_X1 MEM_stage_inst_dmem_U16973 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n18374), .ZN(MEM_stage_inst_dmem_n18345) );
NAND2_X1 MEM_stage_inst_dmem_U16972 ( .A1(MEM_stage_inst_dmem_ram_2990), .A2(MEM_stage_inst_dmem_n18373), .ZN(MEM_stage_inst_dmem_n18346) );
NAND2_X1 MEM_stage_inst_dmem_U16971 ( .A1(MEM_stage_inst_dmem_n18344), .A2(MEM_stage_inst_dmem_n18343), .ZN(MEM_stage_inst_dmem_n10218) );
NAND2_X1 MEM_stage_inst_dmem_U16970 ( .A1(MEM_stage_inst_dmem_n21320), .A2(MEM_stage_inst_dmem_n18374), .ZN(MEM_stage_inst_dmem_n18343) );
NAND2_X1 MEM_stage_inst_dmem_U16969 ( .A1(MEM_stage_inst_dmem_ram_2991), .A2(MEM_stage_inst_dmem_n18373), .ZN(MEM_stage_inst_dmem_n18344) );
NAND2_X1 MEM_stage_inst_dmem_U16968 ( .A1(MEM_stage_inst_dmem_n21109), .A2(MEM_stage_inst_dmem_n18683), .ZN(MEM_stage_inst_dmem_n18373) );
NAND2_X1 MEM_stage_inst_dmem_U16967 ( .A1(MEM_stage_inst_dmem_n18342), .A2(MEM_stage_inst_dmem_n18341), .ZN(MEM_stage_inst_dmem_n10219) );
NAND2_X1 MEM_stage_inst_dmem_U16966 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n18340), .ZN(MEM_stage_inst_dmem_n18341) );
NAND2_X1 MEM_stage_inst_dmem_U16965 ( .A1(MEM_stage_inst_dmem_ram_2992), .A2(MEM_stage_inst_dmem_n18339), .ZN(MEM_stage_inst_dmem_n18342) );
NAND2_X1 MEM_stage_inst_dmem_U16964 ( .A1(MEM_stage_inst_dmem_n18338), .A2(MEM_stage_inst_dmem_n18337), .ZN(MEM_stage_inst_dmem_n10220) );
NAND2_X1 MEM_stage_inst_dmem_U16963 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n18340), .ZN(MEM_stage_inst_dmem_n18337) );
NAND2_X1 MEM_stage_inst_dmem_U16962 ( .A1(MEM_stage_inst_dmem_ram_2993), .A2(MEM_stage_inst_dmem_n18339), .ZN(MEM_stage_inst_dmem_n18338) );
NAND2_X1 MEM_stage_inst_dmem_U16961 ( .A1(MEM_stage_inst_dmem_n18336), .A2(MEM_stage_inst_dmem_n18335), .ZN(MEM_stage_inst_dmem_n10221) );
NAND2_X1 MEM_stage_inst_dmem_U16960 ( .A1(MEM_stage_inst_dmem_n18887), .A2(MEM_stage_inst_dmem_n18340), .ZN(MEM_stage_inst_dmem_n18335) );
NAND2_X1 MEM_stage_inst_dmem_U16959 ( .A1(MEM_stage_inst_dmem_ram_2994), .A2(MEM_stage_inst_dmem_n18339), .ZN(MEM_stage_inst_dmem_n18336) );
NAND2_X1 MEM_stage_inst_dmem_U16958 ( .A1(MEM_stage_inst_dmem_n18334), .A2(MEM_stage_inst_dmem_n18333), .ZN(MEM_stage_inst_dmem_n10222) );
NAND2_X1 MEM_stage_inst_dmem_U16957 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n18340), .ZN(MEM_stage_inst_dmem_n18333) );
NAND2_X1 MEM_stage_inst_dmem_U16956 ( .A1(MEM_stage_inst_dmem_ram_2995), .A2(MEM_stage_inst_dmem_n18339), .ZN(MEM_stage_inst_dmem_n18334) );
NAND2_X1 MEM_stage_inst_dmem_U16955 ( .A1(MEM_stage_inst_dmem_n18332), .A2(MEM_stage_inst_dmem_n18331), .ZN(MEM_stage_inst_dmem_n10223) );
NAND2_X1 MEM_stage_inst_dmem_U16954 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n18340), .ZN(MEM_stage_inst_dmem_n18331) );
NAND2_X1 MEM_stage_inst_dmem_U16953 ( .A1(MEM_stage_inst_dmem_ram_2996), .A2(MEM_stage_inst_dmem_n18339), .ZN(MEM_stage_inst_dmem_n18332) );
NAND2_X1 MEM_stage_inst_dmem_U16952 ( .A1(MEM_stage_inst_dmem_n18330), .A2(MEM_stage_inst_dmem_n18329), .ZN(MEM_stage_inst_dmem_n10224) );
NAND2_X1 MEM_stage_inst_dmem_U16951 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n18340), .ZN(MEM_stage_inst_dmem_n18329) );
NAND2_X1 MEM_stage_inst_dmem_U16950 ( .A1(MEM_stage_inst_dmem_ram_2997), .A2(MEM_stage_inst_dmem_n18339), .ZN(MEM_stage_inst_dmem_n18330) );
NAND2_X1 MEM_stage_inst_dmem_U16949 ( .A1(MEM_stage_inst_dmem_n18328), .A2(MEM_stage_inst_dmem_n18327), .ZN(MEM_stage_inst_dmem_n10225) );
NAND2_X1 MEM_stage_inst_dmem_U16948 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n18340), .ZN(MEM_stage_inst_dmem_n18327) );
NAND2_X1 MEM_stage_inst_dmem_U16947 ( .A1(MEM_stage_inst_dmem_ram_2998), .A2(MEM_stage_inst_dmem_n18339), .ZN(MEM_stage_inst_dmem_n18328) );
NAND2_X1 MEM_stage_inst_dmem_U16946 ( .A1(MEM_stage_inst_dmem_n18326), .A2(MEM_stage_inst_dmem_n18325), .ZN(MEM_stage_inst_dmem_n10226) );
NAND2_X1 MEM_stage_inst_dmem_U16945 ( .A1(MEM_stage_inst_dmem_n18875), .A2(MEM_stage_inst_dmem_n18340), .ZN(MEM_stage_inst_dmem_n18325) );
NAND2_X1 MEM_stage_inst_dmem_U16944 ( .A1(MEM_stage_inst_dmem_ram_2999), .A2(MEM_stage_inst_dmem_n18339), .ZN(MEM_stage_inst_dmem_n18326) );
NAND2_X1 MEM_stage_inst_dmem_U16943 ( .A1(MEM_stage_inst_dmem_n18324), .A2(MEM_stage_inst_dmem_n18323), .ZN(MEM_stage_inst_dmem_n10227) );
NAND2_X1 MEM_stage_inst_dmem_U16942 ( .A1(MEM_stage_inst_dmem_n111), .A2(MEM_stage_inst_dmem_n18340), .ZN(MEM_stage_inst_dmem_n18323) );
NAND2_X1 MEM_stage_inst_dmem_U16941 ( .A1(MEM_stage_inst_dmem_ram_3000), .A2(MEM_stage_inst_dmem_n18339), .ZN(MEM_stage_inst_dmem_n18324) );
NAND2_X1 MEM_stage_inst_dmem_U16940 ( .A1(MEM_stage_inst_dmem_n18322), .A2(MEM_stage_inst_dmem_n18321), .ZN(MEM_stage_inst_dmem_n10228) );
NAND2_X1 MEM_stage_inst_dmem_U16939 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n18340), .ZN(MEM_stage_inst_dmem_n18321) );
NAND2_X1 MEM_stage_inst_dmem_U16938 ( .A1(MEM_stage_inst_dmem_ram_3001), .A2(MEM_stage_inst_dmem_n18339), .ZN(MEM_stage_inst_dmem_n18322) );
NAND2_X1 MEM_stage_inst_dmem_U16937 ( .A1(MEM_stage_inst_dmem_n18320), .A2(MEM_stage_inst_dmem_n18319), .ZN(MEM_stage_inst_dmem_n10229) );
NAND2_X1 MEM_stage_inst_dmem_U16936 ( .A1(MEM_stage_inst_dmem_n18867), .A2(MEM_stage_inst_dmem_n18340), .ZN(MEM_stage_inst_dmem_n18319) );
NAND2_X1 MEM_stage_inst_dmem_U16935 ( .A1(MEM_stage_inst_dmem_ram_3002), .A2(MEM_stage_inst_dmem_n18339), .ZN(MEM_stage_inst_dmem_n18320) );
NAND2_X1 MEM_stage_inst_dmem_U16934 ( .A1(MEM_stage_inst_dmem_n18318), .A2(MEM_stage_inst_dmem_n18317), .ZN(MEM_stage_inst_dmem_n10230) );
NAND2_X1 MEM_stage_inst_dmem_U16933 ( .A1(MEM_stage_inst_dmem_n18864), .A2(MEM_stage_inst_dmem_n18340), .ZN(MEM_stage_inst_dmem_n18317) );
NAND2_X1 MEM_stage_inst_dmem_U16932 ( .A1(MEM_stage_inst_dmem_ram_3003), .A2(MEM_stage_inst_dmem_n18339), .ZN(MEM_stage_inst_dmem_n18318) );
NAND2_X1 MEM_stage_inst_dmem_U16931 ( .A1(MEM_stage_inst_dmem_n18316), .A2(MEM_stage_inst_dmem_n18315), .ZN(MEM_stage_inst_dmem_n10231) );
NAND2_X1 MEM_stage_inst_dmem_U16930 ( .A1(MEM_stage_inst_dmem_n18861), .A2(MEM_stage_inst_dmem_n18340), .ZN(MEM_stage_inst_dmem_n18315) );
NAND2_X1 MEM_stage_inst_dmem_U16929 ( .A1(MEM_stage_inst_dmem_ram_3004), .A2(MEM_stage_inst_dmem_n18339), .ZN(MEM_stage_inst_dmem_n18316) );
NAND2_X1 MEM_stage_inst_dmem_U16928 ( .A1(MEM_stage_inst_dmem_n18314), .A2(MEM_stage_inst_dmem_n18313), .ZN(MEM_stage_inst_dmem_n10232) );
NAND2_X1 MEM_stage_inst_dmem_U16927 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n18340), .ZN(MEM_stage_inst_dmem_n18313) );
NAND2_X1 MEM_stage_inst_dmem_U16926 ( .A1(MEM_stage_inst_dmem_ram_3005), .A2(MEM_stage_inst_dmem_n18339), .ZN(MEM_stage_inst_dmem_n18314) );
NAND2_X1 MEM_stage_inst_dmem_U16925 ( .A1(MEM_stage_inst_dmem_n18312), .A2(MEM_stage_inst_dmem_n18311), .ZN(MEM_stage_inst_dmem_n10233) );
NAND2_X1 MEM_stage_inst_dmem_U16924 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n18340), .ZN(MEM_stage_inst_dmem_n18311) );
NAND2_X1 MEM_stage_inst_dmem_U16923 ( .A1(MEM_stage_inst_dmem_ram_3006), .A2(MEM_stage_inst_dmem_n18339), .ZN(MEM_stage_inst_dmem_n18312) );
NAND2_X1 MEM_stage_inst_dmem_U16922 ( .A1(MEM_stage_inst_dmem_n18310), .A2(MEM_stage_inst_dmem_n18309), .ZN(MEM_stage_inst_dmem_n10234) );
NAND2_X1 MEM_stage_inst_dmem_U16921 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n18340), .ZN(MEM_stage_inst_dmem_n18309) );
INV_X1 MEM_stage_inst_dmem_U16920 ( .A(MEM_stage_inst_dmem_n18339), .ZN(MEM_stage_inst_dmem_n18340) );
NAND2_X1 MEM_stage_inst_dmem_U16919 ( .A1(MEM_stage_inst_dmem_ram_3007), .A2(MEM_stage_inst_dmem_n18339), .ZN(MEM_stage_inst_dmem_n18310) );
NAND2_X1 MEM_stage_inst_dmem_U16918 ( .A1(MEM_stage_inst_dmem_n21074), .A2(MEM_stage_inst_dmem_n18683), .ZN(MEM_stage_inst_dmem_n18339) );
NAND2_X1 MEM_stage_inst_dmem_U16917 ( .A1(MEM_stage_inst_dmem_n18308), .A2(MEM_stage_inst_dmem_n18307), .ZN(MEM_stage_inst_dmem_n10235) );
NAND2_X1 MEM_stage_inst_dmem_U16916 ( .A1(MEM_stage_inst_dmem_n20551), .A2(MEM_stage_inst_dmem_n18306), .ZN(MEM_stage_inst_dmem_n18307) );
NAND2_X1 MEM_stage_inst_dmem_U16915 ( .A1(MEM_stage_inst_dmem_ram_3008), .A2(MEM_stage_inst_dmem_n18305), .ZN(MEM_stage_inst_dmem_n18308) );
NAND2_X1 MEM_stage_inst_dmem_U16914 ( .A1(MEM_stage_inst_dmem_n18304), .A2(MEM_stage_inst_dmem_n18303), .ZN(MEM_stage_inst_dmem_n10236) );
NAND2_X1 MEM_stage_inst_dmem_U16913 ( .A1(MEM_stage_inst_dmem_n20547), .A2(MEM_stage_inst_dmem_n18306), .ZN(MEM_stage_inst_dmem_n18303) );
NAND2_X1 MEM_stage_inst_dmem_U16912 ( .A1(MEM_stage_inst_dmem_ram_3009), .A2(MEM_stage_inst_dmem_n18305), .ZN(MEM_stage_inst_dmem_n18304) );
NAND2_X1 MEM_stage_inst_dmem_U16911 ( .A1(MEM_stage_inst_dmem_n18302), .A2(MEM_stage_inst_dmem_n18301), .ZN(MEM_stage_inst_dmem_n10237) );
NAND2_X1 MEM_stage_inst_dmem_U16910 ( .A1(MEM_stage_inst_dmem_n20544), .A2(MEM_stage_inst_dmem_n18306), .ZN(MEM_stage_inst_dmem_n18301) );
NAND2_X1 MEM_stage_inst_dmem_U16909 ( .A1(MEM_stage_inst_dmem_ram_3010), .A2(MEM_stage_inst_dmem_n18305), .ZN(MEM_stage_inst_dmem_n18302) );
NAND2_X1 MEM_stage_inst_dmem_U16908 ( .A1(MEM_stage_inst_dmem_n18300), .A2(MEM_stage_inst_dmem_n18299), .ZN(MEM_stage_inst_dmem_n10238) );
NAND2_X1 MEM_stage_inst_dmem_U16907 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n18306), .ZN(MEM_stage_inst_dmem_n18299) );
NAND2_X1 MEM_stage_inst_dmem_U16906 ( .A1(MEM_stage_inst_dmem_ram_3011), .A2(MEM_stage_inst_dmem_n18305), .ZN(MEM_stage_inst_dmem_n18300) );
NAND2_X1 MEM_stage_inst_dmem_U16905 ( .A1(MEM_stage_inst_dmem_n18298), .A2(MEM_stage_inst_dmem_n18297), .ZN(MEM_stage_inst_dmem_n10239) );
NAND2_X1 MEM_stage_inst_dmem_U16904 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n18306), .ZN(MEM_stage_inst_dmem_n18297) );
NAND2_X1 MEM_stage_inst_dmem_U16903 ( .A1(MEM_stage_inst_dmem_ram_3012), .A2(MEM_stage_inst_dmem_n18305), .ZN(MEM_stage_inst_dmem_n18298) );
NAND2_X1 MEM_stage_inst_dmem_U16902 ( .A1(MEM_stage_inst_dmem_n18296), .A2(MEM_stage_inst_dmem_n18295), .ZN(MEM_stage_inst_dmem_n10240) );
NAND2_X1 MEM_stage_inst_dmem_U16901 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n18306), .ZN(MEM_stage_inst_dmem_n18295) );
NAND2_X1 MEM_stage_inst_dmem_U16900 ( .A1(MEM_stage_inst_dmem_ram_3013), .A2(MEM_stage_inst_dmem_n18305), .ZN(MEM_stage_inst_dmem_n18296) );
NAND2_X1 MEM_stage_inst_dmem_U16899 ( .A1(MEM_stage_inst_dmem_n18294), .A2(MEM_stage_inst_dmem_n18293), .ZN(MEM_stage_inst_dmem_n10241) );
NAND2_X1 MEM_stage_inst_dmem_U16898 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n18306), .ZN(MEM_stage_inst_dmem_n18293) );
NAND2_X1 MEM_stage_inst_dmem_U16897 ( .A1(MEM_stage_inst_dmem_ram_3014), .A2(MEM_stage_inst_dmem_n18305), .ZN(MEM_stage_inst_dmem_n18294) );
NAND2_X1 MEM_stage_inst_dmem_U16896 ( .A1(MEM_stage_inst_dmem_n18292), .A2(MEM_stage_inst_dmem_n18291), .ZN(MEM_stage_inst_dmem_n10242) );
NAND2_X1 MEM_stage_inst_dmem_U16895 ( .A1(MEM_stage_inst_dmem_n20530), .A2(MEM_stage_inst_dmem_n18306), .ZN(MEM_stage_inst_dmem_n18291) );
NAND2_X1 MEM_stage_inst_dmem_U16894 ( .A1(MEM_stage_inst_dmem_ram_3015), .A2(MEM_stage_inst_dmem_n18305), .ZN(MEM_stage_inst_dmem_n18292) );
NAND2_X1 MEM_stage_inst_dmem_U16893 ( .A1(MEM_stage_inst_dmem_n18290), .A2(MEM_stage_inst_dmem_n18289), .ZN(MEM_stage_inst_dmem_n10243) );
NAND2_X1 MEM_stage_inst_dmem_U16892 ( .A1(MEM_stage_inst_dmem_n20527), .A2(MEM_stage_inst_dmem_n18306), .ZN(MEM_stage_inst_dmem_n18289) );
NAND2_X1 MEM_stage_inst_dmem_U16891 ( .A1(MEM_stage_inst_dmem_ram_3016), .A2(MEM_stage_inst_dmem_n18305), .ZN(MEM_stage_inst_dmem_n18290) );
NAND2_X1 MEM_stage_inst_dmem_U16890 ( .A1(MEM_stage_inst_dmem_n18288), .A2(MEM_stage_inst_dmem_n18287), .ZN(MEM_stage_inst_dmem_n10244) );
NAND2_X1 MEM_stage_inst_dmem_U16889 ( .A1(MEM_stage_inst_dmem_n20524), .A2(MEM_stage_inst_dmem_n18306), .ZN(MEM_stage_inst_dmem_n18287) );
NAND2_X1 MEM_stage_inst_dmem_U16888 ( .A1(MEM_stage_inst_dmem_ram_3017), .A2(MEM_stage_inst_dmem_n18305), .ZN(MEM_stage_inst_dmem_n18288) );
NAND2_X1 MEM_stage_inst_dmem_U16887 ( .A1(MEM_stage_inst_dmem_n18286), .A2(MEM_stage_inst_dmem_n18285), .ZN(MEM_stage_inst_dmem_n10245) );
NAND2_X1 MEM_stage_inst_dmem_U16886 ( .A1(MEM_stage_inst_dmem_n20521), .A2(MEM_stage_inst_dmem_n18306), .ZN(MEM_stage_inst_dmem_n18285) );
NAND2_X1 MEM_stage_inst_dmem_U16885 ( .A1(MEM_stage_inst_dmem_ram_3018), .A2(MEM_stage_inst_dmem_n18305), .ZN(MEM_stage_inst_dmem_n18286) );
NAND2_X1 MEM_stage_inst_dmem_U16884 ( .A1(MEM_stage_inst_dmem_n18284), .A2(MEM_stage_inst_dmem_n18283), .ZN(MEM_stage_inst_dmem_n10246) );
NAND2_X1 MEM_stage_inst_dmem_U16883 ( .A1(MEM_stage_inst_dmem_n20518), .A2(MEM_stage_inst_dmem_n18306), .ZN(MEM_stage_inst_dmem_n18283) );
NAND2_X1 MEM_stage_inst_dmem_U16882 ( .A1(MEM_stage_inst_dmem_ram_3019), .A2(MEM_stage_inst_dmem_n18305), .ZN(MEM_stage_inst_dmem_n18284) );
NAND2_X1 MEM_stage_inst_dmem_U16881 ( .A1(MEM_stage_inst_dmem_n18282), .A2(MEM_stage_inst_dmem_n18281), .ZN(MEM_stage_inst_dmem_n10247) );
NAND2_X1 MEM_stage_inst_dmem_U16880 ( .A1(MEM_stage_inst_dmem_n20515), .A2(MEM_stage_inst_dmem_n18306), .ZN(MEM_stage_inst_dmem_n18281) );
NAND2_X1 MEM_stage_inst_dmem_U16879 ( .A1(MEM_stage_inst_dmem_ram_3020), .A2(MEM_stage_inst_dmem_n18305), .ZN(MEM_stage_inst_dmem_n18282) );
NAND2_X1 MEM_stage_inst_dmem_U16878 ( .A1(MEM_stage_inst_dmem_n18280), .A2(MEM_stage_inst_dmem_n18279), .ZN(MEM_stage_inst_dmem_n10248) );
NAND2_X1 MEM_stage_inst_dmem_U16877 ( .A1(MEM_stage_inst_dmem_n20512), .A2(MEM_stage_inst_dmem_n18306), .ZN(MEM_stage_inst_dmem_n18279) );
NAND2_X1 MEM_stage_inst_dmem_U16876 ( .A1(MEM_stage_inst_dmem_ram_3021), .A2(MEM_stage_inst_dmem_n18305), .ZN(MEM_stage_inst_dmem_n18280) );
NAND2_X1 MEM_stage_inst_dmem_U16875 ( .A1(MEM_stage_inst_dmem_n18278), .A2(MEM_stage_inst_dmem_n18277), .ZN(MEM_stage_inst_dmem_n10249) );
NAND2_X1 MEM_stage_inst_dmem_U16874 ( .A1(MEM_stage_inst_dmem_n20509), .A2(MEM_stage_inst_dmem_n18306), .ZN(MEM_stage_inst_dmem_n18277) );
NAND2_X1 MEM_stage_inst_dmem_U16873 ( .A1(MEM_stage_inst_dmem_ram_3022), .A2(MEM_stage_inst_dmem_n18305), .ZN(MEM_stage_inst_dmem_n18278) );
NAND2_X1 MEM_stage_inst_dmem_U16872 ( .A1(MEM_stage_inst_dmem_n18276), .A2(MEM_stage_inst_dmem_n18275), .ZN(MEM_stage_inst_dmem_n10250) );
NAND2_X1 MEM_stage_inst_dmem_U16871 ( .A1(MEM_stage_inst_dmem_n20506), .A2(MEM_stage_inst_dmem_n18306), .ZN(MEM_stage_inst_dmem_n18275) );
INV_X1 MEM_stage_inst_dmem_U16870 ( .A(MEM_stage_inst_dmem_n18305), .ZN(MEM_stage_inst_dmem_n18306) );
NAND2_X1 MEM_stage_inst_dmem_U16869 ( .A1(MEM_stage_inst_dmem_ram_3023), .A2(MEM_stage_inst_dmem_n18305), .ZN(MEM_stage_inst_dmem_n18276) );
NAND2_X1 MEM_stage_inst_dmem_U16868 ( .A1(MEM_stage_inst_dmem_n21039), .A2(MEM_stage_inst_dmem_n18683), .ZN(MEM_stage_inst_dmem_n18305) );
NAND2_X1 MEM_stage_inst_dmem_U16867 ( .A1(MEM_stage_inst_dmem_n18274), .A2(MEM_stage_inst_dmem_n18273), .ZN(MEM_stage_inst_dmem_n10251) );
NAND2_X1 MEM_stage_inst_dmem_U16866 ( .A1(MEM_stage_inst_dmem_n19275), .A2(MEM_stage_inst_dmem_n18272), .ZN(MEM_stage_inst_dmem_n18273) );
NAND2_X1 MEM_stage_inst_dmem_U16865 ( .A1(MEM_stage_inst_dmem_ram_3024), .A2(MEM_stage_inst_dmem_n18271), .ZN(MEM_stage_inst_dmem_n18274) );
NAND2_X1 MEM_stage_inst_dmem_U16864 ( .A1(MEM_stage_inst_dmem_n18270), .A2(MEM_stage_inst_dmem_n18269), .ZN(MEM_stage_inst_dmem_n10252) );
NAND2_X1 MEM_stage_inst_dmem_U16863 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n18272), .ZN(MEM_stage_inst_dmem_n18269) );
NAND2_X1 MEM_stage_inst_dmem_U16862 ( .A1(MEM_stage_inst_dmem_ram_3025), .A2(MEM_stage_inst_dmem_n18271), .ZN(MEM_stage_inst_dmem_n18270) );
NAND2_X1 MEM_stage_inst_dmem_U16861 ( .A1(MEM_stage_inst_dmem_n18268), .A2(MEM_stage_inst_dmem_n18267), .ZN(MEM_stage_inst_dmem_n10253) );
NAND2_X1 MEM_stage_inst_dmem_U16860 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n18272), .ZN(MEM_stage_inst_dmem_n18267) );
NAND2_X1 MEM_stage_inst_dmem_U16859 ( .A1(MEM_stage_inst_dmem_ram_3026), .A2(MEM_stage_inst_dmem_n18271), .ZN(MEM_stage_inst_dmem_n18268) );
NAND2_X1 MEM_stage_inst_dmem_U16858 ( .A1(MEM_stage_inst_dmem_n18266), .A2(MEM_stage_inst_dmem_n18265), .ZN(MEM_stage_inst_dmem_n10254) );
NAND2_X1 MEM_stage_inst_dmem_U16857 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n18272), .ZN(MEM_stage_inst_dmem_n18265) );
NAND2_X1 MEM_stage_inst_dmem_U16856 ( .A1(MEM_stage_inst_dmem_ram_3027), .A2(MEM_stage_inst_dmem_n18271), .ZN(MEM_stage_inst_dmem_n18266) );
NAND2_X1 MEM_stage_inst_dmem_U16855 ( .A1(MEM_stage_inst_dmem_n18264), .A2(MEM_stage_inst_dmem_n18263), .ZN(MEM_stage_inst_dmem_n10255) );
NAND2_X1 MEM_stage_inst_dmem_U16854 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n18272), .ZN(MEM_stage_inst_dmem_n18263) );
NAND2_X1 MEM_stage_inst_dmem_U16853 ( .A1(MEM_stage_inst_dmem_ram_3028), .A2(MEM_stage_inst_dmem_n18271), .ZN(MEM_stage_inst_dmem_n18264) );
NAND2_X1 MEM_stage_inst_dmem_U16852 ( .A1(MEM_stage_inst_dmem_n18262), .A2(MEM_stage_inst_dmem_n18261), .ZN(MEM_stage_inst_dmem_n10256) );
NAND2_X1 MEM_stage_inst_dmem_U16851 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n18272), .ZN(MEM_stage_inst_dmem_n18261) );
NAND2_X1 MEM_stage_inst_dmem_U16850 ( .A1(MEM_stage_inst_dmem_ram_3029), .A2(MEM_stage_inst_dmem_n18271), .ZN(MEM_stage_inst_dmem_n18262) );
NAND2_X1 MEM_stage_inst_dmem_U16849 ( .A1(MEM_stage_inst_dmem_n18260), .A2(MEM_stage_inst_dmem_n18259), .ZN(MEM_stage_inst_dmem_n10257) );
NAND2_X1 MEM_stage_inst_dmem_U16848 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n18272), .ZN(MEM_stage_inst_dmem_n18259) );
NAND2_X1 MEM_stage_inst_dmem_U16847 ( .A1(MEM_stage_inst_dmem_ram_3030), .A2(MEM_stage_inst_dmem_n18271), .ZN(MEM_stage_inst_dmem_n18260) );
NAND2_X1 MEM_stage_inst_dmem_U16846 ( .A1(MEM_stage_inst_dmem_n18258), .A2(MEM_stage_inst_dmem_n18257), .ZN(MEM_stage_inst_dmem_n10258) );
NAND2_X1 MEM_stage_inst_dmem_U16845 ( .A1(MEM_stage_inst_dmem_n20530), .A2(MEM_stage_inst_dmem_n18272), .ZN(MEM_stage_inst_dmem_n18257) );
NAND2_X1 MEM_stage_inst_dmem_U16844 ( .A1(MEM_stage_inst_dmem_ram_3031), .A2(MEM_stage_inst_dmem_n18271), .ZN(MEM_stage_inst_dmem_n18258) );
NAND2_X1 MEM_stage_inst_dmem_U16843 ( .A1(MEM_stage_inst_dmem_n18256), .A2(MEM_stage_inst_dmem_n18255), .ZN(MEM_stage_inst_dmem_n10259) );
NAND2_X1 MEM_stage_inst_dmem_U16842 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n18272), .ZN(MEM_stage_inst_dmem_n18255) );
NAND2_X1 MEM_stage_inst_dmem_U16841 ( .A1(MEM_stage_inst_dmem_ram_3032), .A2(MEM_stage_inst_dmem_n18271), .ZN(MEM_stage_inst_dmem_n18256) );
NAND2_X1 MEM_stage_inst_dmem_U16840 ( .A1(MEM_stage_inst_dmem_n18254), .A2(MEM_stage_inst_dmem_n18253), .ZN(MEM_stage_inst_dmem_n10260) );
NAND2_X1 MEM_stage_inst_dmem_U16839 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n18272), .ZN(MEM_stage_inst_dmem_n18253) );
NAND2_X1 MEM_stage_inst_dmem_U16838 ( .A1(MEM_stage_inst_dmem_ram_3033), .A2(MEM_stage_inst_dmem_n18271), .ZN(MEM_stage_inst_dmem_n18254) );
NAND2_X1 MEM_stage_inst_dmem_U16837 ( .A1(MEM_stage_inst_dmem_n18252), .A2(MEM_stage_inst_dmem_n18251), .ZN(MEM_stage_inst_dmem_n10261) );
NAND2_X1 MEM_stage_inst_dmem_U16836 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n18272), .ZN(MEM_stage_inst_dmem_n18251) );
NAND2_X1 MEM_stage_inst_dmem_U16835 ( .A1(MEM_stage_inst_dmem_ram_3034), .A2(MEM_stage_inst_dmem_n18271), .ZN(MEM_stage_inst_dmem_n18252) );
NAND2_X1 MEM_stage_inst_dmem_U16834 ( .A1(MEM_stage_inst_dmem_n18250), .A2(MEM_stage_inst_dmem_n18249), .ZN(MEM_stage_inst_dmem_n10262) );
NAND2_X1 MEM_stage_inst_dmem_U16833 ( .A1(MEM_stage_inst_dmem_n14705), .A2(MEM_stage_inst_dmem_n18272), .ZN(MEM_stage_inst_dmem_n18249) );
NAND2_X1 MEM_stage_inst_dmem_U16832 ( .A1(MEM_stage_inst_dmem_ram_3035), .A2(MEM_stage_inst_dmem_n18271), .ZN(MEM_stage_inst_dmem_n18250) );
NAND2_X1 MEM_stage_inst_dmem_U16831 ( .A1(MEM_stage_inst_dmem_n18248), .A2(MEM_stage_inst_dmem_n18247), .ZN(MEM_stage_inst_dmem_n10263) );
NAND2_X1 MEM_stage_inst_dmem_U16830 ( .A1(MEM_stage_inst_dmem_n14702), .A2(MEM_stage_inst_dmem_n18272), .ZN(MEM_stage_inst_dmem_n18247) );
NAND2_X1 MEM_stage_inst_dmem_U16829 ( .A1(MEM_stage_inst_dmem_ram_3036), .A2(MEM_stage_inst_dmem_n18271), .ZN(MEM_stage_inst_dmem_n18248) );
NAND2_X1 MEM_stage_inst_dmem_U16828 ( .A1(MEM_stage_inst_dmem_n18246), .A2(MEM_stage_inst_dmem_n18245), .ZN(MEM_stage_inst_dmem_n10264) );
NAND2_X1 MEM_stage_inst_dmem_U16827 ( .A1(MEM_stage_inst_dmem_n19242), .A2(MEM_stage_inst_dmem_n18272), .ZN(MEM_stage_inst_dmem_n18245) );
NAND2_X1 MEM_stage_inst_dmem_U16826 ( .A1(MEM_stage_inst_dmem_ram_3037), .A2(MEM_stage_inst_dmem_n18271), .ZN(MEM_stage_inst_dmem_n18246) );
NAND2_X1 MEM_stage_inst_dmem_U16825 ( .A1(MEM_stage_inst_dmem_n18244), .A2(MEM_stage_inst_dmem_n18243), .ZN(MEM_stage_inst_dmem_n10265) );
NAND2_X1 MEM_stage_inst_dmem_U16824 ( .A1(MEM_stage_inst_dmem_n115), .A2(MEM_stage_inst_dmem_n18272), .ZN(MEM_stage_inst_dmem_n18243) );
NAND2_X1 MEM_stage_inst_dmem_U16823 ( .A1(MEM_stage_inst_dmem_ram_3038), .A2(MEM_stage_inst_dmem_n18271), .ZN(MEM_stage_inst_dmem_n18244) );
NAND2_X1 MEM_stage_inst_dmem_U16822 ( .A1(MEM_stage_inst_dmem_n18242), .A2(MEM_stage_inst_dmem_n18241), .ZN(MEM_stage_inst_dmem_n10266) );
NAND2_X1 MEM_stage_inst_dmem_U16821 ( .A1(MEM_stage_inst_dmem_n15110), .A2(MEM_stage_inst_dmem_n18272), .ZN(MEM_stage_inst_dmem_n18241) );
INV_X1 MEM_stage_inst_dmem_U16820 ( .A(MEM_stage_inst_dmem_n18271), .ZN(MEM_stage_inst_dmem_n18272) );
NAND2_X1 MEM_stage_inst_dmem_U16819 ( .A1(MEM_stage_inst_dmem_ram_3039), .A2(MEM_stage_inst_dmem_n18271), .ZN(MEM_stage_inst_dmem_n18242) );
NAND2_X1 MEM_stage_inst_dmem_U16818 ( .A1(MEM_stage_inst_dmem_n21004), .A2(MEM_stage_inst_dmem_n18683), .ZN(MEM_stage_inst_dmem_n18271) );
NAND2_X1 MEM_stage_inst_dmem_U16817 ( .A1(MEM_stage_inst_dmem_n18240), .A2(MEM_stage_inst_dmem_n18239), .ZN(MEM_stage_inst_dmem_n10267) );
NAND2_X1 MEM_stage_inst_dmem_U16816 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n18238), .ZN(MEM_stage_inst_dmem_n18239) );
NAND2_X1 MEM_stage_inst_dmem_U16815 ( .A1(MEM_stage_inst_dmem_ram_3040), .A2(MEM_stage_inst_dmem_n18237), .ZN(MEM_stage_inst_dmem_n18240) );
NAND2_X1 MEM_stage_inst_dmem_U16814 ( .A1(MEM_stage_inst_dmem_n18236), .A2(MEM_stage_inst_dmem_n18235), .ZN(MEM_stage_inst_dmem_n10268) );
NAND2_X1 MEM_stage_inst_dmem_U16813 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n18238), .ZN(MEM_stage_inst_dmem_n18235) );
NAND2_X1 MEM_stage_inst_dmem_U16812 ( .A1(MEM_stage_inst_dmem_ram_3041), .A2(MEM_stage_inst_dmem_n18237), .ZN(MEM_stage_inst_dmem_n18236) );
NAND2_X1 MEM_stage_inst_dmem_U16811 ( .A1(MEM_stage_inst_dmem_n18234), .A2(MEM_stage_inst_dmem_n18233), .ZN(MEM_stage_inst_dmem_n10269) );
NAND2_X1 MEM_stage_inst_dmem_U16810 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n18238), .ZN(MEM_stage_inst_dmem_n18233) );
NAND2_X1 MEM_stage_inst_dmem_U16809 ( .A1(MEM_stage_inst_dmem_ram_3042), .A2(MEM_stage_inst_dmem_n18237), .ZN(MEM_stage_inst_dmem_n18234) );
NAND2_X1 MEM_stage_inst_dmem_U16808 ( .A1(MEM_stage_inst_dmem_n18232), .A2(MEM_stage_inst_dmem_n18231), .ZN(MEM_stage_inst_dmem_n10270) );
NAND2_X1 MEM_stage_inst_dmem_U16807 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n18238), .ZN(MEM_stage_inst_dmem_n18231) );
NAND2_X1 MEM_stage_inst_dmem_U16806 ( .A1(MEM_stage_inst_dmem_ram_3043), .A2(MEM_stage_inst_dmem_n18237), .ZN(MEM_stage_inst_dmem_n18232) );
NAND2_X1 MEM_stage_inst_dmem_U16805 ( .A1(MEM_stage_inst_dmem_n18230), .A2(MEM_stage_inst_dmem_n18229), .ZN(MEM_stage_inst_dmem_n10271) );
NAND2_X1 MEM_stage_inst_dmem_U16804 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n18238), .ZN(MEM_stage_inst_dmem_n18229) );
NAND2_X1 MEM_stage_inst_dmem_U16803 ( .A1(MEM_stage_inst_dmem_ram_3044), .A2(MEM_stage_inst_dmem_n18237), .ZN(MEM_stage_inst_dmem_n18230) );
NAND2_X1 MEM_stage_inst_dmem_U16802 ( .A1(MEM_stage_inst_dmem_n18228), .A2(MEM_stage_inst_dmem_n18227), .ZN(MEM_stage_inst_dmem_n10272) );
NAND2_X1 MEM_stage_inst_dmem_U16801 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n18238), .ZN(MEM_stage_inst_dmem_n18227) );
NAND2_X1 MEM_stage_inst_dmem_U16800 ( .A1(MEM_stage_inst_dmem_ram_3045), .A2(MEM_stage_inst_dmem_n18237), .ZN(MEM_stage_inst_dmem_n18228) );
NAND2_X1 MEM_stage_inst_dmem_U16799 ( .A1(MEM_stage_inst_dmem_n18226), .A2(MEM_stage_inst_dmem_n18225), .ZN(MEM_stage_inst_dmem_n10273) );
NAND2_X1 MEM_stage_inst_dmem_U16798 ( .A1(MEM_stage_inst_dmem_n21340), .A2(MEM_stage_inst_dmem_n18238), .ZN(MEM_stage_inst_dmem_n18225) );
NAND2_X1 MEM_stage_inst_dmem_U16797 ( .A1(MEM_stage_inst_dmem_ram_3046), .A2(MEM_stage_inst_dmem_n18237), .ZN(MEM_stage_inst_dmem_n18226) );
NAND2_X1 MEM_stage_inst_dmem_U16796 ( .A1(MEM_stage_inst_dmem_n18224), .A2(MEM_stage_inst_dmem_n18223), .ZN(MEM_stage_inst_dmem_n10274) );
NAND2_X1 MEM_stage_inst_dmem_U16795 ( .A1(MEM_stage_inst_dmem_n17), .A2(MEM_stage_inst_dmem_n18238), .ZN(MEM_stage_inst_dmem_n18223) );
NAND2_X1 MEM_stage_inst_dmem_U16794 ( .A1(MEM_stage_inst_dmem_ram_3047), .A2(MEM_stage_inst_dmem_n18237), .ZN(MEM_stage_inst_dmem_n18224) );
NAND2_X1 MEM_stage_inst_dmem_U16793 ( .A1(MEM_stage_inst_dmem_n18222), .A2(MEM_stage_inst_dmem_n18221), .ZN(MEM_stage_inst_dmem_n10275) );
NAND2_X1 MEM_stage_inst_dmem_U16792 ( .A1(MEM_stage_inst_dmem_n21335), .A2(MEM_stage_inst_dmem_n18238), .ZN(MEM_stage_inst_dmem_n18221) );
NAND2_X1 MEM_stage_inst_dmem_U16791 ( .A1(MEM_stage_inst_dmem_ram_3048), .A2(MEM_stage_inst_dmem_n18237), .ZN(MEM_stage_inst_dmem_n18222) );
NAND2_X1 MEM_stage_inst_dmem_U16790 ( .A1(MEM_stage_inst_dmem_n18220), .A2(MEM_stage_inst_dmem_n18219), .ZN(MEM_stage_inst_dmem_n10276) );
NAND2_X1 MEM_stage_inst_dmem_U16789 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n18238), .ZN(MEM_stage_inst_dmem_n18219) );
NAND2_X1 MEM_stage_inst_dmem_U16788 ( .A1(MEM_stage_inst_dmem_ram_3049), .A2(MEM_stage_inst_dmem_n18237), .ZN(MEM_stage_inst_dmem_n18220) );
NAND2_X1 MEM_stage_inst_dmem_U16787 ( .A1(MEM_stage_inst_dmem_n18218), .A2(MEM_stage_inst_dmem_n18217), .ZN(MEM_stage_inst_dmem_n10277) );
NAND2_X1 MEM_stage_inst_dmem_U16786 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n18238), .ZN(MEM_stage_inst_dmem_n18217) );
NAND2_X1 MEM_stage_inst_dmem_U16785 ( .A1(MEM_stage_inst_dmem_ram_3050), .A2(MEM_stage_inst_dmem_n18237), .ZN(MEM_stage_inst_dmem_n18218) );
NAND2_X1 MEM_stage_inst_dmem_U16784 ( .A1(MEM_stage_inst_dmem_n18216), .A2(MEM_stage_inst_dmem_n18215), .ZN(MEM_stage_inst_dmem_n10278) );
NAND2_X1 MEM_stage_inst_dmem_U16783 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n18238), .ZN(MEM_stage_inst_dmem_n18215) );
NAND2_X1 MEM_stage_inst_dmem_U16782 ( .A1(MEM_stage_inst_dmem_ram_3051), .A2(MEM_stage_inst_dmem_n18237), .ZN(MEM_stage_inst_dmem_n18216) );
NAND2_X1 MEM_stage_inst_dmem_U16781 ( .A1(MEM_stage_inst_dmem_n18214), .A2(MEM_stage_inst_dmem_n18213), .ZN(MEM_stage_inst_dmem_n10279) );
NAND2_X1 MEM_stage_inst_dmem_U16780 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n18238), .ZN(MEM_stage_inst_dmem_n18213) );
NAND2_X1 MEM_stage_inst_dmem_U16779 ( .A1(MEM_stage_inst_dmem_ram_3052), .A2(MEM_stage_inst_dmem_n18237), .ZN(MEM_stage_inst_dmem_n18214) );
NAND2_X1 MEM_stage_inst_dmem_U16778 ( .A1(MEM_stage_inst_dmem_n18212), .A2(MEM_stage_inst_dmem_n18211), .ZN(MEM_stage_inst_dmem_n10280) );
NAND2_X1 MEM_stage_inst_dmem_U16777 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n18238), .ZN(MEM_stage_inst_dmem_n18211) );
NAND2_X1 MEM_stage_inst_dmem_U16776 ( .A1(MEM_stage_inst_dmem_ram_3053), .A2(MEM_stage_inst_dmem_n18237), .ZN(MEM_stage_inst_dmem_n18212) );
NAND2_X1 MEM_stage_inst_dmem_U16775 ( .A1(MEM_stage_inst_dmem_n18210), .A2(MEM_stage_inst_dmem_n18209), .ZN(MEM_stage_inst_dmem_n10281) );
NAND2_X1 MEM_stage_inst_dmem_U16774 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n18238), .ZN(MEM_stage_inst_dmem_n18209) );
NAND2_X1 MEM_stage_inst_dmem_U16773 ( .A1(MEM_stage_inst_dmem_ram_3054), .A2(MEM_stage_inst_dmem_n18237), .ZN(MEM_stage_inst_dmem_n18210) );
NAND2_X1 MEM_stage_inst_dmem_U16772 ( .A1(MEM_stage_inst_dmem_n18208), .A2(MEM_stage_inst_dmem_n18207), .ZN(MEM_stage_inst_dmem_n10282) );
NAND2_X1 MEM_stage_inst_dmem_U16771 ( .A1(MEM_stage_inst_dmem_n21320), .A2(MEM_stage_inst_dmem_n18238), .ZN(MEM_stage_inst_dmem_n18207) );
INV_X1 MEM_stage_inst_dmem_U16770 ( .A(MEM_stage_inst_dmem_n18237), .ZN(MEM_stage_inst_dmem_n18238) );
NAND2_X1 MEM_stage_inst_dmem_U16769 ( .A1(MEM_stage_inst_dmem_ram_3055), .A2(MEM_stage_inst_dmem_n18237), .ZN(MEM_stage_inst_dmem_n18208) );
NAND2_X1 MEM_stage_inst_dmem_U16768 ( .A1(MEM_stage_inst_dmem_n20969), .A2(MEM_stage_inst_dmem_n18683), .ZN(MEM_stage_inst_dmem_n18237) );
NAND2_X1 MEM_stage_inst_dmem_U16767 ( .A1(MEM_stage_inst_dmem_n18206), .A2(MEM_stage_inst_dmem_n18205), .ZN(MEM_stage_inst_dmem_n10283) );
NAND2_X1 MEM_stage_inst_dmem_U16766 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n18204), .ZN(MEM_stage_inst_dmem_n18205) );
NAND2_X1 MEM_stage_inst_dmem_U16765 ( .A1(MEM_stage_inst_dmem_ram_3056), .A2(MEM_stage_inst_dmem_n18203), .ZN(MEM_stage_inst_dmem_n18206) );
NAND2_X1 MEM_stage_inst_dmem_U16764 ( .A1(MEM_stage_inst_dmem_n18202), .A2(MEM_stage_inst_dmem_n18201), .ZN(MEM_stage_inst_dmem_n10284) );
NAND2_X1 MEM_stage_inst_dmem_U16763 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n18204), .ZN(MEM_stage_inst_dmem_n18201) );
NAND2_X1 MEM_stage_inst_dmem_U16762 ( .A1(MEM_stage_inst_dmem_ram_3057), .A2(MEM_stage_inst_dmem_n18203), .ZN(MEM_stage_inst_dmem_n18202) );
NAND2_X1 MEM_stage_inst_dmem_U16761 ( .A1(MEM_stage_inst_dmem_n18200), .A2(MEM_stage_inst_dmem_n18199), .ZN(MEM_stage_inst_dmem_n10285) );
NAND2_X1 MEM_stage_inst_dmem_U16760 ( .A1(MEM_stage_inst_dmem_n18887), .A2(MEM_stage_inst_dmem_n18204), .ZN(MEM_stage_inst_dmem_n18199) );
NAND2_X1 MEM_stage_inst_dmem_U16759 ( .A1(MEM_stage_inst_dmem_ram_3058), .A2(MEM_stage_inst_dmem_n18203), .ZN(MEM_stage_inst_dmem_n18200) );
NAND2_X1 MEM_stage_inst_dmem_U16758 ( .A1(MEM_stage_inst_dmem_n18198), .A2(MEM_stage_inst_dmem_n18197), .ZN(MEM_stage_inst_dmem_n10286) );
NAND2_X1 MEM_stage_inst_dmem_U16757 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n18204), .ZN(MEM_stage_inst_dmem_n18197) );
NAND2_X1 MEM_stage_inst_dmem_U16756 ( .A1(MEM_stage_inst_dmem_ram_3059), .A2(MEM_stage_inst_dmem_n18203), .ZN(MEM_stage_inst_dmem_n18198) );
NAND2_X1 MEM_stage_inst_dmem_U16755 ( .A1(MEM_stage_inst_dmem_n18196), .A2(MEM_stage_inst_dmem_n18195), .ZN(MEM_stage_inst_dmem_n10287) );
NAND2_X1 MEM_stage_inst_dmem_U16754 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n18204), .ZN(MEM_stage_inst_dmem_n18195) );
NAND2_X1 MEM_stage_inst_dmem_U16753 ( .A1(MEM_stage_inst_dmem_ram_3060), .A2(MEM_stage_inst_dmem_n18203), .ZN(MEM_stage_inst_dmem_n18196) );
NAND2_X1 MEM_stage_inst_dmem_U16752 ( .A1(MEM_stage_inst_dmem_n18194), .A2(MEM_stage_inst_dmem_n18193), .ZN(MEM_stage_inst_dmem_n10288) );
NAND2_X1 MEM_stage_inst_dmem_U16751 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n18204), .ZN(MEM_stage_inst_dmem_n18193) );
NAND2_X1 MEM_stage_inst_dmem_U16750 ( .A1(MEM_stage_inst_dmem_ram_3061), .A2(MEM_stage_inst_dmem_n18203), .ZN(MEM_stage_inst_dmem_n18194) );
NAND2_X1 MEM_stage_inst_dmem_U16749 ( .A1(MEM_stage_inst_dmem_n18192), .A2(MEM_stage_inst_dmem_n18191), .ZN(MEM_stage_inst_dmem_n10289) );
NAND2_X1 MEM_stage_inst_dmem_U16748 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n18204), .ZN(MEM_stage_inst_dmem_n18191) );
NAND2_X1 MEM_stage_inst_dmem_U16747 ( .A1(MEM_stage_inst_dmem_ram_3062), .A2(MEM_stage_inst_dmem_n18203), .ZN(MEM_stage_inst_dmem_n18192) );
NAND2_X1 MEM_stage_inst_dmem_U16746 ( .A1(MEM_stage_inst_dmem_n18190), .A2(MEM_stage_inst_dmem_n18189), .ZN(MEM_stage_inst_dmem_n10290) );
NAND2_X1 MEM_stage_inst_dmem_U16745 ( .A1(MEM_stage_inst_dmem_n18875), .A2(MEM_stage_inst_dmem_n18204), .ZN(MEM_stage_inst_dmem_n18189) );
NAND2_X1 MEM_stage_inst_dmem_U16744 ( .A1(MEM_stage_inst_dmem_ram_3063), .A2(MEM_stage_inst_dmem_n18203), .ZN(MEM_stage_inst_dmem_n18190) );
NAND2_X1 MEM_stage_inst_dmem_U16743 ( .A1(MEM_stage_inst_dmem_n18188), .A2(MEM_stage_inst_dmem_n18187), .ZN(MEM_stage_inst_dmem_n10291) );
NAND2_X1 MEM_stage_inst_dmem_U16742 ( .A1(MEM_stage_inst_dmem_n111), .A2(MEM_stage_inst_dmem_n18204), .ZN(MEM_stage_inst_dmem_n18187) );
NAND2_X1 MEM_stage_inst_dmem_U16741 ( .A1(MEM_stage_inst_dmem_ram_3064), .A2(MEM_stage_inst_dmem_n18203), .ZN(MEM_stage_inst_dmem_n18188) );
NAND2_X1 MEM_stage_inst_dmem_U16740 ( .A1(MEM_stage_inst_dmem_n18186), .A2(MEM_stage_inst_dmem_n18185), .ZN(MEM_stage_inst_dmem_n10292) );
NAND2_X1 MEM_stage_inst_dmem_U16739 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n18204), .ZN(MEM_stage_inst_dmem_n18185) );
NAND2_X1 MEM_stage_inst_dmem_U16738 ( .A1(MEM_stage_inst_dmem_ram_3065), .A2(MEM_stage_inst_dmem_n18203), .ZN(MEM_stage_inst_dmem_n18186) );
NAND2_X1 MEM_stage_inst_dmem_U16737 ( .A1(MEM_stage_inst_dmem_n18184), .A2(MEM_stage_inst_dmem_n18183), .ZN(MEM_stage_inst_dmem_n10293) );
NAND2_X1 MEM_stage_inst_dmem_U16736 ( .A1(MEM_stage_inst_dmem_n18867), .A2(MEM_stage_inst_dmem_n18204), .ZN(MEM_stage_inst_dmem_n18183) );
NAND2_X1 MEM_stage_inst_dmem_U16735 ( .A1(MEM_stage_inst_dmem_ram_3066), .A2(MEM_stage_inst_dmem_n18203), .ZN(MEM_stage_inst_dmem_n18184) );
NAND2_X1 MEM_stage_inst_dmem_U16734 ( .A1(MEM_stage_inst_dmem_n18182), .A2(MEM_stage_inst_dmem_n18181), .ZN(MEM_stage_inst_dmem_n10294) );
NAND2_X1 MEM_stage_inst_dmem_U16733 ( .A1(MEM_stage_inst_dmem_n18864), .A2(MEM_stage_inst_dmem_n18204), .ZN(MEM_stage_inst_dmem_n18181) );
NAND2_X1 MEM_stage_inst_dmem_U16732 ( .A1(MEM_stage_inst_dmem_ram_3067), .A2(MEM_stage_inst_dmem_n18203), .ZN(MEM_stage_inst_dmem_n18182) );
NAND2_X1 MEM_stage_inst_dmem_U16731 ( .A1(MEM_stage_inst_dmem_n18180), .A2(MEM_stage_inst_dmem_n18179), .ZN(MEM_stage_inst_dmem_n10295) );
NAND2_X1 MEM_stage_inst_dmem_U16730 ( .A1(MEM_stage_inst_dmem_n18861), .A2(MEM_stage_inst_dmem_n18204), .ZN(MEM_stage_inst_dmem_n18179) );
NAND2_X1 MEM_stage_inst_dmem_U16729 ( .A1(MEM_stage_inst_dmem_ram_3068), .A2(MEM_stage_inst_dmem_n18203), .ZN(MEM_stage_inst_dmem_n18180) );
NAND2_X1 MEM_stage_inst_dmem_U16728 ( .A1(MEM_stage_inst_dmem_n18178), .A2(MEM_stage_inst_dmem_n18177), .ZN(MEM_stage_inst_dmem_n10296) );
NAND2_X1 MEM_stage_inst_dmem_U16727 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n18204), .ZN(MEM_stage_inst_dmem_n18177) );
NAND2_X1 MEM_stage_inst_dmem_U16726 ( .A1(MEM_stage_inst_dmem_ram_3069), .A2(MEM_stage_inst_dmem_n18203), .ZN(MEM_stage_inst_dmem_n18178) );
NAND2_X1 MEM_stage_inst_dmem_U16725 ( .A1(MEM_stage_inst_dmem_n18176), .A2(MEM_stage_inst_dmem_n18175), .ZN(MEM_stage_inst_dmem_n10297) );
NAND2_X1 MEM_stage_inst_dmem_U16724 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n18204), .ZN(MEM_stage_inst_dmem_n18175) );
NAND2_X1 MEM_stage_inst_dmem_U16723 ( .A1(MEM_stage_inst_dmem_ram_3070), .A2(MEM_stage_inst_dmem_n18203), .ZN(MEM_stage_inst_dmem_n18176) );
NAND2_X1 MEM_stage_inst_dmem_U16722 ( .A1(MEM_stage_inst_dmem_n18174), .A2(MEM_stage_inst_dmem_n18173), .ZN(MEM_stage_inst_dmem_n10298) );
NAND2_X1 MEM_stage_inst_dmem_U16721 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n18204), .ZN(MEM_stage_inst_dmem_n18173) );
INV_X1 MEM_stage_inst_dmem_U16720 ( .A(MEM_stage_inst_dmem_n18203), .ZN(MEM_stage_inst_dmem_n18204) );
NAND2_X1 MEM_stage_inst_dmem_U16719 ( .A1(MEM_stage_inst_dmem_ram_3071), .A2(MEM_stage_inst_dmem_n18203), .ZN(MEM_stage_inst_dmem_n18174) );
NAND2_X1 MEM_stage_inst_dmem_U16718 ( .A1(MEM_stage_inst_dmem_n20934), .A2(MEM_stage_inst_dmem_n18683), .ZN(MEM_stage_inst_dmem_n18203) );
NOR2_X2 MEM_stage_inst_dmem_U16717 ( .A1(MEM_stage_inst_dmem_n18718), .A2(MEM_stage_inst_dmem_n20369), .ZN(MEM_stage_inst_dmem_n18683) );
NAND2_X1 MEM_stage_inst_dmem_U16716 ( .A1(MEM_stage_inst_dmem_n18172), .A2(MEM_stage_inst_dmem_n18171), .ZN(MEM_stage_inst_dmem_n10299) );
NAND2_X1 MEM_stage_inst_dmem_U16715 ( .A1(MEM_stage_inst_dmem_n20551), .A2(MEM_stage_inst_dmem_n18170), .ZN(MEM_stage_inst_dmem_n18171) );
NAND2_X1 MEM_stage_inst_dmem_U16714 ( .A1(MEM_stage_inst_dmem_ram_2048), .A2(MEM_stage_inst_dmem_n18169), .ZN(MEM_stage_inst_dmem_n18172) );
NAND2_X1 MEM_stage_inst_dmem_U16713 ( .A1(MEM_stage_inst_dmem_n18168), .A2(MEM_stage_inst_dmem_n18167), .ZN(MEM_stage_inst_dmem_n10300) );
NAND2_X1 MEM_stage_inst_dmem_U16712 ( .A1(MEM_stage_inst_dmem_n20547), .A2(MEM_stage_inst_dmem_n18170), .ZN(MEM_stage_inst_dmem_n18167) );
NAND2_X1 MEM_stage_inst_dmem_U16711 ( .A1(MEM_stage_inst_dmem_ram_2049), .A2(MEM_stage_inst_dmem_n18169), .ZN(MEM_stage_inst_dmem_n18168) );
NAND2_X1 MEM_stage_inst_dmem_U16710 ( .A1(MEM_stage_inst_dmem_n18166), .A2(MEM_stage_inst_dmem_n18165), .ZN(MEM_stage_inst_dmem_n10301) );
NAND2_X1 MEM_stage_inst_dmem_U16709 ( .A1(MEM_stage_inst_dmem_n20544), .A2(MEM_stage_inst_dmem_n18170), .ZN(MEM_stage_inst_dmem_n18165) );
NAND2_X1 MEM_stage_inst_dmem_U16708 ( .A1(MEM_stage_inst_dmem_ram_2050), .A2(MEM_stage_inst_dmem_n18169), .ZN(MEM_stage_inst_dmem_n18166) );
NAND2_X1 MEM_stage_inst_dmem_U16707 ( .A1(MEM_stage_inst_dmem_n18164), .A2(MEM_stage_inst_dmem_n18163), .ZN(MEM_stage_inst_dmem_n10302) );
NAND2_X1 MEM_stage_inst_dmem_U16706 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n18170), .ZN(MEM_stage_inst_dmem_n18163) );
NAND2_X1 MEM_stage_inst_dmem_U16705 ( .A1(MEM_stage_inst_dmem_ram_2051), .A2(MEM_stage_inst_dmem_n18169), .ZN(MEM_stage_inst_dmem_n18164) );
NAND2_X1 MEM_stage_inst_dmem_U16704 ( .A1(MEM_stage_inst_dmem_n18162), .A2(MEM_stage_inst_dmem_n18161), .ZN(MEM_stage_inst_dmem_n10303) );
NAND2_X1 MEM_stage_inst_dmem_U16703 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n18170), .ZN(MEM_stage_inst_dmem_n18161) );
NAND2_X1 MEM_stage_inst_dmem_U16702 ( .A1(MEM_stage_inst_dmem_ram_2052), .A2(MEM_stage_inst_dmem_n18169), .ZN(MEM_stage_inst_dmem_n18162) );
NAND2_X1 MEM_stage_inst_dmem_U16701 ( .A1(MEM_stage_inst_dmem_n18160), .A2(MEM_stage_inst_dmem_n18159), .ZN(MEM_stage_inst_dmem_n10304) );
NAND2_X1 MEM_stage_inst_dmem_U16700 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n18170), .ZN(MEM_stage_inst_dmem_n18159) );
NAND2_X1 MEM_stage_inst_dmem_U16699 ( .A1(MEM_stage_inst_dmem_ram_2053), .A2(MEM_stage_inst_dmem_n18169), .ZN(MEM_stage_inst_dmem_n18160) );
NAND2_X1 MEM_stage_inst_dmem_U16698 ( .A1(MEM_stage_inst_dmem_n18158), .A2(MEM_stage_inst_dmem_n18157), .ZN(MEM_stage_inst_dmem_n10305) );
NAND2_X1 MEM_stage_inst_dmem_U16697 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n18170), .ZN(MEM_stage_inst_dmem_n18157) );
NAND2_X1 MEM_stage_inst_dmem_U16696 ( .A1(MEM_stage_inst_dmem_ram_2054), .A2(MEM_stage_inst_dmem_n18169), .ZN(MEM_stage_inst_dmem_n18158) );
NAND2_X1 MEM_stage_inst_dmem_U16695 ( .A1(MEM_stage_inst_dmem_n18156), .A2(MEM_stage_inst_dmem_n18155), .ZN(MEM_stage_inst_dmem_n10306) );
NAND2_X1 MEM_stage_inst_dmem_U16694 ( .A1(MEM_stage_inst_dmem_n20530), .A2(MEM_stage_inst_dmem_n18170), .ZN(MEM_stage_inst_dmem_n18155) );
NAND2_X1 MEM_stage_inst_dmem_U16693 ( .A1(MEM_stage_inst_dmem_ram_2055), .A2(MEM_stage_inst_dmem_n18169), .ZN(MEM_stage_inst_dmem_n18156) );
NAND2_X1 MEM_stage_inst_dmem_U16692 ( .A1(MEM_stage_inst_dmem_n18154), .A2(MEM_stage_inst_dmem_n18153), .ZN(MEM_stage_inst_dmem_n10307) );
NAND2_X1 MEM_stage_inst_dmem_U16691 ( .A1(MEM_stage_inst_dmem_n20527), .A2(MEM_stage_inst_dmem_n18170), .ZN(MEM_stage_inst_dmem_n18153) );
NAND2_X1 MEM_stage_inst_dmem_U16690 ( .A1(MEM_stage_inst_dmem_ram_2056), .A2(MEM_stage_inst_dmem_n18169), .ZN(MEM_stage_inst_dmem_n18154) );
NAND2_X1 MEM_stage_inst_dmem_U16689 ( .A1(MEM_stage_inst_dmem_n18152), .A2(MEM_stage_inst_dmem_n18151), .ZN(MEM_stage_inst_dmem_n10308) );
NAND2_X1 MEM_stage_inst_dmem_U16688 ( .A1(MEM_stage_inst_dmem_n20524), .A2(MEM_stage_inst_dmem_n18170), .ZN(MEM_stage_inst_dmem_n18151) );
NAND2_X1 MEM_stage_inst_dmem_U16687 ( .A1(MEM_stage_inst_dmem_ram_2057), .A2(MEM_stage_inst_dmem_n18169), .ZN(MEM_stage_inst_dmem_n18152) );
NAND2_X1 MEM_stage_inst_dmem_U16686 ( .A1(MEM_stage_inst_dmem_n18150), .A2(MEM_stage_inst_dmem_n18149), .ZN(MEM_stage_inst_dmem_n10309) );
NAND2_X1 MEM_stage_inst_dmem_U16685 ( .A1(MEM_stage_inst_dmem_n20521), .A2(MEM_stage_inst_dmem_n18170), .ZN(MEM_stage_inst_dmem_n18149) );
NAND2_X1 MEM_stage_inst_dmem_U16684 ( .A1(MEM_stage_inst_dmem_ram_2058), .A2(MEM_stage_inst_dmem_n18169), .ZN(MEM_stage_inst_dmem_n18150) );
NAND2_X1 MEM_stage_inst_dmem_U16683 ( .A1(MEM_stage_inst_dmem_n18148), .A2(MEM_stage_inst_dmem_n18147), .ZN(MEM_stage_inst_dmem_n10310) );
NAND2_X1 MEM_stage_inst_dmem_U16682 ( .A1(MEM_stage_inst_dmem_n20518), .A2(MEM_stage_inst_dmem_n18170), .ZN(MEM_stage_inst_dmem_n18147) );
NAND2_X1 MEM_stage_inst_dmem_U16681 ( .A1(MEM_stage_inst_dmem_ram_2059), .A2(MEM_stage_inst_dmem_n18169), .ZN(MEM_stage_inst_dmem_n18148) );
NAND2_X1 MEM_stage_inst_dmem_U16680 ( .A1(MEM_stage_inst_dmem_n18146), .A2(MEM_stage_inst_dmem_n18145), .ZN(MEM_stage_inst_dmem_n10311) );
NAND2_X1 MEM_stage_inst_dmem_U16679 ( .A1(MEM_stage_inst_dmem_n20515), .A2(MEM_stage_inst_dmem_n18170), .ZN(MEM_stage_inst_dmem_n18145) );
NAND2_X1 MEM_stage_inst_dmem_U16678 ( .A1(MEM_stage_inst_dmem_ram_2060), .A2(MEM_stage_inst_dmem_n18169), .ZN(MEM_stage_inst_dmem_n18146) );
NAND2_X1 MEM_stage_inst_dmem_U16677 ( .A1(MEM_stage_inst_dmem_n18144), .A2(MEM_stage_inst_dmem_n18143), .ZN(MEM_stage_inst_dmem_n10312) );
NAND2_X1 MEM_stage_inst_dmem_U16676 ( .A1(MEM_stage_inst_dmem_n20512), .A2(MEM_stage_inst_dmem_n18170), .ZN(MEM_stage_inst_dmem_n18143) );
NAND2_X1 MEM_stage_inst_dmem_U16675 ( .A1(MEM_stage_inst_dmem_ram_2061), .A2(MEM_stage_inst_dmem_n18169), .ZN(MEM_stage_inst_dmem_n18144) );
NAND2_X1 MEM_stage_inst_dmem_U16674 ( .A1(MEM_stage_inst_dmem_n18142), .A2(MEM_stage_inst_dmem_n18141), .ZN(MEM_stage_inst_dmem_n10313) );
NAND2_X1 MEM_stage_inst_dmem_U16673 ( .A1(MEM_stage_inst_dmem_n20509), .A2(MEM_stage_inst_dmem_n18170), .ZN(MEM_stage_inst_dmem_n18141) );
NAND2_X1 MEM_stage_inst_dmem_U16672 ( .A1(MEM_stage_inst_dmem_ram_2062), .A2(MEM_stage_inst_dmem_n18169), .ZN(MEM_stage_inst_dmem_n18142) );
NAND2_X1 MEM_stage_inst_dmem_U16671 ( .A1(MEM_stage_inst_dmem_n18140), .A2(MEM_stage_inst_dmem_n18139), .ZN(MEM_stage_inst_dmem_n10314) );
NAND2_X1 MEM_stage_inst_dmem_U16670 ( .A1(MEM_stage_inst_dmem_n20506), .A2(MEM_stage_inst_dmem_n18170), .ZN(MEM_stage_inst_dmem_n18139) );
INV_X1 MEM_stage_inst_dmem_U16669 ( .A(MEM_stage_inst_dmem_n18169), .ZN(MEM_stage_inst_dmem_n18170) );
NAND2_X1 MEM_stage_inst_dmem_U16668 ( .A1(MEM_stage_inst_dmem_ram_2063), .A2(MEM_stage_inst_dmem_n18169), .ZN(MEM_stage_inst_dmem_n18140) );
NAND2_X1 MEM_stage_inst_dmem_U16667 ( .A1(MEM_stage_inst_dmem_n21465), .A2(MEM_stage_inst_dmem_n18138), .ZN(MEM_stage_inst_dmem_n18169) );
NAND2_X1 MEM_stage_inst_dmem_U16666 ( .A1(MEM_stage_inst_dmem_n18137), .A2(MEM_stage_inst_dmem_n18136), .ZN(MEM_stage_inst_dmem_n10315) );
NAND2_X1 MEM_stage_inst_dmem_U16665 ( .A1(MEM_stage_inst_dmem_n19275), .A2(MEM_stage_inst_dmem_n18135), .ZN(MEM_stage_inst_dmem_n18136) );
NAND2_X1 MEM_stage_inst_dmem_U16664 ( .A1(MEM_stage_inst_dmem_ram_2064), .A2(MEM_stage_inst_dmem_n18134), .ZN(MEM_stage_inst_dmem_n18137) );
NAND2_X1 MEM_stage_inst_dmem_U16663 ( .A1(MEM_stage_inst_dmem_n18133), .A2(MEM_stage_inst_dmem_n18132), .ZN(MEM_stage_inst_dmem_n10316) );
NAND2_X1 MEM_stage_inst_dmem_U16662 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n18135), .ZN(MEM_stage_inst_dmem_n18132) );
NAND2_X1 MEM_stage_inst_dmem_U16661 ( .A1(MEM_stage_inst_dmem_ram_2065), .A2(MEM_stage_inst_dmem_n18134), .ZN(MEM_stage_inst_dmem_n18133) );
NAND2_X1 MEM_stage_inst_dmem_U16660 ( .A1(MEM_stage_inst_dmem_n18131), .A2(MEM_stage_inst_dmem_n18130), .ZN(MEM_stage_inst_dmem_n10317) );
NAND2_X1 MEM_stage_inst_dmem_U16659 ( .A1(MEM_stage_inst_dmem_n18027), .A2(MEM_stage_inst_dmem_n18135), .ZN(MEM_stage_inst_dmem_n18130) );
NAND2_X1 MEM_stage_inst_dmem_U16658 ( .A1(MEM_stage_inst_dmem_ram_2066), .A2(MEM_stage_inst_dmem_n18134), .ZN(MEM_stage_inst_dmem_n18131) );
NAND2_X1 MEM_stage_inst_dmem_U16657 ( .A1(MEM_stage_inst_dmem_n18129), .A2(MEM_stage_inst_dmem_n18128), .ZN(MEM_stage_inst_dmem_n10318) );
NAND2_X1 MEM_stage_inst_dmem_U16656 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n18135), .ZN(MEM_stage_inst_dmem_n18128) );
NAND2_X1 MEM_stage_inst_dmem_U16655 ( .A1(MEM_stage_inst_dmem_ram_2067), .A2(MEM_stage_inst_dmem_n18134), .ZN(MEM_stage_inst_dmem_n18129) );
NAND2_X1 MEM_stage_inst_dmem_U16654 ( .A1(MEM_stage_inst_dmem_n18127), .A2(MEM_stage_inst_dmem_n18126), .ZN(MEM_stage_inst_dmem_n10319) );
NAND2_X1 MEM_stage_inst_dmem_U16653 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n18135), .ZN(MEM_stage_inst_dmem_n18126) );
NAND2_X1 MEM_stage_inst_dmem_U16652 ( .A1(MEM_stage_inst_dmem_ram_2068), .A2(MEM_stage_inst_dmem_n18134), .ZN(MEM_stage_inst_dmem_n18127) );
NAND2_X1 MEM_stage_inst_dmem_U16651 ( .A1(MEM_stage_inst_dmem_n18125), .A2(MEM_stage_inst_dmem_n18124), .ZN(MEM_stage_inst_dmem_n10320) );
NAND2_X1 MEM_stage_inst_dmem_U16650 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n18135), .ZN(MEM_stage_inst_dmem_n18124) );
NAND2_X1 MEM_stage_inst_dmem_U16649 ( .A1(MEM_stage_inst_dmem_ram_2069), .A2(MEM_stage_inst_dmem_n18134), .ZN(MEM_stage_inst_dmem_n18125) );
NAND2_X1 MEM_stage_inst_dmem_U16648 ( .A1(MEM_stage_inst_dmem_n18123), .A2(MEM_stage_inst_dmem_n18122), .ZN(MEM_stage_inst_dmem_n10321) );
NAND2_X1 MEM_stage_inst_dmem_U16647 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n18135), .ZN(MEM_stage_inst_dmem_n18122) );
NAND2_X1 MEM_stage_inst_dmem_U16646 ( .A1(MEM_stage_inst_dmem_ram_2070), .A2(MEM_stage_inst_dmem_n18134), .ZN(MEM_stage_inst_dmem_n18123) );
NAND2_X1 MEM_stage_inst_dmem_U16645 ( .A1(MEM_stage_inst_dmem_n18121), .A2(MEM_stage_inst_dmem_n18120), .ZN(MEM_stage_inst_dmem_n10322) );
NAND2_X1 MEM_stage_inst_dmem_U16644 ( .A1(MEM_stage_inst_dmem_n20530), .A2(MEM_stage_inst_dmem_n18135), .ZN(MEM_stage_inst_dmem_n18120) );
NAND2_X1 MEM_stage_inst_dmem_U16643 ( .A1(MEM_stage_inst_dmem_ram_2071), .A2(MEM_stage_inst_dmem_n18134), .ZN(MEM_stage_inst_dmem_n18121) );
NAND2_X1 MEM_stage_inst_dmem_U16642 ( .A1(MEM_stage_inst_dmem_n18119), .A2(MEM_stage_inst_dmem_n18118), .ZN(MEM_stage_inst_dmem_n10323) );
NAND2_X1 MEM_stage_inst_dmem_U16641 ( .A1(MEM_stage_inst_dmem_n20527), .A2(MEM_stage_inst_dmem_n18135), .ZN(MEM_stage_inst_dmem_n18118) );
NAND2_X1 MEM_stage_inst_dmem_U16640 ( .A1(MEM_stage_inst_dmem_ram_2072), .A2(MEM_stage_inst_dmem_n18134), .ZN(MEM_stage_inst_dmem_n18119) );
NAND2_X1 MEM_stage_inst_dmem_U16639 ( .A1(MEM_stage_inst_dmem_n18117), .A2(MEM_stage_inst_dmem_n18116), .ZN(MEM_stage_inst_dmem_n10324) );
NAND2_X1 MEM_stage_inst_dmem_U16638 ( .A1(MEM_stage_inst_dmem_n19251), .A2(MEM_stage_inst_dmem_n18135), .ZN(MEM_stage_inst_dmem_n18116) );
NAND2_X1 MEM_stage_inst_dmem_U16637 ( .A1(MEM_stage_inst_dmem_ram_2073), .A2(MEM_stage_inst_dmem_n18134), .ZN(MEM_stage_inst_dmem_n18117) );
NAND2_X1 MEM_stage_inst_dmem_U16636 ( .A1(MEM_stage_inst_dmem_n18115), .A2(MEM_stage_inst_dmem_n18114), .ZN(MEM_stage_inst_dmem_n10325) );
NAND2_X1 MEM_stage_inst_dmem_U16635 ( .A1(MEM_stage_inst_dmem_n18007), .A2(MEM_stage_inst_dmem_n18135), .ZN(MEM_stage_inst_dmem_n18114) );
NAND2_X1 MEM_stage_inst_dmem_U16634 ( .A1(MEM_stage_inst_dmem_ram_2074), .A2(MEM_stage_inst_dmem_n18134), .ZN(MEM_stage_inst_dmem_n18115) );
NAND2_X1 MEM_stage_inst_dmem_U16633 ( .A1(MEM_stage_inst_dmem_n18113), .A2(MEM_stage_inst_dmem_n18112), .ZN(MEM_stage_inst_dmem_n10326) );
NAND2_X1 MEM_stage_inst_dmem_U16632 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n18135), .ZN(MEM_stage_inst_dmem_n18112) );
NAND2_X1 MEM_stage_inst_dmem_U16631 ( .A1(MEM_stage_inst_dmem_ram_2075), .A2(MEM_stage_inst_dmem_n18134), .ZN(MEM_stage_inst_dmem_n18113) );
NAND2_X1 MEM_stage_inst_dmem_U16630 ( .A1(MEM_stage_inst_dmem_n18111), .A2(MEM_stage_inst_dmem_n18110), .ZN(MEM_stage_inst_dmem_n10327) );
NAND2_X1 MEM_stage_inst_dmem_U16629 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n18135), .ZN(MEM_stage_inst_dmem_n18110) );
NAND2_X1 MEM_stage_inst_dmem_U16628 ( .A1(MEM_stage_inst_dmem_ram_2076), .A2(MEM_stage_inst_dmem_n18134), .ZN(MEM_stage_inst_dmem_n18111) );
NAND2_X1 MEM_stage_inst_dmem_U16627 ( .A1(MEM_stage_inst_dmem_n18109), .A2(MEM_stage_inst_dmem_n18108), .ZN(MEM_stage_inst_dmem_n10328) );
NAND2_X1 MEM_stage_inst_dmem_U16626 ( .A1(MEM_stage_inst_dmem_n19242), .A2(MEM_stage_inst_dmem_n18135), .ZN(MEM_stage_inst_dmem_n18108) );
NAND2_X1 MEM_stage_inst_dmem_U16625 ( .A1(MEM_stage_inst_dmem_ram_2077), .A2(MEM_stage_inst_dmem_n18134), .ZN(MEM_stage_inst_dmem_n18109) );
NAND2_X1 MEM_stage_inst_dmem_U16624 ( .A1(MEM_stage_inst_dmem_n18107), .A2(MEM_stage_inst_dmem_n18106), .ZN(MEM_stage_inst_dmem_n10329) );
NAND2_X1 MEM_stage_inst_dmem_U16623 ( .A1(MEM_stage_inst_dmem_n115), .A2(MEM_stage_inst_dmem_n18135), .ZN(MEM_stage_inst_dmem_n18106) );
NAND2_X1 MEM_stage_inst_dmem_U16622 ( .A1(MEM_stage_inst_dmem_ram_2078), .A2(MEM_stage_inst_dmem_n18134), .ZN(MEM_stage_inst_dmem_n18107) );
NAND2_X1 MEM_stage_inst_dmem_U16621 ( .A1(MEM_stage_inst_dmem_n18105), .A2(MEM_stage_inst_dmem_n18104), .ZN(MEM_stage_inst_dmem_n10330) );
NAND2_X1 MEM_stage_inst_dmem_U16620 ( .A1(MEM_stage_inst_dmem_n20506), .A2(MEM_stage_inst_dmem_n18135), .ZN(MEM_stage_inst_dmem_n18104) );
INV_X1 MEM_stage_inst_dmem_U16619 ( .A(MEM_stage_inst_dmem_n18134), .ZN(MEM_stage_inst_dmem_n18135) );
NAND2_X1 MEM_stage_inst_dmem_U16618 ( .A1(MEM_stage_inst_dmem_ram_2079), .A2(MEM_stage_inst_dmem_n18134), .ZN(MEM_stage_inst_dmem_n18105) );
NAND2_X1 MEM_stage_inst_dmem_U16617 ( .A1(MEM_stage_inst_dmem_n21429), .A2(MEM_stage_inst_dmem_n18138), .ZN(MEM_stage_inst_dmem_n18134) );
NAND2_X1 MEM_stage_inst_dmem_U16616 ( .A1(MEM_stage_inst_dmem_n18103), .A2(MEM_stage_inst_dmem_n18102), .ZN(MEM_stage_inst_dmem_n10331) );
NAND2_X1 MEM_stage_inst_dmem_U16615 ( .A1(MEM_stage_inst_dmem_n15145), .A2(MEM_stage_inst_dmem_n18101), .ZN(MEM_stage_inst_dmem_n18102) );
NAND2_X1 MEM_stage_inst_dmem_U16614 ( .A1(MEM_stage_inst_dmem_ram_2080), .A2(MEM_stage_inst_dmem_n18100), .ZN(MEM_stage_inst_dmem_n18103) );
NAND2_X1 MEM_stage_inst_dmem_U16613 ( .A1(MEM_stage_inst_dmem_n18099), .A2(MEM_stage_inst_dmem_n18098), .ZN(MEM_stage_inst_dmem_n10332) );
NAND2_X1 MEM_stage_inst_dmem_U16612 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n18101), .ZN(MEM_stage_inst_dmem_n18098) );
NAND2_X1 MEM_stage_inst_dmem_U16611 ( .A1(MEM_stage_inst_dmem_ram_2081), .A2(MEM_stage_inst_dmem_n18100), .ZN(MEM_stage_inst_dmem_n18099) );
NAND2_X1 MEM_stage_inst_dmem_U16610 ( .A1(MEM_stage_inst_dmem_n18097), .A2(MEM_stage_inst_dmem_n18096), .ZN(MEM_stage_inst_dmem_n10333) );
NAND2_X1 MEM_stage_inst_dmem_U16609 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n18101), .ZN(MEM_stage_inst_dmem_n18096) );
NAND2_X1 MEM_stage_inst_dmem_U16608 ( .A1(MEM_stage_inst_dmem_ram_2082), .A2(MEM_stage_inst_dmem_n18100), .ZN(MEM_stage_inst_dmem_n18097) );
NAND2_X1 MEM_stage_inst_dmem_U16607 ( .A1(MEM_stage_inst_dmem_n18095), .A2(MEM_stage_inst_dmem_n18094), .ZN(MEM_stage_inst_dmem_n10334) );
NAND2_X1 MEM_stage_inst_dmem_U16606 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n18101), .ZN(MEM_stage_inst_dmem_n18094) );
NAND2_X1 MEM_stage_inst_dmem_U16605 ( .A1(MEM_stage_inst_dmem_ram_2083), .A2(MEM_stage_inst_dmem_n18100), .ZN(MEM_stage_inst_dmem_n18095) );
NAND2_X1 MEM_stage_inst_dmem_U16604 ( .A1(MEM_stage_inst_dmem_n18093), .A2(MEM_stage_inst_dmem_n18092), .ZN(MEM_stage_inst_dmem_n10335) );
NAND2_X1 MEM_stage_inst_dmem_U16603 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n18101), .ZN(MEM_stage_inst_dmem_n18092) );
NAND2_X1 MEM_stage_inst_dmem_U16602 ( .A1(MEM_stage_inst_dmem_ram_2084), .A2(MEM_stage_inst_dmem_n18100), .ZN(MEM_stage_inst_dmem_n18093) );
NAND2_X1 MEM_stage_inst_dmem_U16601 ( .A1(MEM_stage_inst_dmem_n18091), .A2(MEM_stage_inst_dmem_n18090), .ZN(MEM_stage_inst_dmem_n10336) );
NAND2_X1 MEM_stage_inst_dmem_U16600 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n18101), .ZN(MEM_stage_inst_dmem_n18090) );
NAND2_X1 MEM_stage_inst_dmem_U16599 ( .A1(MEM_stage_inst_dmem_ram_2085), .A2(MEM_stage_inst_dmem_n18100), .ZN(MEM_stage_inst_dmem_n18091) );
NAND2_X1 MEM_stage_inst_dmem_U16598 ( .A1(MEM_stage_inst_dmem_n18089), .A2(MEM_stage_inst_dmem_n18088), .ZN(MEM_stage_inst_dmem_n10337) );
NAND2_X1 MEM_stage_inst_dmem_U16597 ( .A1(MEM_stage_inst_dmem_n21340), .A2(MEM_stage_inst_dmem_n18101), .ZN(MEM_stage_inst_dmem_n18088) );
NAND2_X1 MEM_stage_inst_dmem_U16596 ( .A1(MEM_stage_inst_dmem_ram_2086), .A2(MEM_stage_inst_dmem_n18100), .ZN(MEM_stage_inst_dmem_n18089) );
NAND2_X1 MEM_stage_inst_dmem_U16595 ( .A1(MEM_stage_inst_dmem_n18087), .A2(MEM_stage_inst_dmem_n18086), .ZN(MEM_stage_inst_dmem_n10338) );
NAND2_X1 MEM_stage_inst_dmem_U16594 ( .A1(MEM_stage_inst_dmem_n18), .A2(MEM_stage_inst_dmem_n18101), .ZN(MEM_stage_inst_dmem_n18086) );
NAND2_X1 MEM_stage_inst_dmem_U16593 ( .A1(MEM_stage_inst_dmem_ram_2087), .A2(MEM_stage_inst_dmem_n18100), .ZN(MEM_stage_inst_dmem_n18087) );
NAND2_X1 MEM_stage_inst_dmem_U16592 ( .A1(MEM_stage_inst_dmem_n18085), .A2(MEM_stage_inst_dmem_n18084), .ZN(MEM_stage_inst_dmem_n10339) );
NAND2_X1 MEM_stage_inst_dmem_U16591 ( .A1(MEM_stage_inst_dmem_n21335), .A2(MEM_stage_inst_dmem_n18101), .ZN(MEM_stage_inst_dmem_n18084) );
BUF_X1 MEM_stage_inst_dmem_U16590 ( .A(MEM_stage_inst_dmem_n104), .Z(MEM_stage_inst_dmem_n21335) );
NAND2_X1 MEM_stage_inst_dmem_U16589 ( .A1(MEM_stage_inst_dmem_ram_2088), .A2(MEM_stage_inst_dmem_n18100), .ZN(MEM_stage_inst_dmem_n18085) );
NAND2_X1 MEM_stage_inst_dmem_U16588 ( .A1(MEM_stage_inst_dmem_n18083), .A2(MEM_stage_inst_dmem_n18082), .ZN(MEM_stage_inst_dmem_n10340) );
NAND2_X1 MEM_stage_inst_dmem_U16587 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n18101), .ZN(MEM_stage_inst_dmem_n18082) );
NAND2_X1 MEM_stage_inst_dmem_U16586 ( .A1(MEM_stage_inst_dmem_ram_2089), .A2(MEM_stage_inst_dmem_n18100), .ZN(MEM_stage_inst_dmem_n18083) );
NAND2_X1 MEM_stage_inst_dmem_U16585 ( .A1(MEM_stage_inst_dmem_n18081), .A2(MEM_stage_inst_dmem_n18080), .ZN(MEM_stage_inst_dmem_n10341) );
NAND2_X1 MEM_stage_inst_dmem_U16584 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n18101), .ZN(MEM_stage_inst_dmem_n18080) );
NAND2_X1 MEM_stage_inst_dmem_U16583 ( .A1(MEM_stage_inst_dmem_ram_2090), .A2(MEM_stage_inst_dmem_n18100), .ZN(MEM_stage_inst_dmem_n18081) );
NAND2_X1 MEM_stage_inst_dmem_U16582 ( .A1(MEM_stage_inst_dmem_n18079), .A2(MEM_stage_inst_dmem_n18078), .ZN(MEM_stage_inst_dmem_n10342) );
NAND2_X1 MEM_stage_inst_dmem_U16581 ( .A1(MEM_stage_inst_dmem_n20904), .A2(MEM_stage_inst_dmem_n18101), .ZN(MEM_stage_inst_dmem_n18078) );
NAND2_X1 MEM_stage_inst_dmem_U16580 ( .A1(MEM_stage_inst_dmem_ram_2091), .A2(MEM_stage_inst_dmem_n18100), .ZN(MEM_stage_inst_dmem_n18079) );
NAND2_X1 MEM_stage_inst_dmem_U16579 ( .A1(MEM_stage_inst_dmem_n18077), .A2(MEM_stage_inst_dmem_n18076), .ZN(MEM_stage_inst_dmem_n10343) );
NAND2_X1 MEM_stage_inst_dmem_U16578 ( .A1(MEM_stage_inst_dmem_n21474), .A2(MEM_stage_inst_dmem_n18101), .ZN(MEM_stage_inst_dmem_n18076) );
NAND2_X1 MEM_stage_inst_dmem_U16577 ( .A1(MEM_stage_inst_dmem_ram_2092), .A2(MEM_stage_inst_dmem_n18100), .ZN(MEM_stage_inst_dmem_n18077) );
NAND2_X1 MEM_stage_inst_dmem_U16576 ( .A1(MEM_stage_inst_dmem_n18075), .A2(MEM_stage_inst_dmem_n18074), .ZN(MEM_stage_inst_dmem_n10344) );
NAND2_X1 MEM_stage_inst_dmem_U16575 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n18101), .ZN(MEM_stage_inst_dmem_n18074) );
NAND2_X1 MEM_stage_inst_dmem_U16574 ( .A1(MEM_stage_inst_dmem_ram_2093), .A2(MEM_stage_inst_dmem_n18100), .ZN(MEM_stage_inst_dmem_n18075) );
NAND2_X1 MEM_stage_inst_dmem_U16573 ( .A1(MEM_stage_inst_dmem_n18073), .A2(MEM_stage_inst_dmem_n18072), .ZN(MEM_stage_inst_dmem_n10345) );
NAND2_X1 MEM_stage_inst_dmem_U16572 ( .A1(MEM_stage_inst_dmem_n15113), .A2(MEM_stage_inst_dmem_n18101), .ZN(MEM_stage_inst_dmem_n18072) );
NAND2_X1 MEM_stage_inst_dmem_U16571 ( .A1(MEM_stage_inst_dmem_ram_2094), .A2(MEM_stage_inst_dmem_n18100), .ZN(MEM_stage_inst_dmem_n18073) );
NAND2_X1 MEM_stage_inst_dmem_U16570 ( .A1(MEM_stage_inst_dmem_n18071), .A2(MEM_stage_inst_dmem_n18070), .ZN(MEM_stage_inst_dmem_n10346) );
NAND2_X1 MEM_stage_inst_dmem_U16569 ( .A1(MEM_stage_inst_dmem_n21320), .A2(MEM_stage_inst_dmem_n18101), .ZN(MEM_stage_inst_dmem_n18070) );
INV_X1 MEM_stage_inst_dmem_U16568 ( .A(MEM_stage_inst_dmem_n18100), .ZN(MEM_stage_inst_dmem_n18101) );
NAND2_X1 MEM_stage_inst_dmem_U16567 ( .A1(MEM_stage_inst_dmem_ram_2095), .A2(MEM_stage_inst_dmem_n18100), .ZN(MEM_stage_inst_dmem_n18071) );
NAND2_X1 MEM_stage_inst_dmem_U16566 ( .A1(MEM_stage_inst_dmem_n21394), .A2(MEM_stage_inst_dmem_n18138), .ZN(MEM_stage_inst_dmem_n18100) );
NAND2_X1 MEM_stage_inst_dmem_U16565 ( .A1(MEM_stage_inst_dmem_n18069), .A2(MEM_stage_inst_dmem_n18068), .ZN(MEM_stage_inst_dmem_n10347) );
NAND2_X1 MEM_stage_inst_dmem_U16564 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n18067), .ZN(MEM_stage_inst_dmem_n18068) );
NAND2_X1 MEM_stage_inst_dmem_U16563 ( .A1(MEM_stage_inst_dmem_ram_2096), .A2(MEM_stage_inst_dmem_n18066), .ZN(MEM_stage_inst_dmem_n18069) );
NAND2_X1 MEM_stage_inst_dmem_U16562 ( .A1(MEM_stage_inst_dmem_n18065), .A2(MEM_stage_inst_dmem_n18064), .ZN(MEM_stage_inst_dmem_n10348) );
NAND2_X1 MEM_stage_inst_dmem_U16561 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n18067), .ZN(MEM_stage_inst_dmem_n18064) );
NAND2_X1 MEM_stage_inst_dmem_U16560 ( .A1(MEM_stage_inst_dmem_ram_2097), .A2(MEM_stage_inst_dmem_n18066), .ZN(MEM_stage_inst_dmem_n18065) );
NAND2_X1 MEM_stage_inst_dmem_U16559 ( .A1(MEM_stage_inst_dmem_n18063), .A2(MEM_stage_inst_dmem_n18062), .ZN(MEM_stage_inst_dmem_n10349) );
NAND2_X1 MEM_stage_inst_dmem_U16558 ( .A1(MEM_stage_inst_dmem_n18887), .A2(MEM_stage_inst_dmem_n18067), .ZN(MEM_stage_inst_dmem_n18062) );
NAND2_X1 MEM_stage_inst_dmem_U16557 ( .A1(MEM_stage_inst_dmem_ram_2098), .A2(MEM_stage_inst_dmem_n18066), .ZN(MEM_stage_inst_dmem_n18063) );
NAND2_X1 MEM_stage_inst_dmem_U16556 ( .A1(MEM_stage_inst_dmem_n18061), .A2(MEM_stage_inst_dmem_n18060), .ZN(MEM_stage_inst_dmem_n10350) );
NAND2_X1 MEM_stage_inst_dmem_U16555 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n18067), .ZN(MEM_stage_inst_dmem_n18060) );
NAND2_X1 MEM_stage_inst_dmem_U16554 ( .A1(MEM_stage_inst_dmem_ram_2099), .A2(MEM_stage_inst_dmem_n18066), .ZN(MEM_stage_inst_dmem_n18061) );
NAND2_X1 MEM_stage_inst_dmem_U16553 ( .A1(MEM_stage_inst_dmem_n18059), .A2(MEM_stage_inst_dmem_n18058), .ZN(MEM_stage_inst_dmem_n10351) );
NAND2_X1 MEM_stage_inst_dmem_U16552 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n18067), .ZN(MEM_stage_inst_dmem_n18058) );
NAND2_X1 MEM_stage_inst_dmem_U16551 ( .A1(MEM_stage_inst_dmem_ram_2100), .A2(MEM_stage_inst_dmem_n18066), .ZN(MEM_stage_inst_dmem_n18059) );
NAND2_X1 MEM_stage_inst_dmem_U16550 ( .A1(MEM_stage_inst_dmem_n18057), .A2(MEM_stage_inst_dmem_n18056), .ZN(MEM_stage_inst_dmem_n10352) );
NAND2_X1 MEM_stage_inst_dmem_U16549 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n18067), .ZN(MEM_stage_inst_dmem_n18056) );
NAND2_X1 MEM_stage_inst_dmem_U16548 ( .A1(MEM_stage_inst_dmem_ram_2101), .A2(MEM_stage_inst_dmem_n18066), .ZN(MEM_stage_inst_dmem_n18057) );
NAND2_X1 MEM_stage_inst_dmem_U16547 ( .A1(MEM_stage_inst_dmem_n18055), .A2(MEM_stage_inst_dmem_n18054), .ZN(MEM_stage_inst_dmem_n10353) );
NAND2_X1 MEM_stage_inst_dmem_U16546 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n18067), .ZN(MEM_stage_inst_dmem_n18054) );
NAND2_X1 MEM_stage_inst_dmem_U16545 ( .A1(MEM_stage_inst_dmem_ram_2102), .A2(MEM_stage_inst_dmem_n18066), .ZN(MEM_stage_inst_dmem_n18055) );
NAND2_X1 MEM_stage_inst_dmem_U16544 ( .A1(MEM_stage_inst_dmem_n18053), .A2(MEM_stage_inst_dmem_n18052), .ZN(MEM_stage_inst_dmem_n10354) );
NAND2_X1 MEM_stage_inst_dmem_U16543 ( .A1(MEM_stage_inst_dmem_n18875), .A2(MEM_stage_inst_dmem_n18067), .ZN(MEM_stage_inst_dmem_n18052) );
NAND2_X1 MEM_stage_inst_dmem_U16542 ( .A1(MEM_stage_inst_dmem_ram_2103), .A2(MEM_stage_inst_dmem_n18066), .ZN(MEM_stage_inst_dmem_n18053) );
NAND2_X1 MEM_stage_inst_dmem_U16541 ( .A1(MEM_stage_inst_dmem_n18051), .A2(MEM_stage_inst_dmem_n18050), .ZN(MEM_stage_inst_dmem_n10355) );
NAND2_X1 MEM_stage_inst_dmem_U16540 ( .A1(MEM_stage_inst_dmem_n111), .A2(MEM_stage_inst_dmem_n18067), .ZN(MEM_stage_inst_dmem_n18050) );
NAND2_X1 MEM_stage_inst_dmem_U16539 ( .A1(MEM_stage_inst_dmem_ram_2104), .A2(MEM_stage_inst_dmem_n18066), .ZN(MEM_stage_inst_dmem_n18051) );
NAND2_X1 MEM_stage_inst_dmem_U16538 ( .A1(MEM_stage_inst_dmem_n18049), .A2(MEM_stage_inst_dmem_n18048), .ZN(MEM_stage_inst_dmem_n10356) );
NAND2_X1 MEM_stage_inst_dmem_U16537 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n18067), .ZN(MEM_stage_inst_dmem_n18048) );
NAND2_X1 MEM_stage_inst_dmem_U16536 ( .A1(MEM_stage_inst_dmem_ram_2105), .A2(MEM_stage_inst_dmem_n18066), .ZN(MEM_stage_inst_dmem_n18049) );
NAND2_X1 MEM_stage_inst_dmem_U16535 ( .A1(MEM_stage_inst_dmem_n18047), .A2(MEM_stage_inst_dmem_n18046), .ZN(MEM_stage_inst_dmem_n10357) );
NAND2_X1 MEM_stage_inst_dmem_U16534 ( .A1(MEM_stage_inst_dmem_n18867), .A2(MEM_stage_inst_dmem_n18067), .ZN(MEM_stage_inst_dmem_n18046) );
NAND2_X1 MEM_stage_inst_dmem_U16533 ( .A1(MEM_stage_inst_dmem_ram_2106), .A2(MEM_stage_inst_dmem_n18066), .ZN(MEM_stage_inst_dmem_n18047) );
NAND2_X1 MEM_stage_inst_dmem_U16532 ( .A1(MEM_stage_inst_dmem_n18045), .A2(MEM_stage_inst_dmem_n18044), .ZN(MEM_stage_inst_dmem_n10358) );
NAND2_X1 MEM_stage_inst_dmem_U16531 ( .A1(MEM_stage_inst_dmem_n18864), .A2(MEM_stage_inst_dmem_n18067), .ZN(MEM_stage_inst_dmem_n18044) );
NAND2_X1 MEM_stage_inst_dmem_U16530 ( .A1(MEM_stage_inst_dmem_ram_2107), .A2(MEM_stage_inst_dmem_n18066), .ZN(MEM_stage_inst_dmem_n18045) );
NAND2_X1 MEM_stage_inst_dmem_U16529 ( .A1(MEM_stage_inst_dmem_n18043), .A2(MEM_stage_inst_dmem_n18042), .ZN(MEM_stage_inst_dmem_n10359) );
NAND2_X1 MEM_stage_inst_dmem_U16528 ( .A1(MEM_stage_inst_dmem_n18861), .A2(MEM_stage_inst_dmem_n18067), .ZN(MEM_stage_inst_dmem_n18042) );
NAND2_X1 MEM_stage_inst_dmem_U16527 ( .A1(MEM_stage_inst_dmem_ram_2108), .A2(MEM_stage_inst_dmem_n18066), .ZN(MEM_stage_inst_dmem_n18043) );
NAND2_X1 MEM_stage_inst_dmem_U16526 ( .A1(MEM_stage_inst_dmem_n18041), .A2(MEM_stage_inst_dmem_n18040), .ZN(MEM_stage_inst_dmem_n10360) );
NAND2_X1 MEM_stage_inst_dmem_U16525 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n18067), .ZN(MEM_stage_inst_dmem_n18040) );
NAND2_X1 MEM_stage_inst_dmem_U16524 ( .A1(MEM_stage_inst_dmem_ram_2109), .A2(MEM_stage_inst_dmem_n18066), .ZN(MEM_stage_inst_dmem_n18041) );
NAND2_X1 MEM_stage_inst_dmem_U16523 ( .A1(MEM_stage_inst_dmem_n18039), .A2(MEM_stage_inst_dmem_n18038), .ZN(MEM_stage_inst_dmem_n10361) );
NAND2_X1 MEM_stage_inst_dmem_U16522 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n18067), .ZN(MEM_stage_inst_dmem_n18038) );
NAND2_X1 MEM_stage_inst_dmem_U16521 ( .A1(MEM_stage_inst_dmem_ram_2110), .A2(MEM_stage_inst_dmem_n18066), .ZN(MEM_stage_inst_dmem_n18039) );
NAND2_X1 MEM_stage_inst_dmem_U16520 ( .A1(MEM_stage_inst_dmem_n18037), .A2(MEM_stage_inst_dmem_n18036), .ZN(MEM_stage_inst_dmem_n10362) );
NAND2_X1 MEM_stage_inst_dmem_U16519 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n18067), .ZN(MEM_stage_inst_dmem_n18036) );
INV_X1 MEM_stage_inst_dmem_U16518 ( .A(MEM_stage_inst_dmem_n18066), .ZN(MEM_stage_inst_dmem_n18067) );
NAND2_X1 MEM_stage_inst_dmem_U16517 ( .A1(MEM_stage_inst_dmem_ram_2111), .A2(MEM_stage_inst_dmem_n18066), .ZN(MEM_stage_inst_dmem_n18037) );
NAND2_X1 MEM_stage_inst_dmem_U16516 ( .A1(MEM_stage_inst_dmem_n21359), .A2(MEM_stage_inst_dmem_n18138), .ZN(MEM_stage_inst_dmem_n18066) );
NAND2_X1 MEM_stage_inst_dmem_U16515 ( .A1(MEM_stage_inst_dmem_n18035), .A2(MEM_stage_inst_dmem_n18034), .ZN(MEM_stage_inst_dmem_n10363) );
NAND2_X1 MEM_stage_inst_dmem_U16514 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n18033), .ZN(MEM_stage_inst_dmem_n18034) );
NAND2_X1 MEM_stage_inst_dmem_U16513 ( .A1(MEM_stage_inst_dmem_ram_2112), .A2(MEM_stage_inst_dmem_n18032), .ZN(MEM_stage_inst_dmem_n18035) );
NAND2_X1 MEM_stage_inst_dmem_U16512 ( .A1(MEM_stage_inst_dmem_n18031), .A2(MEM_stage_inst_dmem_n18030), .ZN(MEM_stage_inst_dmem_n10364) );
NAND2_X1 MEM_stage_inst_dmem_U16511 ( .A1(MEM_stage_inst_dmem_n20547), .A2(MEM_stage_inst_dmem_n18033), .ZN(MEM_stage_inst_dmem_n18030) );
NAND2_X1 MEM_stage_inst_dmem_U16510 ( .A1(MEM_stage_inst_dmem_ram_2113), .A2(MEM_stage_inst_dmem_n18032), .ZN(MEM_stage_inst_dmem_n18031) );
NAND2_X1 MEM_stage_inst_dmem_U16509 ( .A1(MEM_stage_inst_dmem_n18029), .A2(MEM_stage_inst_dmem_n18028), .ZN(MEM_stage_inst_dmem_n10365) );
NAND2_X1 MEM_stage_inst_dmem_U16508 ( .A1(MEM_stage_inst_dmem_n18027), .A2(MEM_stage_inst_dmem_n18033), .ZN(MEM_stage_inst_dmem_n18028) );
NAND2_X1 MEM_stage_inst_dmem_U16507 ( .A1(MEM_stage_inst_dmem_ram_2114), .A2(MEM_stage_inst_dmem_n18032), .ZN(MEM_stage_inst_dmem_n18029) );
NAND2_X1 MEM_stage_inst_dmem_U16506 ( .A1(MEM_stage_inst_dmem_n18026), .A2(MEM_stage_inst_dmem_n18025), .ZN(MEM_stage_inst_dmem_n10366) );
NAND2_X1 MEM_stage_inst_dmem_U16505 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n18033), .ZN(MEM_stage_inst_dmem_n18025) );
NAND2_X1 MEM_stage_inst_dmem_U16504 ( .A1(MEM_stage_inst_dmem_ram_2115), .A2(MEM_stage_inst_dmem_n18032), .ZN(MEM_stage_inst_dmem_n18026) );
NAND2_X1 MEM_stage_inst_dmem_U16503 ( .A1(MEM_stage_inst_dmem_n18024), .A2(MEM_stage_inst_dmem_n18023), .ZN(MEM_stage_inst_dmem_n10367) );
NAND2_X1 MEM_stage_inst_dmem_U16502 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n18033), .ZN(MEM_stage_inst_dmem_n18023) );
NAND2_X1 MEM_stage_inst_dmem_U16501 ( .A1(MEM_stage_inst_dmem_ram_2116), .A2(MEM_stage_inst_dmem_n18032), .ZN(MEM_stage_inst_dmem_n18024) );
NAND2_X1 MEM_stage_inst_dmem_U16500 ( .A1(MEM_stage_inst_dmem_n18021), .A2(MEM_stage_inst_dmem_n18020), .ZN(MEM_stage_inst_dmem_n10368) );
NAND2_X1 MEM_stage_inst_dmem_U16499 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n18033), .ZN(MEM_stage_inst_dmem_n18020) );
NAND2_X1 MEM_stage_inst_dmem_U16498 ( .A1(MEM_stage_inst_dmem_ram_2117), .A2(MEM_stage_inst_dmem_n18032), .ZN(MEM_stage_inst_dmem_n18021) );
NAND2_X1 MEM_stage_inst_dmem_U16497 ( .A1(MEM_stage_inst_dmem_n18019), .A2(MEM_stage_inst_dmem_n18018), .ZN(MEM_stage_inst_dmem_n10369) );
NAND2_X1 MEM_stage_inst_dmem_U16496 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n18033), .ZN(MEM_stage_inst_dmem_n18018) );
NAND2_X1 MEM_stage_inst_dmem_U16495 ( .A1(MEM_stage_inst_dmem_ram_2118), .A2(MEM_stage_inst_dmem_n18032), .ZN(MEM_stage_inst_dmem_n18019) );
NAND2_X1 MEM_stage_inst_dmem_U16494 ( .A1(MEM_stage_inst_dmem_n18017), .A2(MEM_stage_inst_dmem_n18016), .ZN(MEM_stage_inst_dmem_n10370) );
NAND2_X1 MEM_stage_inst_dmem_U16493 ( .A1(MEM_stage_inst_dmem_n18), .A2(MEM_stage_inst_dmem_n18033), .ZN(MEM_stage_inst_dmem_n18016) );
NAND2_X1 MEM_stage_inst_dmem_U16492 ( .A1(MEM_stage_inst_dmem_ram_2119), .A2(MEM_stage_inst_dmem_n18032), .ZN(MEM_stage_inst_dmem_n18017) );
NAND2_X1 MEM_stage_inst_dmem_U16491 ( .A1(MEM_stage_inst_dmem_n18015), .A2(MEM_stage_inst_dmem_n18014), .ZN(MEM_stage_inst_dmem_n10371) );
NAND2_X1 MEM_stage_inst_dmem_U16490 ( .A1(MEM_stage_inst_dmem_n18013), .A2(MEM_stage_inst_dmem_n18033), .ZN(MEM_stage_inst_dmem_n18014) );
NAND2_X1 MEM_stage_inst_dmem_U16489 ( .A1(MEM_stage_inst_dmem_ram_2120), .A2(MEM_stage_inst_dmem_n18032), .ZN(MEM_stage_inst_dmem_n18015) );
NAND2_X1 MEM_stage_inst_dmem_U16488 ( .A1(MEM_stage_inst_dmem_n18012), .A2(MEM_stage_inst_dmem_n18011), .ZN(MEM_stage_inst_dmem_n10372) );
NAND2_X1 MEM_stage_inst_dmem_U16487 ( .A1(MEM_stage_inst_dmem_n96), .A2(MEM_stage_inst_dmem_n18033), .ZN(MEM_stage_inst_dmem_n18011) );
NAND2_X1 MEM_stage_inst_dmem_U16486 ( .A1(MEM_stage_inst_dmem_ram_2121), .A2(MEM_stage_inst_dmem_n18032), .ZN(MEM_stage_inst_dmem_n18012) );
NAND2_X1 MEM_stage_inst_dmem_U16485 ( .A1(MEM_stage_inst_dmem_n18009), .A2(MEM_stage_inst_dmem_n18008), .ZN(MEM_stage_inst_dmem_n10373) );
NAND2_X1 MEM_stage_inst_dmem_U16484 ( .A1(MEM_stage_inst_dmem_n18007), .A2(MEM_stage_inst_dmem_n18033), .ZN(MEM_stage_inst_dmem_n18008) );
NAND2_X1 MEM_stage_inst_dmem_U16483 ( .A1(MEM_stage_inst_dmem_ram_2122), .A2(MEM_stage_inst_dmem_n18032), .ZN(MEM_stage_inst_dmem_n18009) );
NAND2_X1 MEM_stage_inst_dmem_U16482 ( .A1(MEM_stage_inst_dmem_n18006), .A2(MEM_stage_inst_dmem_n18005), .ZN(MEM_stage_inst_dmem_n10374) );
NAND2_X1 MEM_stage_inst_dmem_U16481 ( .A1(MEM_stage_inst_dmem_n18004), .A2(MEM_stage_inst_dmem_n18033), .ZN(MEM_stage_inst_dmem_n18005) );
NAND2_X1 MEM_stage_inst_dmem_U16480 ( .A1(MEM_stage_inst_dmem_ram_2123), .A2(MEM_stage_inst_dmem_n18032), .ZN(MEM_stage_inst_dmem_n18006) );
NAND2_X1 MEM_stage_inst_dmem_U16479 ( .A1(MEM_stage_inst_dmem_n18003), .A2(MEM_stage_inst_dmem_n18002), .ZN(MEM_stage_inst_dmem_n10375) );
NAND2_X1 MEM_stage_inst_dmem_U16478 ( .A1(MEM_stage_inst_dmem_n18001), .A2(MEM_stage_inst_dmem_n18033), .ZN(MEM_stage_inst_dmem_n18002) );
NAND2_X1 MEM_stage_inst_dmem_U16477 ( .A1(MEM_stage_inst_dmem_ram_2124), .A2(MEM_stage_inst_dmem_n18032), .ZN(MEM_stage_inst_dmem_n18003) );
NAND2_X1 MEM_stage_inst_dmem_U16476 ( .A1(MEM_stage_inst_dmem_n18000), .A2(MEM_stage_inst_dmem_n17999), .ZN(MEM_stage_inst_dmem_n10376) );
NAND2_X1 MEM_stage_inst_dmem_U16475 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n18033), .ZN(MEM_stage_inst_dmem_n17999) );
NAND2_X1 MEM_stage_inst_dmem_U16474 ( .A1(MEM_stage_inst_dmem_ram_2125), .A2(MEM_stage_inst_dmem_n18032), .ZN(MEM_stage_inst_dmem_n18000) );
NAND2_X1 MEM_stage_inst_dmem_U16473 ( .A1(MEM_stage_inst_dmem_n17998), .A2(MEM_stage_inst_dmem_n17997), .ZN(MEM_stage_inst_dmem_n10377) );
NAND2_X1 MEM_stage_inst_dmem_U16472 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n18033), .ZN(MEM_stage_inst_dmem_n17997) );
NAND2_X1 MEM_stage_inst_dmem_U16471 ( .A1(MEM_stage_inst_dmem_ram_2126), .A2(MEM_stage_inst_dmem_n18032), .ZN(MEM_stage_inst_dmem_n17998) );
NAND2_X1 MEM_stage_inst_dmem_U16470 ( .A1(MEM_stage_inst_dmem_n17996), .A2(MEM_stage_inst_dmem_n17995), .ZN(MEM_stage_inst_dmem_n10378) );
NAND2_X1 MEM_stage_inst_dmem_U16469 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n18033), .ZN(MEM_stage_inst_dmem_n17995) );
INV_X1 MEM_stage_inst_dmem_U16468 ( .A(MEM_stage_inst_dmem_n18032), .ZN(MEM_stage_inst_dmem_n18033) );
NAND2_X1 MEM_stage_inst_dmem_U16467 ( .A1(MEM_stage_inst_dmem_ram_2127), .A2(MEM_stage_inst_dmem_n18032), .ZN(MEM_stage_inst_dmem_n17996) );
NAND2_X1 MEM_stage_inst_dmem_U16466 ( .A1(MEM_stage_inst_dmem_n21319), .A2(MEM_stage_inst_dmem_n18138), .ZN(MEM_stage_inst_dmem_n18032) );
NAND2_X1 MEM_stage_inst_dmem_U16465 ( .A1(MEM_stage_inst_dmem_n17993), .A2(MEM_stage_inst_dmem_n17992), .ZN(MEM_stage_inst_dmem_n10379) );
NAND2_X1 MEM_stage_inst_dmem_U16464 ( .A1(EX_pipeline_reg_out_5), .A2(MEM_stage_inst_dmem_n17991), .ZN(MEM_stage_inst_dmem_n17992) );
NAND2_X1 MEM_stage_inst_dmem_U16463 ( .A1(MEM_stage_inst_dmem_ram_2128), .A2(MEM_stage_inst_dmem_n17990), .ZN(MEM_stage_inst_dmem_n17993) );
NAND2_X1 MEM_stage_inst_dmem_U16462 ( .A1(MEM_stage_inst_dmem_n17989), .A2(MEM_stage_inst_dmem_n17988), .ZN(MEM_stage_inst_dmem_n10380) );
NAND2_X1 MEM_stage_inst_dmem_U16461 ( .A1(EX_pipeline_reg_out_6), .A2(MEM_stage_inst_dmem_n17991), .ZN(MEM_stage_inst_dmem_n17988) );
NAND2_X1 MEM_stage_inst_dmem_U16460 ( .A1(MEM_stage_inst_dmem_ram_2129), .A2(MEM_stage_inst_dmem_n17990), .ZN(MEM_stage_inst_dmem_n17989) );
NAND2_X1 MEM_stage_inst_dmem_U16459 ( .A1(MEM_stage_inst_dmem_n17987), .A2(MEM_stage_inst_dmem_n17986), .ZN(MEM_stage_inst_dmem_n10381) );
NAND2_X1 MEM_stage_inst_dmem_U16458 ( .A1(EX_pipeline_reg_out_7), .A2(MEM_stage_inst_dmem_n17991), .ZN(MEM_stage_inst_dmem_n17986) );
NAND2_X1 MEM_stage_inst_dmem_U16457 ( .A1(MEM_stage_inst_dmem_ram_2130), .A2(MEM_stage_inst_dmem_n17990), .ZN(MEM_stage_inst_dmem_n17987) );
NAND2_X1 MEM_stage_inst_dmem_U16456 ( .A1(MEM_stage_inst_dmem_n17985), .A2(MEM_stage_inst_dmem_n17984), .ZN(MEM_stage_inst_dmem_n10382) );
NAND2_X1 MEM_stage_inst_dmem_U16455 ( .A1(EX_pipeline_reg_out_8), .A2(MEM_stage_inst_dmem_n17991), .ZN(MEM_stage_inst_dmem_n17984) );
NAND2_X1 MEM_stage_inst_dmem_U16454 ( .A1(MEM_stage_inst_dmem_ram_2131), .A2(MEM_stage_inst_dmem_n17990), .ZN(MEM_stage_inst_dmem_n17985) );
NAND2_X1 MEM_stage_inst_dmem_U16453 ( .A1(MEM_stage_inst_dmem_n17983), .A2(MEM_stage_inst_dmem_n17982), .ZN(MEM_stage_inst_dmem_n10383) );
NAND2_X1 MEM_stage_inst_dmem_U16452 ( .A1(EX_pipeline_reg_out_9), .A2(MEM_stage_inst_dmem_n17991), .ZN(MEM_stage_inst_dmem_n17982) );
NAND2_X1 MEM_stage_inst_dmem_U16451 ( .A1(MEM_stage_inst_dmem_ram_2132), .A2(MEM_stage_inst_dmem_n17990), .ZN(MEM_stage_inst_dmem_n17983) );
NAND2_X1 MEM_stage_inst_dmem_U16450 ( .A1(MEM_stage_inst_dmem_n17981), .A2(MEM_stage_inst_dmem_n17980), .ZN(MEM_stage_inst_dmem_n10384) );
NAND2_X1 MEM_stage_inst_dmem_U16449 ( .A1(EX_pipeline_reg_out_10), .A2(MEM_stage_inst_dmem_n17991), .ZN(MEM_stage_inst_dmem_n17980) );
NAND2_X1 MEM_stage_inst_dmem_U16448 ( .A1(MEM_stage_inst_dmem_ram_2133), .A2(MEM_stage_inst_dmem_n17990), .ZN(MEM_stage_inst_dmem_n17981) );
NAND2_X1 MEM_stage_inst_dmem_U16447 ( .A1(MEM_stage_inst_dmem_n17979), .A2(MEM_stage_inst_dmem_n17978), .ZN(MEM_stage_inst_dmem_n10385) );
NAND2_X1 MEM_stage_inst_dmem_U16446 ( .A1(EX_pipeline_reg_out_11), .A2(MEM_stage_inst_dmem_n17991), .ZN(MEM_stage_inst_dmem_n17978) );
NAND2_X1 MEM_stage_inst_dmem_U16445 ( .A1(MEM_stage_inst_dmem_ram_2134), .A2(MEM_stage_inst_dmem_n17990), .ZN(MEM_stage_inst_dmem_n17979) );
NAND2_X1 MEM_stage_inst_dmem_U16444 ( .A1(MEM_stage_inst_dmem_n17977), .A2(MEM_stage_inst_dmem_n17976), .ZN(MEM_stage_inst_dmem_n10386) );
NAND2_X1 MEM_stage_inst_dmem_U16443 ( .A1(EX_pipeline_reg_out_12), .A2(MEM_stage_inst_dmem_n17991), .ZN(MEM_stage_inst_dmem_n17976) );
NAND2_X1 MEM_stage_inst_dmem_U16442 ( .A1(MEM_stage_inst_dmem_ram_2135), .A2(MEM_stage_inst_dmem_n17990), .ZN(MEM_stage_inst_dmem_n17977) );
NAND2_X1 MEM_stage_inst_dmem_U16441 ( .A1(MEM_stage_inst_dmem_n17975), .A2(MEM_stage_inst_dmem_n17974), .ZN(MEM_stage_inst_dmem_n10387) );
NAND2_X1 MEM_stage_inst_dmem_U16440 ( .A1(EX_pipeline_reg_out_13), .A2(MEM_stage_inst_dmem_n17991), .ZN(MEM_stage_inst_dmem_n17974) );
NAND2_X1 MEM_stage_inst_dmem_U16439 ( .A1(MEM_stage_inst_dmem_ram_2136), .A2(MEM_stage_inst_dmem_n17990), .ZN(MEM_stage_inst_dmem_n17975) );
NAND2_X1 MEM_stage_inst_dmem_U16438 ( .A1(MEM_stage_inst_dmem_n17973), .A2(MEM_stage_inst_dmem_n17972), .ZN(MEM_stage_inst_dmem_n10388) );
NAND2_X1 MEM_stage_inst_dmem_U16437 ( .A1(EX_pipeline_reg_out_14), .A2(MEM_stage_inst_dmem_n17991), .ZN(MEM_stage_inst_dmem_n17972) );
NAND2_X1 MEM_stage_inst_dmem_U16436 ( .A1(MEM_stage_inst_dmem_ram_2137), .A2(MEM_stage_inst_dmem_n17990), .ZN(MEM_stage_inst_dmem_n17973) );
NAND2_X1 MEM_stage_inst_dmem_U16435 ( .A1(MEM_stage_inst_dmem_n17971), .A2(MEM_stage_inst_dmem_n17970), .ZN(MEM_stage_inst_dmem_n10389) );
NAND2_X1 MEM_stage_inst_dmem_U16434 ( .A1(EX_pipeline_reg_out_15), .A2(MEM_stage_inst_dmem_n17991), .ZN(MEM_stage_inst_dmem_n17970) );
NAND2_X1 MEM_stage_inst_dmem_U16433 ( .A1(MEM_stage_inst_dmem_ram_2138), .A2(MEM_stage_inst_dmem_n17990), .ZN(MEM_stage_inst_dmem_n17971) );
NAND2_X1 MEM_stage_inst_dmem_U16432 ( .A1(MEM_stage_inst_dmem_n17969), .A2(MEM_stage_inst_dmem_n17968), .ZN(MEM_stage_inst_dmem_n10390) );
NAND2_X1 MEM_stage_inst_dmem_U16431 ( .A1(EX_pipeline_reg_out_16), .A2(MEM_stage_inst_dmem_n17991), .ZN(MEM_stage_inst_dmem_n17968) );
NAND2_X1 MEM_stage_inst_dmem_U16430 ( .A1(MEM_stage_inst_dmem_ram_2139), .A2(MEM_stage_inst_dmem_n17990), .ZN(MEM_stage_inst_dmem_n17969) );
NAND2_X1 MEM_stage_inst_dmem_U16429 ( .A1(MEM_stage_inst_dmem_n17967), .A2(MEM_stage_inst_dmem_n17966), .ZN(MEM_stage_inst_dmem_n10391) );
NAND2_X1 MEM_stage_inst_dmem_U16428 ( .A1(EX_pipeline_reg_out_17), .A2(MEM_stage_inst_dmem_n17991), .ZN(MEM_stage_inst_dmem_n17966) );
NAND2_X1 MEM_stage_inst_dmem_U16427 ( .A1(MEM_stage_inst_dmem_ram_2140), .A2(MEM_stage_inst_dmem_n17990), .ZN(MEM_stage_inst_dmem_n17967) );
NAND2_X1 MEM_stage_inst_dmem_U16426 ( .A1(MEM_stage_inst_dmem_n17965), .A2(MEM_stage_inst_dmem_n17964), .ZN(MEM_stage_inst_dmem_n10392) );
NAND2_X1 MEM_stage_inst_dmem_U16425 ( .A1(EX_pipeline_reg_out_18), .A2(MEM_stage_inst_dmem_n17991), .ZN(MEM_stage_inst_dmem_n17964) );
NAND2_X1 MEM_stage_inst_dmem_U16424 ( .A1(MEM_stage_inst_dmem_ram_2141), .A2(MEM_stage_inst_dmem_n17990), .ZN(MEM_stage_inst_dmem_n17965) );
NAND2_X1 MEM_stage_inst_dmem_U16423 ( .A1(MEM_stage_inst_dmem_n17963), .A2(MEM_stage_inst_dmem_n17962), .ZN(MEM_stage_inst_dmem_n10393) );
NAND2_X1 MEM_stage_inst_dmem_U16422 ( .A1(EX_pipeline_reg_out_19), .A2(MEM_stage_inst_dmem_n17991), .ZN(MEM_stage_inst_dmem_n17962) );
NAND2_X1 MEM_stage_inst_dmem_U16421 ( .A1(MEM_stage_inst_dmem_ram_2142), .A2(MEM_stage_inst_dmem_n17990), .ZN(MEM_stage_inst_dmem_n17963) );
NAND2_X1 MEM_stage_inst_dmem_U16420 ( .A1(MEM_stage_inst_dmem_n17961), .A2(MEM_stage_inst_dmem_n17960), .ZN(MEM_stage_inst_dmem_n10394) );
NAND2_X1 MEM_stage_inst_dmem_U16419 ( .A1(EX_pipeline_reg_out_20), .A2(MEM_stage_inst_dmem_n17991), .ZN(MEM_stage_inst_dmem_n17960) );
INV_X1 MEM_stage_inst_dmem_U16418 ( .A(MEM_stage_inst_dmem_n17990), .ZN(MEM_stage_inst_dmem_n17991) );
NAND2_X1 MEM_stage_inst_dmem_U16417 ( .A1(MEM_stage_inst_dmem_ram_2143), .A2(MEM_stage_inst_dmem_n17990), .ZN(MEM_stage_inst_dmem_n17961) );
NAND2_X1 MEM_stage_inst_dmem_U16416 ( .A1(MEM_stage_inst_dmem_n21284), .A2(MEM_stage_inst_dmem_n18138), .ZN(MEM_stage_inst_dmem_n17990) );
NAND2_X1 MEM_stage_inst_dmem_U16415 ( .A1(MEM_stage_inst_dmem_n17959), .A2(MEM_stage_inst_dmem_n17958), .ZN(MEM_stage_inst_dmem_n10395) );
NAND2_X1 MEM_stage_inst_dmem_U16414 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n17957), .ZN(MEM_stage_inst_dmem_n17958) );
NAND2_X1 MEM_stage_inst_dmem_U16413 ( .A1(MEM_stage_inst_dmem_ram_2144), .A2(MEM_stage_inst_dmem_n17956), .ZN(MEM_stage_inst_dmem_n17959) );
NAND2_X1 MEM_stage_inst_dmem_U16412 ( .A1(MEM_stage_inst_dmem_n17955), .A2(MEM_stage_inst_dmem_n17954), .ZN(MEM_stage_inst_dmem_n10396) );
NAND2_X1 MEM_stage_inst_dmem_U16411 ( .A1(EX_pipeline_reg_out_6), .A2(MEM_stage_inst_dmem_n17957), .ZN(MEM_stage_inst_dmem_n17954) );
NAND2_X1 MEM_stage_inst_dmem_U16410 ( .A1(MEM_stage_inst_dmem_ram_2145), .A2(MEM_stage_inst_dmem_n17956), .ZN(MEM_stage_inst_dmem_n17955) );
NAND2_X1 MEM_stage_inst_dmem_U16409 ( .A1(MEM_stage_inst_dmem_n17953), .A2(MEM_stage_inst_dmem_n17952), .ZN(MEM_stage_inst_dmem_n10397) );
NAND2_X1 MEM_stage_inst_dmem_U16408 ( .A1(MEM_stage_inst_dmem_n18027), .A2(MEM_stage_inst_dmem_n17957), .ZN(MEM_stage_inst_dmem_n17952) );
NAND2_X1 MEM_stage_inst_dmem_U16407 ( .A1(MEM_stage_inst_dmem_ram_2146), .A2(MEM_stage_inst_dmem_n17956), .ZN(MEM_stage_inst_dmem_n17953) );
NAND2_X1 MEM_stage_inst_dmem_U16406 ( .A1(MEM_stage_inst_dmem_n17951), .A2(MEM_stage_inst_dmem_n17950), .ZN(MEM_stage_inst_dmem_n10398) );
NAND2_X1 MEM_stage_inst_dmem_U16405 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n17957), .ZN(MEM_stage_inst_dmem_n17950) );
NAND2_X1 MEM_stage_inst_dmem_U16404 ( .A1(MEM_stage_inst_dmem_ram_2147), .A2(MEM_stage_inst_dmem_n17956), .ZN(MEM_stage_inst_dmem_n17951) );
NAND2_X1 MEM_stage_inst_dmem_U16403 ( .A1(MEM_stage_inst_dmem_n17949), .A2(MEM_stage_inst_dmem_n17948), .ZN(MEM_stage_inst_dmem_n10399) );
NAND2_X1 MEM_stage_inst_dmem_U16402 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n17957), .ZN(MEM_stage_inst_dmem_n17948) );
NAND2_X1 MEM_stage_inst_dmem_U16401 ( .A1(MEM_stage_inst_dmem_ram_2148), .A2(MEM_stage_inst_dmem_n17956), .ZN(MEM_stage_inst_dmem_n17949) );
NAND2_X1 MEM_stage_inst_dmem_U16400 ( .A1(MEM_stage_inst_dmem_n17947), .A2(MEM_stage_inst_dmem_n17946), .ZN(MEM_stage_inst_dmem_n10400) );
NAND2_X1 MEM_stage_inst_dmem_U16399 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n17957), .ZN(MEM_stage_inst_dmem_n17946) );
NAND2_X1 MEM_stage_inst_dmem_U16398 ( .A1(MEM_stage_inst_dmem_ram_2149), .A2(MEM_stage_inst_dmem_n17956), .ZN(MEM_stage_inst_dmem_n17947) );
NAND2_X1 MEM_stage_inst_dmem_U16397 ( .A1(MEM_stage_inst_dmem_n17945), .A2(MEM_stage_inst_dmem_n17944), .ZN(MEM_stage_inst_dmem_n10401) );
NAND2_X1 MEM_stage_inst_dmem_U16396 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n17957), .ZN(MEM_stage_inst_dmem_n17944) );
NAND2_X1 MEM_stage_inst_dmem_U16395 ( .A1(MEM_stage_inst_dmem_ram_2150), .A2(MEM_stage_inst_dmem_n17956), .ZN(MEM_stage_inst_dmem_n17945) );
NAND2_X1 MEM_stage_inst_dmem_U16394 ( .A1(MEM_stage_inst_dmem_n17943), .A2(MEM_stage_inst_dmem_n17942), .ZN(MEM_stage_inst_dmem_n10402) );
NAND2_X1 MEM_stage_inst_dmem_U16393 ( .A1(MEM_stage_inst_dmem_n16361), .A2(MEM_stage_inst_dmem_n17957), .ZN(MEM_stage_inst_dmem_n17942) );
NAND2_X1 MEM_stage_inst_dmem_U16392 ( .A1(MEM_stage_inst_dmem_ram_2151), .A2(MEM_stage_inst_dmem_n17956), .ZN(MEM_stage_inst_dmem_n17943) );
NAND2_X1 MEM_stage_inst_dmem_U16391 ( .A1(MEM_stage_inst_dmem_n17941), .A2(MEM_stage_inst_dmem_n17940), .ZN(MEM_stage_inst_dmem_n10403) );
NAND2_X1 MEM_stage_inst_dmem_U16390 ( .A1(MEM_stage_inst_dmem_n18013), .A2(MEM_stage_inst_dmem_n17957), .ZN(MEM_stage_inst_dmem_n17940) );
NAND2_X1 MEM_stage_inst_dmem_U16389 ( .A1(MEM_stage_inst_dmem_ram_2152), .A2(MEM_stage_inst_dmem_n17956), .ZN(MEM_stage_inst_dmem_n17941) );
NAND2_X1 MEM_stage_inst_dmem_U16388 ( .A1(MEM_stage_inst_dmem_n17939), .A2(MEM_stage_inst_dmem_n17938), .ZN(MEM_stage_inst_dmem_n10404) );
NAND2_X1 MEM_stage_inst_dmem_U16387 ( .A1(MEM_stage_inst_dmem_n96), .A2(MEM_stage_inst_dmem_n17957), .ZN(MEM_stage_inst_dmem_n17938) );
NAND2_X1 MEM_stage_inst_dmem_U16386 ( .A1(MEM_stage_inst_dmem_ram_2153), .A2(MEM_stage_inst_dmem_n17956), .ZN(MEM_stage_inst_dmem_n17939) );
NAND2_X1 MEM_stage_inst_dmem_U16385 ( .A1(MEM_stage_inst_dmem_n17937), .A2(MEM_stage_inst_dmem_n17936), .ZN(MEM_stage_inst_dmem_n10405) );
NAND2_X1 MEM_stage_inst_dmem_U16384 ( .A1(MEM_stage_inst_dmem_n18007), .A2(MEM_stage_inst_dmem_n17957), .ZN(MEM_stage_inst_dmem_n17936) );
NAND2_X1 MEM_stage_inst_dmem_U16383 ( .A1(MEM_stage_inst_dmem_ram_2154), .A2(MEM_stage_inst_dmem_n17956), .ZN(MEM_stage_inst_dmem_n17937) );
NAND2_X1 MEM_stage_inst_dmem_U16382 ( .A1(MEM_stage_inst_dmem_n17935), .A2(MEM_stage_inst_dmem_n17934), .ZN(MEM_stage_inst_dmem_n10406) );
NAND2_X1 MEM_stage_inst_dmem_U16381 ( .A1(MEM_stage_inst_dmem_n18004), .A2(MEM_stage_inst_dmem_n17957), .ZN(MEM_stage_inst_dmem_n17934) );
NAND2_X1 MEM_stage_inst_dmem_U16380 ( .A1(MEM_stage_inst_dmem_ram_2155), .A2(MEM_stage_inst_dmem_n17956), .ZN(MEM_stage_inst_dmem_n17935) );
NAND2_X1 MEM_stage_inst_dmem_U16379 ( .A1(MEM_stage_inst_dmem_n17933), .A2(MEM_stage_inst_dmem_n17932), .ZN(MEM_stage_inst_dmem_n10407) );
NAND2_X1 MEM_stage_inst_dmem_U16378 ( .A1(MEM_stage_inst_dmem_n18001), .A2(MEM_stage_inst_dmem_n17957), .ZN(MEM_stage_inst_dmem_n17932) );
NAND2_X1 MEM_stage_inst_dmem_U16377 ( .A1(MEM_stage_inst_dmem_ram_2156), .A2(MEM_stage_inst_dmem_n17956), .ZN(MEM_stage_inst_dmem_n17933) );
NAND2_X1 MEM_stage_inst_dmem_U16376 ( .A1(MEM_stage_inst_dmem_n17931), .A2(MEM_stage_inst_dmem_n17930), .ZN(MEM_stage_inst_dmem_n10408) );
NAND2_X1 MEM_stage_inst_dmem_U16375 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n17957), .ZN(MEM_stage_inst_dmem_n17930) );
NAND2_X1 MEM_stage_inst_dmem_U16374 ( .A1(MEM_stage_inst_dmem_ram_2157), .A2(MEM_stage_inst_dmem_n17956), .ZN(MEM_stage_inst_dmem_n17931) );
NAND2_X1 MEM_stage_inst_dmem_U16373 ( .A1(MEM_stage_inst_dmem_n17929), .A2(MEM_stage_inst_dmem_n17928), .ZN(MEM_stage_inst_dmem_n10409) );
NAND2_X1 MEM_stage_inst_dmem_U16372 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n17957), .ZN(MEM_stage_inst_dmem_n17928) );
NAND2_X1 MEM_stage_inst_dmem_U16371 ( .A1(MEM_stage_inst_dmem_ram_2158), .A2(MEM_stage_inst_dmem_n17956), .ZN(MEM_stage_inst_dmem_n17929) );
NAND2_X1 MEM_stage_inst_dmem_U16370 ( .A1(MEM_stage_inst_dmem_n17927), .A2(MEM_stage_inst_dmem_n17926), .ZN(MEM_stage_inst_dmem_n10410) );
NAND2_X1 MEM_stage_inst_dmem_U16369 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n17957), .ZN(MEM_stage_inst_dmem_n17926) );
INV_X1 MEM_stage_inst_dmem_U16368 ( .A(MEM_stage_inst_dmem_n17956), .ZN(MEM_stage_inst_dmem_n17957) );
NAND2_X1 MEM_stage_inst_dmem_U16367 ( .A1(MEM_stage_inst_dmem_ram_2159), .A2(MEM_stage_inst_dmem_n17956), .ZN(MEM_stage_inst_dmem_n17927) );
NAND2_X1 MEM_stage_inst_dmem_U16366 ( .A1(MEM_stage_inst_dmem_n21249), .A2(MEM_stage_inst_dmem_n18138), .ZN(MEM_stage_inst_dmem_n17956) );
NAND2_X1 MEM_stage_inst_dmem_U16365 ( .A1(MEM_stage_inst_dmem_n17925), .A2(MEM_stage_inst_dmem_n17924), .ZN(MEM_stage_inst_dmem_n10411) );
NAND2_X1 MEM_stage_inst_dmem_U16364 ( .A1(EX_pipeline_reg_out_5), .A2(MEM_stage_inst_dmem_n17923), .ZN(MEM_stage_inst_dmem_n17924) );
NAND2_X1 MEM_stage_inst_dmem_U16363 ( .A1(MEM_stage_inst_dmem_ram_2160), .A2(MEM_stage_inst_dmem_n17922), .ZN(MEM_stage_inst_dmem_n17925) );
NAND2_X1 MEM_stage_inst_dmem_U16362 ( .A1(MEM_stage_inst_dmem_n17921), .A2(MEM_stage_inst_dmem_n17920), .ZN(MEM_stage_inst_dmem_n10412) );
NAND2_X1 MEM_stage_inst_dmem_U16361 ( .A1(EX_pipeline_reg_out_6), .A2(MEM_stage_inst_dmem_n17923), .ZN(MEM_stage_inst_dmem_n17920) );
NAND2_X1 MEM_stage_inst_dmem_U16360 ( .A1(MEM_stage_inst_dmem_ram_2161), .A2(MEM_stage_inst_dmem_n17922), .ZN(MEM_stage_inst_dmem_n17921) );
NAND2_X1 MEM_stage_inst_dmem_U16359 ( .A1(MEM_stage_inst_dmem_n17919), .A2(MEM_stage_inst_dmem_n17918), .ZN(MEM_stage_inst_dmem_n10413) );
NAND2_X1 MEM_stage_inst_dmem_U16358 ( .A1(EX_pipeline_reg_out_7), .A2(MEM_stage_inst_dmem_n17923), .ZN(MEM_stage_inst_dmem_n17918) );
NAND2_X1 MEM_stage_inst_dmem_U16357 ( .A1(MEM_stage_inst_dmem_ram_2162), .A2(MEM_stage_inst_dmem_n17922), .ZN(MEM_stage_inst_dmem_n17919) );
NAND2_X1 MEM_stage_inst_dmem_U16356 ( .A1(MEM_stage_inst_dmem_n17917), .A2(MEM_stage_inst_dmem_n17916), .ZN(MEM_stage_inst_dmem_n10414) );
NAND2_X1 MEM_stage_inst_dmem_U16355 ( .A1(EX_pipeline_reg_out_8), .A2(MEM_stage_inst_dmem_n17923), .ZN(MEM_stage_inst_dmem_n17916) );
NAND2_X1 MEM_stage_inst_dmem_U16354 ( .A1(MEM_stage_inst_dmem_ram_2163), .A2(MEM_stage_inst_dmem_n17922), .ZN(MEM_stage_inst_dmem_n17917) );
NAND2_X1 MEM_stage_inst_dmem_U16353 ( .A1(MEM_stage_inst_dmem_n17915), .A2(MEM_stage_inst_dmem_n17914), .ZN(MEM_stage_inst_dmem_n10415) );
NAND2_X1 MEM_stage_inst_dmem_U16352 ( .A1(EX_pipeline_reg_out_9), .A2(MEM_stage_inst_dmem_n17923), .ZN(MEM_stage_inst_dmem_n17914) );
NAND2_X1 MEM_stage_inst_dmem_U16351 ( .A1(MEM_stage_inst_dmem_ram_2164), .A2(MEM_stage_inst_dmem_n17922), .ZN(MEM_stage_inst_dmem_n17915) );
NAND2_X1 MEM_stage_inst_dmem_U16350 ( .A1(MEM_stage_inst_dmem_n17913), .A2(MEM_stage_inst_dmem_n17912), .ZN(MEM_stage_inst_dmem_n10416) );
NAND2_X1 MEM_stage_inst_dmem_U16349 ( .A1(EX_pipeline_reg_out_10), .A2(MEM_stage_inst_dmem_n17923), .ZN(MEM_stage_inst_dmem_n17912) );
NAND2_X1 MEM_stage_inst_dmem_U16348 ( .A1(MEM_stage_inst_dmem_ram_2165), .A2(MEM_stage_inst_dmem_n17922), .ZN(MEM_stage_inst_dmem_n17913) );
NAND2_X1 MEM_stage_inst_dmem_U16347 ( .A1(MEM_stage_inst_dmem_n17911), .A2(MEM_stage_inst_dmem_n17910), .ZN(MEM_stage_inst_dmem_n10417) );
NAND2_X1 MEM_stage_inst_dmem_U16346 ( .A1(EX_pipeline_reg_out_11), .A2(MEM_stage_inst_dmem_n17923), .ZN(MEM_stage_inst_dmem_n17910) );
NAND2_X1 MEM_stage_inst_dmem_U16345 ( .A1(MEM_stage_inst_dmem_ram_2166), .A2(MEM_stage_inst_dmem_n17922), .ZN(MEM_stage_inst_dmem_n17911) );
NAND2_X1 MEM_stage_inst_dmem_U16344 ( .A1(MEM_stage_inst_dmem_n17909), .A2(MEM_stage_inst_dmem_n17908), .ZN(MEM_stage_inst_dmem_n10418) );
NAND2_X1 MEM_stage_inst_dmem_U16343 ( .A1(EX_pipeline_reg_out_12), .A2(MEM_stage_inst_dmem_n17923), .ZN(MEM_stage_inst_dmem_n17908) );
NAND2_X1 MEM_stage_inst_dmem_U16342 ( .A1(MEM_stage_inst_dmem_ram_2167), .A2(MEM_stage_inst_dmem_n17922), .ZN(MEM_stage_inst_dmem_n17909) );
NAND2_X1 MEM_stage_inst_dmem_U16341 ( .A1(MEM_stage_inst_dmem_n17907), .A2(MEM_stage_inst_dmem_n17906), .ZN(MEM_stage_inst_dmem_n10419) );
NAND2_X1 MEM_stage_inst_dmem_U16340 ( .A1(EX_pipeline_reg_out_13), .A2(MEM_stage_inst_dmem_n17923), .ZN(MEM_stage_inst_dmem_n17906) );
NAND2_X1 MEM_stage_inst_dmem_U16339 ( .A1(MEM_stage_inst_dmem_ram_2168), .A2(MEM_stage_inst_dmem_n17922), .ZN(MEM_stage_inst_dmem_n17907) );
NAND2_X1 MEM_stage_inst_dmem_U16338 ( .A1(MEM_stage_inst_dmem_n17905), .A2(MEM_stage_inst_dmem_n17904), .ZN(MEM_stage_inst_dmem_n10420) );
NAND2_X1 MEM_stage_inst_dmem_U16337 ( .A1(EX_pipeline_reg_out_14), .A2(MEM_stage_inst_dmem_n17923), .ZN(MEM_stage_inst_dmem_n17904) );
NAND2_X1 MEM_stage_inst_dmem_U16336 ( .A1(MEM_stage_inst_dmem_ram_2169), .A2(MEM_stage_inst_dmem_n17922), .ZN(MEM_stage_inst_dmem_n17905) );
NAND2_X1 MEM_stage_inst_dmem_U16335 ( .A1(MEM_stage_inst_dmem_n17903), .A2(MEM_stage_inst_dmem_n17902), .ZN(MEM_stage_inst_dmem_n10421) );
NAND2_X1 MEM_stage_inst_dmem_U16334 ( .A1(EX_pipeline_reg_out_15), .A2(MEM_stage_inst_dmem_n17923), .ZN(MEM_stage_inst_dmem_n17902) );
NAND2_X1 MEM_stage_inst_dmem_U16333 ( .A1(MEM_stage_inst_dmem_ram_2170), .A2(MEM_stage_inst_dmem_n17922), .ZN(MEM_stage_inst_dmem_n17903) );
NAND2_X1 MEM_stage_inst_dmem_U16332 ( .A1(MEM_stage_inst_dmem_n17901), .A2(MEM_stage_inst_dmem_n17900), .ZN(MEM_stage_inst_dmem_n10422) );
NAND2_X1 MEM_stage_inst_dmem_U16331 ( .A1(EX_pipeline_reg_out_16), .A2(MEM_stage_inst_dmem_n17923), .ZN(MEM_stage_inst_dmem_n17900) );
NAND2_X1 MEM_stage_inst_dmem_U16330 ( .A1(MEM_stage_inst_dmem_ram_2171), .A2(MEM_stage_inst_dmem_n17922), .ZN(MEM_stage_inst_dmem_n17901) );
NAND2_X1 MEM_stage_inst_dmem_U16329 ( .A1(MEM_stage_inst_dmem_n17899), .A2(MEM_stage_inst_dmem_n17898), .ZN(MEM_stage_inst_dmem_n10423) );
NAND2_X1 MEM_stage_inst_dmem_U16328 ( .A1(EX_pipeline_reg_out_17), .A2(MEM_stage_inst_dmem_n17923), .ZN(MEM_stage_inst_dmem_n17898) );
NAND2_X1 MEM_stage_inst_dmem_U16327 ( .A1(MEM_stage_inst_dmem_ram_2172), .A2(MEM_stage_inst_dmem_n17922), .ZN(MEM_stage_inst_dmem_n17899) );
NAND2_X1 MEM_stage_inst_dmem_U16326 ( .A1(MEM_stage_inst_dmem_n17897), .A2(MEM_stage_inst_dmem_n17896), .ZN(MEM_stage_inst_dmem_n10424) );
NAND2_X1 MEM_stage_inst_dmem_U16325 ( .A1(EX_pipeline_reg_out_18), .A2(MEM_stage_inst_dmem_n17923), .ZN(MEM_stage_inst_dmem_n17896) );
NAND2_X1 MEM_stage_inst_dmem_U16324 ( .A1(MEM_stage_inst_dmem_ram_2173), .A2(MEM_stage_inst_dmem_n17922), .ZN(MEM_stage_inst_dmem_n17897) );
NAND2_X1 MEM_stage_inst_dmem_U16323 ( .A1(MEM_stage_inst_dmem_n17895), .A2(MEM_stage_inst_dmem_n17894), .ZN(MEM_stage_inst_dmem_n10425) );
NAND2_X1 MEM_stage_inst_dmem_U16322 ( .A1(EX_pipeline_reg_out_19), .A2(MEM_stage_inst_dmem_n17923), .ZN(MEM_stage_inst_dmem_n17894) );
NAND2_X1 MEM_stage_inst_dmem_U16321 ( .A1(MEM_stage_inst_dmem_ram_2174), .A2(MEM_stage_inst_dmem_n17922), .ZN(MEM_stage_inst_dmem_n17895) );
NAND2_X1 MEM_stage_inst_dmem_U16320 ( .A1(MEM_stage_inst_dmem_n17893), .A2(MEM_stage_inst_dmem_n17892), .ZN(MEM_stage_inst_dmem_n10426) );
NAND2_X1 MEM_stage_inst_dmem_U16319 ( .A1(EX_pipeline_reg_out_20), .A2(MEM_stage_inst_dmem_n17923), .ZN(MEM_stage_inst_dmem_n17892) );
INV_X1 MEM_stage_inst_dmem_U16318 ( .A(MEM_stage_inst_dmem_n17922), .ZN(MEM_stage_inst_dmem_n17923) );
NAND2_X1 MEM_stage_inst_dmem_U16317 ( .A1(MEM_stage_inst_dmem_ram_2175), .A2(MEM_stage_inst_dmem_n17922), .ZN(MEM_stage_inst_dmem_n17893) );
NAND2_X1 MEM_stage_inst_dmem_U16316 ( .A1(MEM_stage_inst_dmem_n21214), .A2(MEM_stage_inst_dmem_n18138), .ZN(MEM_stage_inst_dmem_n17922) );
NAND2_X1 MEM_stage_inst_dmem_U16315 ( .A1(MEM_stage_inst_dmem_n17891), .A2(MEM_stage_inst_dmem_n17890), .ZN(MEM_stage_inst_dmem_n10427) );
NAND2_X1 MEM_stage_inst_dmem_U16314 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n17889), .ZN(MEM_stage_inst_dmem_n17890) );
NAND2_X1 MEM_stage_inst_dmem_U16313 ( .A1(MEM_stage_inst_dmem_ram_2176), .A2(MEM_stage_inst_dmem_n17888), .ZN(MEM_stage_inst_dmem_n17891) );
NAND2_X1 MEM_stage_inst_dmem_U16312 ( .A1(MEM_stage_inst_dmem_n17887), .A2(MEM_stage_inst_dmem_n17886), .ZN(MEM_stage_inst_dmem_n10428) );
NAND2_X1 MEM_stage_inst_dmem_U16311 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n17889), .ZN(MEM_stage_inst_dmem_n17886) );
NAND2_X1 MEM_stage_inst_dmem_U16310 ( .A1(MEM_stage_inst_dmem_ram_2177), .A2(MEM_stage_inst_dmem_n17888), .ZN(MEM_stage_inst_dmem_n17887) );
NAND2_X1 MEM_stage_inst_dmem_U16309 ( .A1(MEM_stage_inst_dmem_n17885), .A2(MEM_stage_inst_dmem_n17884), .ZN(MEM_stage_inst_dmem_n10429) );
NAND2_X1 MEM_stage_inst_dmem_U16308 ( .A1(MEM_stage_inst_dmem_n18027), .A2(MEM_stage_inst_dmem_n17889), .ZN(MEM_stage_inst_dmem_n17884) );
NAND2_X1 MEM_stage_inst_dmem_U16307 ( .A1(MEM_stage_inst_dmem_ram_2178), .A2(MEM_stage_inst_dmem_n17888), .ZN(MEM_stage_inst_dmem_n17885) );
NAND2_X1 MEM_stage_inst_dmem_U16306 ( .A1(MEM_stage_inst_dmem_n17883), .A2(MEM_stage_inst_dmem_n17882), .ZN(MEM_stage_inst_dmem_n10430) );
NAND2_X1 MEM_stage_inst_dmem_U16305 ( .A1(EX_pipeline_reg_out_8), .A2(MEM_stage_inst_dmem_n17889), .ZN(MEM_stage_inst_dmem_n17882) );
NAND2_X1 MEM_stage_inst_dmem_U16304 ( .A1(MEM_stage_inst_dmem_ram_2179), .A2(MEM_stage_inst_dmem_n17888), .ZN(MEM_stage_inst_dmem_n17883) );
NAND2_X1 MEM_stage_inst_dmem_U16303 ( .A1(MEM_stage_inst_dmem_n17881), .A2(MEM_stage_inst_dmem_n17880), .ZN(MEM_stage_inst_dmem_n10431) );
NAND2_X1 MEM_stage_inst_dmem_U16302 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n17889), .ZN(MEM_stage_inst_dmem_n17880) );
NAND2_X1 MEM_stage_inst_dmem_U16301 ( .A1(MEM_stage_inst_dmem_ram_2180), .A2(MEM_stage_inst_dmem_n17888), .ZN(MEM_stage_inst_dmem_n17881) );
NAND2_X1 MEM_stage_inst_dmem_U16300 ( .A1(MEM_stage_inst_dmem_n17879), .A2(MEM_stage_inst_dmem_n17878), .ZN(MEM_stage_inst_dmem_n10432) );
NAND2_X1 MEM_stage_inst_dmem_U16299 ( .A1(EX_pipeline_reg_out_10), .A2(MEM_stage_inst_dmem_n17889), .ZN(MEM_stage_inst_dmem_n17878) );
NAND2_X1 MEM_stage_inst_dmem_U16298 ( .A1(MEM_stage_inst_dmem_ram_2181), .A2(MEM_stage_inst_dmem_n17888), .ZN(MEM_stage_inst_dmem_n17879) );
NAND2_X1 MEM_stage_inst_dmem_U16297 ( .A1(MEM_stage_inst_dmem_n17877), .A2(MEM_stage_inst_dmem_n17876), .ZN(MEM_stage_inst_dmem_n10433) );
NAND2_X1 MEM_stage_inst_dmem_U16296 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n17889), .ZN(MEM_stage_inst_dmem_n17876) );
NAND2_X1 MEM_stage_inst_dmem_U16295 ( .A1(MEM_stage_inst_dmem_ram_2182), .A2(MEM_stage_inst_dmem_n17888), .ZN(MEM_stage_inst_dmem_n17877) );
NAND2_X1 MEM_stage_inst_dmem_U16294 ( .A1(MEM_stage_inst_dmem_n17875), .A2(MEM_stage_inst_dmem_n17874), .ZN(MEM_stage_inst_dmem_n10434) );
NAND2_X1 MEM_stage_inst_dmem_U16293 ( .A1(MEM_stage_inst_dmem_n112), .A2(MEM_stage_inst_dmem_n17889), .ZN(MEM_stage_inst_dmem_n17874) );
NAND2_X1 MEM_stage_inst_dmem_U16292 ( .A1(MEM_stage_inst_dmem_ram_2183), .A2(MEM_stage_inst_dmem_n17888), .ZN(MEM_stage_inst_dmem_n17875) );
NAND2_X1 MEM_stage_inst_dmem_U16291 ( .A1(MEM_stage_inst_dmem_n17873), .A2(MEM_stage_inst_dmem_n17872), .ZN(MEM_stage_inst_dmem_n10435) );
NAND2_X1 MEM_stage_inst_dmem_U16290 ( .A1(MEM_stage_inst_dmem_n18013), .A2(MEM_stage_inst_dmem_n17889), .ZN(MEM_stage_inst_dmem_n17872) );
NAND2_X1 MEM_stage_inst_dmem_U16289 ( .A1(MEM_stage_inst_dmem_ram_2184), .A2(MEM_stage_inst_dmem_n17888), .ZN(MEM_stage_inst_dmem_n17873) );
NAND2_X1 MEM_stage_inst_dmem_U16288 ( .A1(MEM_stage_inst_dmem_n17871), .A2(MEM_stage_inst_dmem_n17870), .ZN(MEM_stage_inst_dmem_n10436) );
NAND2_X1 MEM_stage_inst_dmem_U16287 ( .A1(MEM_stage_inst_dmem_n96), .A2(MEM_stage_inst_dmem_n17889), .ZN(MEM_stage_inst_dmem_n17870) );
NAND2_X1 MEM_stage_inst_dmem_U16286 ( .A1(MEM_stage_inst_dmem_ram_2185), .A2(MEM_stage_inst_dmem_n17888), .ZN(MEM_stage_inst_dmem_n17871) );
NAND2_X1 MEM_stage_inst_dmem_U16285 ( .A1(MEM_stage_inst_dmem_n17869), .A2(MEM_stage_inst_dmem_n17868), .ZN(MEM_stage_inst_dmem_n10437) );
NAND2_X1 MEM_stage_inst_dmem_U16284 ( .A1(MEM_stage_inst_dmem_n18007), .A2(MEM_stage_inst_dmem_n17889), .ZN(MEM_stage_inst_dmem_n17868) );
NAND2_X1 MEM_stage_inst_dmem_U16283 ( .A1(MEM_stage_inst_dmem_ram_2186), .A2(MEM_stage_inst_dmem_n17888), .ZN(MEM_stage_inst_dmem_n17869) );
NAND2_X1 MEM_stage_inst_dmem_U16282 ( .A1(MEM_stage_inst_dmem_n17867), .A2(MEM_stage_inst_dmem_n17866), .ZN(MEM_stage_inst_dmem_n10438) );
NAND2_X1 MEM_stage_inst_dmem_U16281 ( .A1(MEM_stage_inst_dmem_n18004), .A2(MEM_stage_inst_dmem_n17889), .ZN(MEM_stage_inst_dmem_n17866) );
NAND2_X1 MEM_stage_inst_dmem_U16280 ( .A1(MEM_stage_inst_dmem_ram_2187), .A2(MEM_stage_inst_dmem_n17888), .ZN(MEM_stage_inst_dmem_n17867) );
NAND2_X1 MEM_stage_inst_dmem_U16279 ( .A1(MEM_stage_inst_dmem_n17865), .A2(MEM_stage_inst_dmem_n17864), .ZN(MEM_stage_inst_dmem_n10439) );
NAND2_X1 MEM_stage_inst_dmem_U16278 ( .A1(MEM_stage_inst_dmem_n18001), .A2(MEM_stage_inst_dmem_n17889), .ZN(MEM_stage_inst_dmem_n17864) );
NAND2_X1 MEM_stage_inst_dmem_U16277 ( .A1(MEM_stage_inst_dmem_ram_2188), .A2(MEM_stage_inst_dmem_n17888), .ZN(MEM_stage_inst_dmem_n17865) );
NAND2_X1 MEM_stage_inst_dmem_U16276 ( .A1(MEM_stage_inst_dmem_n17863), .A2(MEM_stage_inst_dmem_n17862), .ZN(MEM_stage_inst_dmem_n10440) );
NAND2_X1 MEM_stage_inst_dmem_U16275 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n17889), .ZN(MEM_stage_inst_dmem_n17862) );
NAND2_X1 MEM_stage_inst_dmem_U16274 ( .A1(MEM_stage_inst_dmem_ram_2189), .A2(MEM_stage_inst_dmem_n17888), .ZN(MEM_stage_inst_dmem_n17863) );
NAND2_X1 MEM_stage_inst_dmem_U16273 ( .A1(MEM_stage_inst_dmem_n17861), .A2(MEM_stage_inst_dmem_n17860), .ZN(MEM_stage_inst_dmem_n10441) );
NAND2_X1 MEM_stage_inst_dmem_U16272 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n17889), .ZN(MEM_stage_inst_dmem_n17860) );
NAND2_X1 MEM_stage_inst_dmem_U16271 ( .A1(MEM_stage_inst_dmem_ram_2190), .A2(MEM_stage_inst_dmem_n17888), .ZN(MEM_stage_inst_dmem_n17861) );
NAND2_X1 MEM_stage_inst_dmem_U16270 ( .A1(MEM_stage_inst_dmem_n17859), .A2(MEM_stage_inst_dmem_n17858), .ZN(MEM_stage_inst_dmem_n10442) );
NAND2_X1 MEM_stage_inst_dmem_U16269 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n17889), .ZN(MEM_stage_inst_dmem_n17858) );
NAND2_X1 MEM_stage_inst_dmem_U16268 ( .A1(MEM_stage_inst_dmem_ram_2191), .A2(MEM_stage_inst_dmem_n17888), .ZN(MEM_stage_inst_dmem_n17859) );
NAND2_X1 MEM_stage_inst_dmem_U16267 ( .A1(MEM_stage_inst_dmem_n21179), .A2(MEM_stage_inst_dmem_n18138), .ZN(MEM_stage_inst_dmem_n17888) );
NAND2_X1 MEM_stage_inst_dmem_U16266 ( .A1(MEM_stage_inst_dmem_n17857), .A2(MEM_stage_inst_dmem_n17856), .ZN(MEM_stage_inst_dmem_n10443) );
NAND2_X1 MEM_stage_inst_dmem_U16265 ( .A1(EX_pipeline_reg_out_5), .A2(MEM_stage_inst_dmem_n17855), .ZN(MEM_stage_inst_dmem_n17856) );
NAND2_X1 MEM_stage_inst_dmem_U16264 ( .A1(MEM_stage_inst_dmem_ram_2192), .A2(MEM_stage_inst_dmem_n17854), .ZN(MEM_stage_inst_dmem_n17857) );
NAND2_X1 MEM_stage_inst_dmem_U16263 ( .A1(MEM_stage_inst_dmem_n17853), .A2(MEM_stage_inst_dmem_n17852), .ZN(MEM_stage_inst_dmem_n10444) );
NAND2_X1 MEM_stage_inst_dmem_U16262 ( .A1(EX_pipeline_reg_out_6), .A2(MEM_stage_inst_dmem_n17855), .ZN(MEM_stage_inst_dmem_n17852) );
NAND2_X1 MEM_stage_inst_dmem_U16261 ( .A1(MEM_stage_inst_dmem_ram_2193), .A2(MEM_stage_inst_dmem_n17854), .ZN(MEM_stage_inst_dmem_n17853) );
NAND2_X1 MEM_stage_inst_dmem_U16260 ( .A1(MEM_stage_inst_dmem_n17851), .A2(MEM_stage_inst_dmem_n17850), .ZN(MEM_stage_inst_dmem_n10445) );
NAND2_X1 MEM_stage_inst_dmem_U16259 ( .A1(EX_pipeline_reg_out_7), .A2(MEM_stage_inst_dmem_n17855), .ZN(MEM_stage_inst_dmem_n17850) );
NAND2_X1 MEM_stage_inst_dmem_U16258 ( .A1(MEM_stage_inst_dmem_ram_2194), .A2(MEM_stage_inst_dmem_n17854), .ZN(MEM_stage_inst_dmem_n17851) );
NAND2_X1 MEM_stage_inst_dmem_U16257 ( .A1(MEM_stage_inst_dmem_n17849), .A2(MEM_stage_inst_dmem_n17848), .ZN(MEM_stage_inst_dmem_n10446) );
NAND2_X1 MEM_stage_inst_dmem_U16256 ( .A1(EX_pipeline_reg_out_8), .A2(MEM_stage_inst_dmem_n17855), .ZN(MEM_stage_inst_dmem_n17848) );
NAND2_X1 MEM_stage_inst_dmem_U16255 ( .A1(MEM_stage_inst_dmem_ram_2195), .A2(MEM_stage_inst_dmem_n17854), .ZN(MEM_stage_inst_dmem_n17849) );
NAND2_X1 MEM_stage_inst_dmem_U16254 ( .A1(MEM_stage_inst_dmem_n17847), .A2(MEM_stage_inst_dmem_n17846), .ZN(MEM_stage_inst_dmem_n10447) );
NAND2_X1 MEM_stage_inst_dmem_U16253 ( .A1(EX_pipeline_reg_out_9), .A2(MEM_stage_inst_dmem_n17855), .ZN(MEM_stage_inst_dmem_n17846) );
NAND2_X1 MEM_stage_inst_dmem_U16252 ( .A1(MEM_stage_inst_dmem_ram_2196), .A2(MEM_stage_inst_dmem_n17854), .ZN(MEM_stage_inst_dmem_n17847) );
NAND2_X1 MEM_stage_inst_dmem_U16251 ( .A1(MEM_stage_inst_dmem_n17845), .A2(MEM_stage_inst_dmem_n17844), .ZN(MEM_stage_inst_dmem_n10448) );
NAND2_X1 MEM_stage_inst_dmem_U16250 ( .A1(EX_pipeline_reg_out_10), .A2(MEM_stage_inst_dmem_n17855), .ZN(MEM_stage_inst_dmem_n17844) );
NAND2_X1 MEM_stage_inst_dmem_U16249 ( .A1(MEM_stage_inst_dmem_ram_2197), .A2(MEM_stage_inst_dmem_n17854), .ZN(MEM_stage_inst_dmem_n17845) );
NAND2_X1 MEM_stage_inst_dmem_U16248 ( .A1(MEM_stage_inst_dmem_n17843), .A2(MEM_stage_inst_dmem_n17842), .ZN(MEM_stage_inst_dmem_n10449) );
NAND2_X1 MEM_stage_inst_dmem_U16247 ( .A1(EX_pipeline_reg_out_11), .A2(MEM_stage_inst_dmem_n17855), .ZN(MEM_stage_inst_dmem_n17842) );
NAND2_X1 MEM_stage_inst_dmem_U16246 ( .A1(MEM_stage_inst_dmem_ram_2198), .A2(MEM_stage_inst_dmem_n17854), .ZN(MEM_stage_inst_dmem_n17843) );
NAND2_X1 MEM_stage_inst_dmem_U16245 ( .A1(MEM_stage_inst_dmem_n17841), .A2(MEM_stage_inst_dmem_n17840), .ZN(MEM_stage_inst_dmem_n10450) );
NAND2_X1 MEM_stage_inst_dmem_U16244 ( .A1(EX_pipeline_reg_out_12), .A2(MEM_stage_inst_dmem_n17855), .ZN(MEM_stage_inst_dmem_n17840) );
NAND2_X1 MEM_stage_inst_dmem_U16243 ( .A1(MEM_stage_inst_dmem_ram_2199), .A2(MEM_stage_inst_dmem_n17854), .ZN(MEM_stage_inst_dmem_n17841) );
NAND2_X1 MEM_stage_inst_dmem_U16242 ( .A1(MEM_stage_inst_dmem_n17839), .A2(MEM_stage_inst_dmem_n17838), .ZN(MEM_stage_inst_dmem_n10451) );
NAND2_X1 MEM_stage_inst_dmem_U16241 ( .A1(EX_pipeline_reg_out_13), .A2(MEM_stage_inst_dmem_n17855), .ZN(MEM_stage_inst_dmem_n17838) );
NAND2_X1 MEM_stage_inst_dmem_U16240 ( .A1(MEM_stage_inst_dmem_ram_2200), .A2(MEM_stage_inst_dmem_n17854), .ZN(MEM_stage_inst_dmem_n17839) );
NAND2_X1 MEM_stage_inst_dmem_U16239 ( .A1(MEM_stage_inst_dmem_n17837), .A2(MEM_stage_inst_dmem_n17836), .ZN(MEM_stage_inst_dmem_n10452) );
NAND2_X1 MEM_stage_inst_dmem_U16238 ( .A1(EX_pipeline_reg_out_14), .A2(MEM_stage_inst_dmem_n17855), .ZN(MEM_stage_inst_dmem_n17836) );
NAND2_X1 MEM_stage_inst_dmem_U16237 ( .A1(MEM_stage_inst_dmem_ram_2201), .A2(MEM_stage_inst_dmem_n17854), .ZN(MEM_stage_inst_dmem_n17837) );
NAND2_X1 MEM_stage_inst_dmem_U16236 ( .A1(MEM_stage_inst_dmem_n17835), .A2(MEM_stage_inst_dmem_n17834), .ZN(MEM_stage_inst_dmem_n10453) );
NAND2_X1 MEM_stage_inst_dmem_U16235 ( .A1(EX_pipeline_reg_out_15), .A2(MEM_stage_inst_dmem_n17855), .ZN(MEM_stage_inst_dmem_n17834) );
NAND2_X1 MEM_stage_inst_dmem_U16234 ( .A1(MEM_stage_inst_dmem_ram_2202), .A2(MEM_stage_inst_dmem_n17854), .ZN(MEM_stage_inst_dmem_n17835) );
NAND2_X1 MEM_stage_inst_dmem_U16233 ( .A1(MEM_stage_inst_dmem_n17833), .A2(MEM_stage_inst_dmem_n17832), .ZN(MEM_stage_inst_dmem_n10454) );
NAND2_X1 MEM_stage_inst_dmem_U16232 ( .A1(EX_pipeline_reg_out_16), .A2(MEM_stage_inst_dmem_n17855), .ZN(MEM_stage_inst_dmem_n17832) );
NAND2_X1 MEM_stage_inst_dmem_U16231 ( .A1(MEM_stage_inst_dmem_ram_2203), .A2(MEM_stage_inst_dmem_n17854), .ZN(MEM_stage_inst_dmem_n17833) );
NAND2_X1 MEM_stage_inst_dmem_U16230 ( .A1(MEM_stage_inst_dmem_n17831), .A2(MEM_stage_inst_dmem_n17830), .ZN(MEM_stage_inst_dmem_n10455) );
NAND2_X1 MEM_stage_inst_dmem_U16229 ( .A1(EX_pipeline_reg_out_17), .A2(MEM_stage_inst_dmem_n17855), .ZN(MEM_stage_inst_dmem_n17830) );
NAND2_X1 MEM_stage_inst_dmem_U16228 ( .A1(MEM_stage_inst_dmem_ram_2204), .A2(MEM_stage_inst_dmem_n17854), .ZN(MEM_stage_inst_dmem_n17831) );
NAND2_X1 MEM_stage_inst_dmem_U16227 ( .A1(MEM_stage_inst_dmem_n17829), .A2(MEM_stage_inst_dmem_n17828), .ZN(MEM_stage_inst_dmem_n10456) );
NAND2_X1 MEM_stage_inst_dmem_U16226 ( .A1(EX_pipeline_reg_out_18), .A2(MEM_stage_inst_dmem_n17855), .ZN(MEM_stage_inst_dmem_n17828) );
NAND2_X1 MEM_stage_inst_dmem_U16225 ( .A1(MEM_stage_inst_dmem_ram_2205), .A2(MEM_stage_inst_dmem_n17854), .ZN(MEM_stage_inst_dmem_n17829) );
NAND2_X1 MEM_stage_inst_dmem_U16224 ( .A1(MEM_stage_inst_dmem_n17827), .A2(MEM_stage_inst_dmem_n17826), .ZN(MEM_stage_inst_dmem_n10457) );
NAND2_X1 MEM_stage_inst_dmem_U16223 ( .A1(EX_pipeline_reg_out_19), .A2(MEM_stage_inst_dmem_n17855), .ZN(MEM_stage_inst_dmem_n17826) );
NAND2_X1 MEM_stage_inst_dmem_U16222 ( .A1(MEM_stage_inst_dmem_ram_2206), .A2(MEM_stage_inst_dmem_n17854), .ZN(MEM_stage_inst_dmem_n17827) );
NAND2_X1 MEM_stage_inst_dmem_U16221 ( .A1(MEM_stage_inst_dmem_n17825), .A2(MEM_stage_inst_dmem_n17824), .ZN(MEM_stage_inst_dmem_n10458) );
NAND2_X1 MEM_stage_inst_dmem_U16220 ( .A1(EX_pipeline_reg_out_20), .A2(MEM_stage_inst_dmem_n17855), .ZN(MEM_stage_inst_dmem_n17824) );
INV_X1 MEM_stage_inst_dmem_U16219 ( .A(MEM_stage_inst_dmem_n17854), .ZN(MEM_stage_inst_dmem_n17855) );
NAND2_X1 MEM_stage_inst_dmem_U16218 ( .A1(MEM_stage_inst_dmem_ram_2207), .A2(MEM_stage_inst_dmem_n17854), .ZN(MEM_stage_inst_dmem_n17825) );
NAND2_X1 MEM_stage_inst_dmem_U16217 ( .A1(MEM_stage_inst_dmem_n21144), .A2(MEM_stage_inst_dmem_n18138), .ZN(MEM_stage_inst_dmem_n17854) );
NAND2_X1 MEM_stage_inst_dmem_U16216 ( .A1(MEM_stage_inst_dmem_n17823), .A2(MEM_stage_inst_dmem_n17822), .ZN(MEM_stage_inst_dmem_n10459) );
NAND2_X1 MEM_stage_inst_dmem_U16215 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n17821), .ZN(MEM_stage_inst_dmem_n17822) );
NAND2_X1 MEM_stage_inst_dmem_U16214 ( .A1(MEM_stage_inst_dmem_ram_2208), .A2(MEM_stage_inst_dmem_n17820), .ZN(MEM_stage_inst_dmem_n17823) );
NAND2_X1 MEM_stage_inst_dmem_U16213 ( .A1(MEM_stage_inst_dmem_n17819), .A2(MEM_stage_inst_dmem_n17818), .ZN(MEM_stage_inst_dmem_n10460) );
NAND2_X1 MEM_stage_inst_dmem_U16212 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n17821), .ZN(MEM_stage_inst_dmem_n17818) );
NAND2_X1 MEM_stage_inst_dmem_U16211 ( .A1(MEM_stage_inst_dmem_ram_2209), .A2(MEM_stage_inst_dmem_n17820), .ZN(MEM_stage_inst_dmem_n17819) );
NAND2_X1 MEM_stage_inst_dmem_U16210 ( .A1(MEM_stage_inst_dmem_n17817), .A2(MEM_stage_inst_dmem_n17816), .ZN(MEM_stage_inst_dmem_n10461) );
NAND2_X1 MEM_stage_inst_dmem_U16209 ( .A1(MEM_stage_inst_dmem_n18027), .A2(MEM_stage_inst_dmem_n17821), .ZN(MEM_stage_inst_dmem_n17816) );
NAND2_X1 MEM_stage_inst_dmem_U16208 ( .A1(MEM_stage_inst_dmem_ram_2210), .A2(MEM_stage_inst_dmem_n17820), .ZN(MEM_stage_inst_dmem_n17817) );
NAND2_X1 MEM_stage_inst_dmem_U16207 ( .A1(MEM_stage_inst_dmem_n17815), .A2(MEM_stage_inst_dmem_n17814), .ZN(MEM_stage_inst_dmem_n10462) );
NAND2_X1 MEM_stage_inst_dmem_U16206 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n17821), .ZN(MEM_stage_inst_dmem_n17814) );
NAND2_X1 MEM_stage_inst_dmem_U16205 ( .A1(MEM_stage_inst_dmem_ram_2211), .A2(MEM_stage_inst_dmem_n17820), .ZN(MEM_stage_inst_dmem_n17815) );
NAND2_X1 MEM_stage_inst_dmem_U16204 ( .A1(MEM_stage_inst_dmem_n17813), .A2(MEM_stage_inst_dmem_n17812), .ZN(MEM_stage_inst_dmem_n10463) );
NAND2_X1 MEM_stage_inst_dmem_U16203 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n17821), .ZN(MEM_stage_inst_dmem_n17812) );
NAND2_X1 MEM_stage_inst_dmem_U16202 ( .A1(MEM_stage_inst_dmem_ram_2212), .A2(MEM_stage_inst_dmem_n17820), .ZN(MEM_stage_inst_dmem_n17813) );
NAND2_X1 MEM_stage_inst_dmem_U16201 ( .A1(MEM_stage_inst_dmem_n17811), .A2(MEM_stage_inst_dmem_n17810), .ZN(MEM_stage_inst_dmem_n10464) );
NAND2_X1 MEM_stage_inst_dmem_U16200 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n17821), .ZN(MEM_stage_inst_dmem_n17810) );
NAND2_X1 MEM_stage_inst_dmem_U16199 ( .A1(MEM_stage_inst_dmem_ram_2213), .A2(MEM_stage_inst_dmem_n17820), .ZN(MEM_stage_inst_dmem_n17811) );
NAND2_X1 MEM_stage_inst_dmem_U16198 ( .A1(MEM_stage_inst_dmem_n17809), .A2(MEM_stage_inst_dmem_n17808), .ZN(MEM_stage_inst_dmem_n10465) );
NAND2_X1 MEM_stage_inst_dmem_U16197 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n17821), .ZN(MEM_stage_inst_dmem_n17808) );
NAND2_X1 MEM_stage_inst_dmem_U16196 ( .A1(MEM_stage_inst_dmem_ram_2214), .A2(MEM_stage_inst_dmem_n17820), .ZN(MEM_stage_inst_dmem_n17809) );
NAND2_X1 MEM_stage_inst_dmem_U16195 ( .A1(MEM_stage_inst_dmem_n17807), .A2(MEM_stage_inst_dmem_n17806), .ZN(MEM_stage_inst_dmem_n10466) );
NAND2_X1 MEM_stage_inst_dmem_U16194 ( .A1(MEM_stage_inst_dmem_n16361), .A2(MEM_stage_inst_dmem_n17821), .ZN(MEM_stage_inst_dmem_n17806) );
NAND2_X1 MEM_stage_inst_dmem_U16193 ( .A1(MEM_stage_inst_dmem_ram_2215), .A2(MEM_stage_inst_dmem_n17820), .ZN(MEM_stage_inst_dmem_n17807) );
NAND2_X1 MEM_stage_inst_dmem_U16192 ( .A1(MEM_stage_inst_dmem_n17805), .A2(MEM_stage_inst_dmem_n17804), .ZN(MEM_stage_inst_dmem_n10467) );
NAND2_X1 MEM_stage_inst_dmem_U16191 ( .A1(MEM_stage_inst_dmem_n18013), .A2(MEM_stage_inst_dmem_n17821), .ZN(MEM_stage_inst_dmem_n17804) );
NAND2_X1 MEM_stage_inst_dmem_U16190 ( .A1(MEM_stage_inst_dmem_ram_2216), .A2(MEM_stage_inst_dmem_n17820), .ZN(MEM_stage_inst_dmem_n17805) );
NAND2_X1 MEM_stage_inst_dmem_U16189 ( .A1(MEM_stage_inst_dmem_n17803), .A2(MEM_stage_inst_dmem_n17802), .ZN(MEM_stage_inst_dmem_n10468) );
NAND2_X1 MEM_stage_inst_dmem_U16188 ( .A1(MEM_stage_inst_dmem_n96), .A2(MEM_stage_inst_dmem_n17821), .ZN(MEM_stage_inst_dmem_n17802) );
NAND2_X1 MEM_stage_inst_dmem_U16187 ( .A1(MEM_stage_inst_dmem_ram_2217), .A2(MEM_stage_inst_dmem_n17820), .ZN(MEM_stage_inst_dmem_n17803) );
NAND2_X1 MEM_stage_inst_dmem_U16186 ( .A1(MEM_stage_inst_dmem_n17801), .A2(MEM_stage_inst_dmem_n17800), .ZN(MEM_stage_inst_dmem_n10469) );
NAND2_X1 MEM_stage_inst_dmem_U16185 ( .A1(MEM_stage_inst_dmem_n18007), .A2(MEM_stage_inst_dmem_n17821), .ZN(MEM_stage_inst_dmem_n17800) );
NAND2_X1 MEM_stage_inst_dmem_U16184 ( .A1(MEM_stage_inst_dmem_ram_2218), .A2(MEM_stage_inst_dmem_n17820), .ZN(MEM_stage_inst_dmem_n17801) );
NAND2_X1 MEM_stage_inst_dmem_U16183 ( .A1(MEM_stage_inst_dmem_n17799), .A2(MEM_stage_inst_dmem_n17798), .ZN(MEM_stage_inst_dmem_n10470) );
NAND2_X1 MEM_stage_inst_dmem_U16182 ( .A1(MEM_stage_inst_dmem_n18004), .A2(MEM_stage_inst_dmem_n17821), .ZN(MEM_stage_inst_dmem_n17798) );
NAND2_X1 MEM_stage_inst_dmem_U16181 ( .A1(MEM_stage_inst_dmem_ram_2219), .A2(MEM_stage_inst_dmem_n17820), .ZN(MEM_stage_inst_dmem_n17799) );
NAND2_X1 MEM_stage_inst_dmem_U16180 ( .A1(MEM_stage_inst_dmem_n17797), .A2(MEM_stage_inst_dmem_n17796), .ZN(MEM_stage_inst_dmem_n10471) );
NAND2_X1 MEM_stage_inst_dmem_U16179 ( .A1(MEM_stage_inst_dmem_n18001), .A2(MEM_stage_inst_dmem_n17821), .ZN(MEM_stage_inst_dmem_n17796) );
NAND2_X1 MEM_stage_inst_dmem_U16178 ( .A1(MEM_stage_inst_dmem_ram_2220), .A2(MEM_stage_inst_dmem_n17820), .ZN(MEM_stage_inst_dmem_n17797) );
NAND2_X1 MEM_stage_inst_dmem_U16177 ( .A1(MEM_stage_inst_dmem_n17795), .A2(MEM_stage_inst_dmem_n17794), .ZN(MEM_stage_inst_dmem_n10472) );
NAND2_X1 MEM_stage_inst_dmem_U16176 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n17821), .ZN(MEM_stage_inst_dmem_n17794) );
NAND2_X1 MEM_stage_inst_dmem_U16175 ( .A1(MEM_stage_inst_dmem_ram_2221), .A2(MEM_stage_inst_dmem_n17820), .ZN(MEM_stage_inst_dmem_n17795) );
NAND2_X1 MEM_stage_inst_dmem_U16174 ( .A1(MEM_stage_inst_dmem_n17793), .A2(MEM_stage_inst_dmem_n17792), .ZN(MEM_stage_inst_dmem_n10473) );
NAND2_X1 MEM_stage_inst_dmem_U16173 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n17821), .ZN(MEM_stage_inst_dmem_n17792) );
NAND2_X1 MEM_stage_inst_dmem_U16172 ( .A1(MEM_stage_inst_dmem_ram_2222), .A2(MEM_stage_inst_dmem_n17820), .ZN(MEM_stage_inst_dmem_n17793) );
NAND2_X1 MEM_stage_inst_dmem_U16171 ( .A1(MEM_stage_inst_dmem_n17791), .A2(MEM_stage_inst_dmem_n17790), .ZN(MEM_stage_inst_dmem_n10474) );
NAND2_X1 MEM_stage_inst_dmem_U16170 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n17821), .ZN(MEM_stage_inst_dmem_n17790) );
INV_X1 MEM_stage_inst_dmem_U16169 ( .A(MEM_stage_inst_dmem_n17820), .ZN(MEM_stage_inst_dmem_n17821) );
NAND2_X1 MEM_stage_inst_dmem_U16168 ( .A1(MEM_stage_inst_dmem_ram_2223), .A2(MEM_stage_inst_dmem_n17820), .ZN(MEM_stage_inst_dmem_n17791) );
NAND2_X1 MEM_stage_inst_dmem_U16167 ( .A1(MEM_stage_inst_dmem_n21109), .A2(MEM_stage_inst_dmem_n18138), .ZN(MEM_stage_inst_dmem_n17820) );
NAND2_X1 MEM_stage_inst_dmem_U16166 ( .A1(MEM_stage_inst_dmem_n17789), .A2(MEM_stage_inst_dmem_n17788), .ZN(MEM_stage_inst_dmem_n10475) );
NAND2_X1 MEM_stage_inst_dmem_U16165 ( .A1(EX_pipeline_reg_out_5), .A2(MEM_stage_inst_dmem_n17787), .ZN(MEM_stage_inst_dmem_n17788) );
NAND2_X1 MEM_stage_inst_dmem_U16164 ( .A1(MEM_stage_inst_dmem_ram_2224), .A2(MEM_stage_inst_dmem_n17786), .ZN(MEM_stage_inst_dmem_n17789) );
NAND2_X1 MEM_stage_inst_dmem_U16163 ( .A1(MEM_stage_inst_dmem_n17785), .A2(MEM_stage_inst_dmem_n17784), .ZN(MEM_stage_inst_dmem_n10476) );
NAND2_X1 MEM_stage_inst_dmem_U16162 ( .A1(EX_pipeline_reg_out_6), .A2(MEM_stage_inst_dmem_n17787), .ZN(MEM_stage_inst_dmem_n17784) );
NAND2_X1 MEM_stage_inst_dmem_U16161 ( .A1(MEM_stage_inst_dmem_ram_2225), .A2(MEM_stage_inst_dmem_n17786), .ZN(MEM_stage_inst_dmem_n17785) );
NAND2_X1 MEM_stage_inst_dmem_U16160 ( .A1(MEM_stage_inst_dmem_n17783), .A2(MEM_stage_inst_dmem_n17782), .ZN(MEM_stage_inst_dmem_n10477) );
NAND2_X1 MEM_stage_inst_dmem_U16159 ( .A1(EX_pipeline_reg_out_7), .A2(MEM_stage_inst_dmem_n17787), .ZN(MEM_stage_inst_dmem_n17782) );
NAND2_X1 MEM_stage_inst_dmem_U16158 ( .A1(MEM_stage_inst_dmem_ram_2226), .A2(MEM_stage_inst_dmem_n17786), .ZN(MEM_stage_inst_dmem_n17783) );
NAND2_X1 MEM_stage_inst_dmem_U16157 ( .A1(MEM_stage_inst_dmem_n17781), .A2(MEM_stage_inst_dmem_n17780), .ZN(MEM_stage_inst_dmem_n10478) );
NAND2_X1 MEM_stage_inst_dmem_U16156 ( .A1(EX_pipeline_reg_out_8), .A2(MEM_stage_inst_dmem_n17787), .ZN(MEM_stage_inst_dmem_n17780) );
NAND2_X1 MEM_stage_inst_dmem_U16155 ( .A1(MEM_stage_inst_dmem_ram_2227), .A2(MEM_stage_inst_dmem_n17786), .ZN(MEM_stage_inst_dmem_n17781) );
NAND2_X1 MEM_stage_inst_dmem_U16154 ( .A1(MEM_stage_inst_dmem_n17779), .A2(MEM_stage_inst_dmem_n17778), .ZN(MEM_stage_inst_dmem_n10479) );
NAND2_X1 MEM_stage_inst_dmem_U16153 ( .A1(EX_pipeline_reg_out_9), .A2(MEM_stage_inst_dmem_n17787), .ZN(MEM_stage_inst_dmem_n17778) );
NAND2_X1 MEM_stage_inst_dmem_U16152 ( .A1(MEM_stage_inst_dmem_ram_2228), .A2(MEM_stage_inst_dmem_n17786), .ZN(MEM_stage_inst_dmem_n17779) );
NAND2_X1 MEM_stage_inst_dmem_U16151 ( .A1(MEM_stage_inst_dmem_n17777), .A2(MEM_stage_inst_dmem_n17776), .ZN(MEM_stage_inst_dmem_n10480) );
NAND2_X1 MEM_stage_inst_dmem_U16150 ( .A1(EX_pipeline_reg_out_10), .A2(MEM_stage_inst_dmem_n17787), .ZN(MEM_stage_inst_dmem_n17776) );
NAND2_X1 MEM_stage_inst_dmem_U16149 ( .A1(MEM_stage_inst_dmem_ram_2229), .A2(MEM_stage_inst_dmem_n17786), .ZN(MEM_stage_inst_dmem_n17777) );
NAND2_X1 MEM_stage_inst_dmem_U16148 ( .A1(MEM_stage_inst_dmem_n17775), .A2(MEM_stage_inst_dmem_n17774), .ZN(MEM_stage_inst_dmem_n10481) );
NAND2_X1 MEM_stage_inst_dmem_U16147 ( .A1(EX_pipeline_reg_out_11), .A2(MEM_stage_inst_dmem_n17787), .ZN(MEM_stage_inst_dmem_n17774) );
NAND2_X1 MEM_stage_inst_dmem_U16146 ( .A1(MEM_stage_inst_dmem_ram_2230), .A2(MEM_stage_inst_dmem_n17786), .ZN(MEM_stage_inst_dmem_n17775) );
NAND2_X1 MEM_stage_inst_dmem_U16145 ( .A1(MEM_stage_inst_dmem_n17773), .A2(MEM_stage_inst_dmem_n17772), .ZN(MEM_stage_inst_dmem_n10482) );
NAND2_X1 MEM_stage_inst_dmem_U16144 ( .A1(EX_pipeline_reg_out_12), .A2(MEM_stage_inst_dmem_n17787), .ZN(MEM_stage_inst_dmem_n17772) );
NAND2_X1 MEM_stage_inst_dmem_U16143 ( .A1(MEM_stage_inst_dmem_ram_2231), .A2(MEM_stage_inst_dmem_n17786), .ZN(MEM_stage_inst_dmem_n17773) );
NAND2_X1 MEM_stage_inst_dmem_U16142 ( .A1(MEM_stage_inst_dmem_n17771), .A2(MEM_stage_inst_dmem_n17770), .ZN(MEM_stage_inst_dmem_n10483) );
NAND2_X1 MEM_stage_inst_dmem_U16141 ( .A1(EX_pipeline_reg_out_13), .A2(MEM_stage_inst_dmem_n17787), .ZN(MEM_stage_inst_dmem_n17770) );
NAND2_X1 MEM_stage_inst_dmem_U16140 ( .A1(MEM_stage_inst_dmem_ram_2232), .A2(MEM_stage_inst_dmem_n17786), .ZN(MEM_stage_inst_dmem_n17771) );
NAND2_X1 MEM_stage_inst_dmem_U16139 ( .A1(MEM_stage_inst_dmem_n17769), .A2(MEM_stage_inst_dmem_n17768), .ZN(MEM_stage_inst_dmem_n10484) );
NAND2_X1 MEM_stage_inst_dmem_U16138 ( .A1(EX_pipeline_reg_out_14), .A2(MEM_stage_inst_dmem_n17787), .ZN(MEM_stage_inst_dmem_n17768) );
NAND2_X1 MEM_stage_inst_dmem_U16137 ( .A1(MEM_stage_inst_dmem_ram_2233), .A2(MEM_stage_inst_dmem_n17786), .ZN(MEM_stage_inst_dmem_n17769) );
NAND2_X1 MEM_stage_inst_dmem_U16136 ( .A1(MEM_stage_inst_dmem_n17767), .A2(MEM_stage_inst_dmem_n17766), .ZN(MEM_stage_inst_dmem_n10485) );
NAND2_X1 MEM_stage_inst_dmem_U16135 ( .A1(EX_pipeline_reg_out_15), .A2(MEM_stage_inst_dmem_n17787), .ZN(MEM_stage_inst_dmem_n17766) );
NAND2_X1 MEM_stage_inst_dmem_U16134 ( .A1(MEM_stage_inst_dmem_ram_2234), .A2(MEM_stage_inst_dmem_n17786), .ZN(MEM_stage_inst_dmem_n17767) );
NAND2_X1 MEM_stage_inst_dmem_U16133 ( .A1(MEM_stage_inst_dmem_n17765), .A2(MEM_stage_inst_dmem_n17764), .ZN(MEM_stage_inst_dmem_n10486) );
NAND2_X1 MEM_stage_inst_dmem_U16132 ( .A1(EX_pipeline_reg_out_16), .A2(MEM_stage_inst_dmem_n17787), .ZN(MEM_stage_inst_dmem_n17764) );
NAND2_X1 MEM_stage_inst_dmem_U16131 ( .A1(MEM_stage_inst_dmem_ram_2235), .A2(MEM_stage_inst_dmem_n17786), .ZN(MEM_stage_inst_dmem_n17765) );
NAND2_X1 MEM_stage_inst_dmem_U16130 ( .A1(MEM_stage_inst_dmem_n17763), .A2(MEM_stage_inst_dmem_n17762), .ZN(MEM_stage_inst_dmem_n10487) );
NAND2_X1 MEM_stage_inst_dmem_U16129 ( .A1(EX_pipeline_reg_out_17), .A2(MEM_stage_inst_dmem_n17787), .ZN(MEM_stage_inst_dmem_n17762) );
NAND2_X1 MEM_stage_inst_dmem_U16128 ( .A1(MEM_stage_inst_dmem_ram_2236), .A2(MEM_stage_inst_dmem_n17786), .ZN(MEM_stage_inst_dmem_n17763) );
NAND2_X1 MEM_stage_inst_dmem_U16127 ( .A1(MEM_stage_inst_dmem_n17761), .A2(MEM_stage_inst_dmem_n17760), .ZN(MEM_stage_inst_dmem_n10488) );
NAND2_X1 MEM_stage_inst_dmem_U16126 ( .A1(EX_pipeline_reg_out_18), .A2(MEM_stage_inst_dmem_n17787), .ZN(MEM_stage_inst_dmem_n17760) );
NAND2_X1 MEM_stage_inst_dmem_U16125 ( .A1(MEM_stage_inst_dmem_ram_2237), .A2(MEM_stage_inst_dmem_n17786), .ZN(MEM_stage_inst_dmem_n17761) );
NAND2_X1 MEM_stage_inst_dmem_U16124 ( .A1(MEM_stage_inst_dmem_n17759), .A2(MEM_stage_inst_dmem_n17758), .ZN(MEM_stage_inst_dmem_n10489) );
NAND2_X1 MEM_stage_inst_dmem_U16123 ( .A1(EX_pipeline_reg_out_19), .A2(MEM_stage_inst_dmem_n17787), .ZN(MEM_stage_inst_dmem_n17758) );
NAND2_X1 MEM_stage_inst_dmem_U16122 ( .A1(MEM_stage_inst_dmem_ram_2238), .A2(MEM_stage_inst_dmem_n17786), .ZN(MEM_stage_inst_dmem_n17759) );
NAND2_X1 MEM_stage_inst_dmem_U16121 ( .A1(MEM_stage_inst_dmem_n17757), .A2(MEM_stage_inst_dmem_n17756), .ZN(MEM_stage_inst_dmem_n10490) );
NAND2_X1 MEM_stage_inst_dmem_U16120 ( .A1(EX_pipeline_reg_out_20), .A2(MEM_stage_inst_dmem_n17787), .ZN(MEM_stage_inst_dmem_n17756) );
INV_X1 MEM_stage_inst_dmem_U16119 ( .A(MEM_stage_inst_dmem_n17786), .ZN(MEM_stage_inst_dmem_n17787) );
NAND2_X1 MEM_stage_inst_dmem_U16118 ( .A1(MEM_stage_inst_dmem_ram_2239), .A2(MEM_stage_inst_dmem_n17786), .ZN(MEM_stage_inst_dmem_n17757) );
NAND2_X1 MEM_stage_inst_dmem_U16117 ( .A1(MEM_stage_inst_dmem_n21074), .A2(MEM_stage_inst_dmem_n18138), .ZN(MEM_stage_inst_dmem_n17786) );
NAND2_X1 MEM_stage_inst_dmem_U16116 ( .A1(MEM_stage_inst_dmem_n17755), .A2(MEM_stage_inst_dmem_n17754), .ZN(MEM_stage_inst_dmem_n10491) );
NAND2_X1 MEM_stage_inst_dmem_U16115 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n17753), .ZN(MEM_stage_inst_dmem_n17754) );
NAND2_X1 MEM_stage_inst_dmem_U16114 ( .A1(MEM_stage_inst_dmem_ram_2240), .A2(MEM_stage_inst_dmem_n17752), .ZN(MEM_stage_inst_dmem_n17755) );
NAND2_X1 MEM_stage_inst_dmem_U16113 ( .A1(MEM_stage_inst_dmem_n17751), .A2(MEM_stage_inst_dmem_n17750), .ZN(MEM_stage_inst_dmem_n10492) );
NAND2_X1 MEM_stage_inst_dmem_U16112 ( .A1(MEM_stage_inst_dmem_n109), .A2(MEM_stage_inst_dmem_n17753), .ZN(MEM_stage_inst_dmem_n17750) );
NAND2_X1 MEM_stage_inst_dmem_U16111 ( .A1(MEM_stage_inst_dmem_ram_2241), .A2(MEM_stage_inst_dmem_n17752), .ZN(MEM_stage_inst_dmem_n17751) );
NAND2_X1 MEM_stage_inst_dmem_U16110 ( .A1(MEM_stage_inst_dmem_n17749), .A2(MEM_stage_inst_dmem_n17748), .ZN(MEM_stage_inst_dmem_n10493) );
NAND2_X1 MEM_stage_inst_dmem_U16109 ( .A1(MEM_stage_inst_dmem_n18027), .A2(MEM_stage_inst_dmem_n17753), .ZN(MEM_stage_inst_dmem_n17748) );
NAND2_X1 MEM_stage_inst_dmem_U16108 ( .A1(MEM_stage_inst_dmem_ram_2242), .A2(MEM_stage_inst_dmem_n17752), .ZN(MEM_stage_inst_dmem_n17749) );
NAND2_X1 MEM_stage_inst_dmem_U16107 ( .A1(MEM_stage_inst_dmem_n17747), .A2(MEM_stage_inst_dmem_n17746), .ZN(MEM_stage_inst_dmem_n10494) );
NAND2_X1 MEM_stage_inst_dmem_U16106 ( .A1(MEM_stage_inst_dmem_n13064), .A2(MEM_stage_inst_dmem_n17753), .ZN(MEM_stage_inst_dmem_n17746) );
NAND2_X1 MEM_stage_inst_dmem_U16105 ( .A1(MEM_stage_inst_dmem_ram_2243), .A2(MEM_stage_inst_dmem_n17752), .ZN(MEM_stage_inst_dmem_n17747) );
NAND2_X1 MEM_stage_inst_dmem_U16104 ( .A1(MEM_stage_inst_dmem_n17745), .A2(MEM_stage_inst_dmem_n17744), .ZN(MEM_stage_inst_dmem_n10495) );
NAND2_X1 MEM_stage_inst_dmem_U16103 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n17753), .ZN(MEM_stage_inst_dmem_n17744) );
NAND2_X1 MEM_stage_inst_dmem_U16102 ( .A1(MEM_stage_inst_dmem_ram_2244), .A2(MEM_stage_inst_dmem_n17752), .ZN(MEM_stage_inst_dmem_n17745) );
NAND2_X1 MEM_stage_inst_dmem_U16101 ( .A1(MEM_stage_inst_dmem_n17743), .A2(MEM_stage_inst_dmem_n17742), .ZN(MEM_stage_inst_dmem_n10496) );
NAND2_X1 MEM_stage_inst_dmem_U16100 ( .A1(MEM_stage_inst_dmem_n13059), .A2(MEM_stage_inst_dmem_n17753), .ZN(MEM_stage_inst_dmem_n17742) );
NAND2_X1 MEM_stage_inst_dmem_U16099 ( .A1(MEM_stage_inst_dmem_ram_2245), .A2(MEM_stage_inst_dmem_n17752), .ZN(MEM_stage_inst_dmem_n17743) );
NAND2_X1 MEM_stage_inst_dmem_U16098 ( .A1(MEM_stage_inst_dmem_n17741), .A2(MEM_stage_inst_dmem_n17740), .ZN(MEM_stage_inst_dmem_n10497) );
NAND2_X1 MEM_stage_inst_dmem_U16097 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n17753), .ZN(MEM_stage_inst_dmem_n17740) );
NAND2_X1 MEM_stage_inst_dmem_U16096 ( .A1(MEM_stage_inst_dmem_ram_2246), .A2(MEM_stage_inst_dmem_n17752), .ZN(MEM_stage_inst_dmem_n17741) );
NAND2_X1 MEM_stage_inst_dmem_U16095 ( .A1(MEM_stage_inst_dmem_n17739), .A2(MEM_stage_inst_dmem_n17738), .ZN(MEM_stage_inst_dmem_n10498) );
NAND2_X1 MEM_stage_inst_dmem_U16094 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n17753), .ZN(MEM_stage_inst_dmem_n17738) );
NAND2_X1 MEM_stage_inst_dmem_U16093 ( .A1(MEM_stage_inst_dmem_ram_2247), .A2(MEM_stage_inst_dmem_n17752), .ZN(MEM_stage_inst_dmem_n17739) );
NAND2_X1 MEM_stage_inst_dmem_U16092 ( .A1(MEM_stage_inst_dmem_n17737), .A2(MEM_stage_inst_dmem_n17736), .ZN(MEM_stage_inst_dmem_n10499) );
NAND2_X1 MEM_stage_inst_dmem_U16091 ( .A1(MEM_stage_inst_dmem_n18013), .A2(MEM_stage_inst_dmem_n17753), .ZN(MEM_stage_inst_dmem_n17736) );
NAND2_X1 MEM_stage_inst_dmem_U16090 ( .A1(MEM_stage_inst_dmem_ram_2248), .A2(MEM_stage_inst_dmem_n17752), .ZN(MEM_stage_inst_dmem_n17737) );
NAND2_X1 MEM_stage_inst_dmem_U16089 ( .A1(MEM_stage_inst_dmem_n17735), .A2(MEM_stage_inst_dmem_n17734), .ZN(MEM_stage_inst_dmem_n10500) );
NAND2_X1 MEM_stage_inst_dmem_U16088 ( .A1(MEM_stage_inst_dmem_n96), .A2(MEM_stage_inst_dmem_n17753), .ZN(MEM_stage_inst_dmem_n17734) );
NAND2_X1 MEM_stage_inst_dmem_U16087 ( .A1(MEM_stage_inst_dmem_ram_2249), .A2(MEM_stage_inst_dmem_n17752), .ZN(MEM_stage_inst_dmem_n17735) );
NAND2_X1 MEM_stage_inst_dmem_U16086 ( .A1(MEM_stage_inst_dmem_n17733), .A2(MEM_stage_inst_dmem_n17732), .ZN(MEM_stage_inst_dmem_n10501) );
NAND2_X1 MEM_stage_inst_dmem_U16085 ( .A1(MEM_stage_inst_dmem_n18007), .A2(MEM_stage_inst_dmem_n17753), .ZN(MEM_stage_inst_dmem_n17732) );
NAND2_X1 MEM_stage_inst_dmem_U16084 ( .A1(MEM_stage_inst_dmem_ram_2250), .A2(MEM_stage_inst_dmem_n17752), .ZN(MEM_stage_inst_dmem_n17733) );
NAND2_X1 MEM_stage_inst_dmem_U16083 ( .A1(MEM_stage_inst_dmem_n17731), .A2(MEM_stage_inst_dmem_n17730), .ZN(MEM_stage_inst_dmem_n10502) );
NAND2_X1 MEM_stage_inst_dmem_U16082 ( .A1(MEM_stage_inst_dmem_n18004), .A2(MEM_stage_inst_dmem_n17753), .ZN(MEM_stage_inst_dmem_n17730) );
NAND2_X1 MEM_stage_inst_dmem_U16081 ( .A1(MEM_stage_inst_dmem_ram_2251), .A2(MEM_stage_inst_dmem_n17752), .ZN(MEM_stage_inst_dmem_n17731) );
NAND2_X1 MEM_stage_inst_dmem_U16080 ( .A1(MEM_stage_inst_dmem_n17729), .A2(MEM_stage_inst_dmem_n17728), .ZN(MEM_stage_inst_dmem_n10503) );
NAND2_X1 MEM_stage_inst_dmem_U16079 ( .A1(MEM_stage_inst_dmem_n18001), .A2(MEM_stage_inst_dmem_n17753), .ZN(MEM_stage_inst_dmem_n17728) );
NAND2_X1 MEM_stage_inst_dmem_U16078 ( .A1(MEM_stage_inst_dmem_ram_2252), .A2(MEM_stage_inst_dmem_n17752), .ZN(MEM_stage_inst_dmem_n17729) );
NAND2_X1 MEM_stage_inst_dmem_U16077 ( .A1(MEM_stage_inst_dmem_n17727), .A2(MEM_stage_inst_dmem_n17726), .ZN(MEM_stage_inst_dmem_n10504) );
NAND2_X1 MEM_stage_inst_dmem_U16076 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n17753), .ZN(MEM_stage_inst_dmem_n17726) );
NAND2_X1 MEM_stage_inst_dmem_U16075 ( .A1(MEM_stage_inst_dmem_ram_2253), .A2(MEM_stage_inst_dmem_n17752), .ZN(MEM_stage_inst_dmem_n17727) );
NAND2_X1 MEM_stage_inst_dmem_U16074 ( .A1(MEM_stage_inst_dmem_n17725), .A2(MEM_stage_inst_dmem_n17724), .ZN(MEM_stage_inst_dmem_n10505) );
NAND2_X1 MEM_stage_inst_dmem_U16073 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n17753), .ZN(MEM_stage_inst_dmem_n17724) );
NAND2_X1 MEM_stage_inst_dmem_U16072 ( .A1(MEM_stage_inst_dmem_ram_2254), .A2(MEM_stage_inst_dmem_n17752), .ZN(MEM_stage_inst_dmem_n17725) );
NAND2_X1 MEM_stage_inst_dmem_U16071 ( .A1(MEM_stage_inst_dmem_n17723), .A2(MEM_stage_inst_dmem_n17722), .ZN(MEM_stage_inst_dmem_n10506) );
NAND2_X1 MEM_stage_inst_dmem_U16070 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n17753), .ZN(MEM_stage_inst_dmem_n17722) );
INV_X1 MEM_stage_inst_dmem_U16069 ( .A(MEM_stage_inst_dmem_n17752), .ZN(MEM_stage_inst_dmem_n17753) );
NAND2_X1 MEM_stage_inst_dmem_U16068 ( .A1(MEM_stage_inst_dmem_ram_2255), .A2(MEM_stage_inst_dmem_n17752), .ZN(MEM_stage_inst_dmem_n17723) );
NAND2_X1 MEM_stage_inst_dmem_U16067 ( .A1(MEM_stage_inst_dmem_n21039), .A2(MEM_stage_inst_dmem_n18138), .ZN(MEM_stage_inst_dmem_n17752) );
NAND2_X1 MEM_stage_inst_dmem_U16066 ( .A1(MEM_stage_inst_dmem_n17721), .A2(MEM_stage_inst_dmem_n17720), .ZN(MEM_stage_inst_dmem_n10507) );
NAND2_X1 MEM_stage_inst_dmem_U16065 ( .A1(EX_pipeline_reg_out_5), .A2(MEM_stage_inst_dmem_n17719), .ZN(MEM_stage_inst_dmem_n17720) );
NAND2_X1 MEM_stage_inst_dmem_U16064 ( .A1(MEM_stage_inst_dmem_ram_2256), .A2(MEM_stage_inst_dmem_n17718), .ZN(MEM_stage_inst_dmem_n17721) );
NAND2_X1 MEM_stage_inst_dmem_U16063 ( .A1(MEM_stage_inst_dmem_n17717), .A2(MEM_stage_inst_dmem_n17716), .ZN(MEM_stage_inst_dmem_n10508) );
NAND2_X1 MEM_stage_inst_dmem_U16062 ( .A1(EX_pipeline_reg_out_6), .A2(MEM_stage_inst_dmem_n17719), .ZN(MEM_stage_inst_dmem_n17716) );
NAND2_X1 MEM_stage_inst_dmem_U16061 ( .A1(MEM_stage_inst_dmem_ram_2257), .A2(MEM_stage_inst_dmem_n17718), .ZN(MEM_stage_inst_dmem_n17717) );
NAND2_X1 MEM_stage_inst_dmem_U16060 ( .A1(MEM_stage_inst_dmem_n17715), .A2(MEM_stage_inst_dmem_n17714), .ZN(MEM_stage_inst_dmem_n10509) );
NAND2_X1 MEM_stage_inst_dmem_U16059 ( .A1(EX_pipeline_reg_out_7), .A2(MEM_stage_inst_dmem_n17719), .ZN(MEM_stage_inst_dmem_n17714) );
NAND2_X1 MEM_stage_inst_dmem_U16058 ( .A1(MEM_stage_inst_dmem_ram_2258), .A2(MEM_stage_inst_dmem_n17718), .ZN(MEM_stage_inst_dmem_n17715) );
NAND2_X1 MEM_stage_inst_dmem_U16057 ( .A1(MEM_stage_inst_dmem_n17713), .A2(MEM_stage_inst_dmem_n17712), .ZN(MEM_stage_inst_dmem_n10510) );
NAND2_X1 MEM_stage_inst_dmem_U16056 ( .A1(EX_pipeline_reg_out_8), .A2(MEM_stage_inst_dmem_n17719), .ZN(MEM_stage_inst_dmem_n17712) );
NAND2_X1 MEM_stage_inst_dmem_U16055 ( .A1(MEM_stage_inst_dmem_ram_2259), .A2(MEM_stage_inst_dmem_n17718), .ZN(MEM_stage_inst_dmem_n17713) );
NAND2_X1 MEM_stage_inst_dmem_U16054 ( .A1(MEM_stage_inst_dmem_n17711), .A2(MEM_stage_inst_dmem_n17710), .ZN(MEM_stage_inst_dmem_n10511) );
NAND2_X1 MEM_stage_inst_dmem_U16053 ( .A1(EX_pipeline_reg_out_9), .A2(MEM_stage_inst_dmem_n17719), .ZN(MEM_stage_inst_dmem_n17710) );
NAND2_X1 MEM_stage_inst_dmem_U16052 ( .A1(MEM_stage_inst_dmem_ram_2260), .A2(MEM_stage_inst_dmem_n17718), .ZN(MEM_stage_inst_dmem_n17711) );
NAND2_X1 MEM_stage_inst_dmem_U16051 ( .A1(MEM_stage_inst_dmem_n17709), .A2(MEM_stage_inst_dmem_n17708), .ZN(MEM_stage_inst_dmem_n10512) );
NAND2_X1 MEM_stage_inst_dmem_U16050 ( .A1(EX_pipeline_reg_out_10), .A2(MEM_stage_inst_dmem_n17719), .ZN(MEM_stage_inst_dmem_n17708) );
NAND2_X1 MEM_stage_inst_dmem_U16049 ( .A1(MEM_stage_inst_dmem_ram_2261), .A2(MEM_stage_inst_dmem_n17718), .ZN(MEM_stage_inst_dmem_n17709) );
NAND2_X1 MEM_stage_inst_dmem_U16048 ( .A1(MEM_stage_inst_dmem_n17707), .A2(MEM_stage_inst_dmem_n17706), .ZN(MEM_stage_inst_dmem_n10513) );
NAND2_X1 MEM_stage_inst_dmem_U16047 ( .A1(EX_pipeline_reg_out_11), .A2(MEM_stage_inst_dmem_n17719), .ZN(MEM_stage_inst_dmem_n17706) );
NAND2_X1 MEM_stage_inst_dmem_U16046 ( .A1(MEM_stage_inst_dmem_ram_2262), .A2(MEM_stage_inst_dmem_n17718), .ZN(MEM_stage_inst_dmem_n17707) );
NAND2_X1 MEM_stage_inst_dmem_U16045 ( .A1(MEM_stage_inst_dmem_n17705), .A2(MEM_stage_inst_dmem_n17704), .ZN(MEM_stage_inst_dmem_n10514) );
NAND2_X1 MEM_stage_inst_dmem_U16044 ( .A1(EX_pipeline_reg_out_12), .A2(MEM_stage_inst_dmem_n17719), .ZN(MEM_stage_inst_dmem_n17704) );
NAND2_X1 MEM_stage_inst_dmem_U16043 ( .A1(MEM_stage_inst_dmem_ram_2263), .A2(MEM_stage_inst_dmem_n17718), .ZN(MEM_stage_inst_dmem_n17705) );
NAND2_X1 MEM_stage_inst_dmem_U16042 ( .A1(MEM_stage_inst_dmem_n17703), .A2(MEM_stage_inst_dmem_n17702), .ZN(MEM_stage_inst_dmem_n10515) );
NAND2_X1 MEM_stage_inst_dmem_U16041 ( .A1(EX_pipeline_reg_out_13), .A2(MEM_stage_inst_dmem_n17719), .ZN(MEM_stage_inst_dmem_n17702) );
NAND2_X1 MEM_stage_inst_dmem_U16040 ( .A1(MEM_stage_inst_dmem_ram_2264), .A2(MEM_stage_inst_dmem_n17718), .ZN(MEM_stage_inst_dmem_n17703) );
NAND2_X1 MEM_stage_inst_dmem_U16039 ( .A1(MEM_stage_inst_dmem_n17701), .A2(MEM_stage_inst_dmem_n17700), .ZN(MEM_stage_inst_dmem_n10516) );
NAND2_X1 MEM_stage_inst_dmem_U16038 ( .A1(EX_pipeline_reg_out_14), .A2(MEM_stage_inst_dmem_n17719), .ZN(MEM_stage_inst_dmem_n17700) );
NAND2_X1 MEM_stage_inst_dmem_U16037 ( .A1(MEM_stage_inst_dmem_ram_2265), .A2(MEM_stage_inst_dmem_n17718), .ZN(MEM_stage_inst_dmem_n17701) );
NAND2_X1 MEM_stage_inst_dmem_U16036 ( .A1(MEM_stage_inst_dmem_n17699), .A2(MEM_stage_inst_dmem_n17698), .ZN(MEM_stage_inst_dmem_n10517) );
NAND2_X1 MEM_stage_inst_dmem_U16035 ( .A1(EX_pipeline_reg_out_15), .A2(MEM_stage_inst_dmem_n17719), .ZN(MEM_stage_inst_dmem_n17698) );
NAND2_X1 MEM_stage_inst_dmem_U16034 ( .A1(MEM_stage_inst_dmem_ram_2266), .A2(MEM_stage_inst_dmem_n17718), .ZN(MEM_stage_inst_dmem_n17699) );
NAND2_X1 MEM_stage_inst_dmem_U16033 ( .A1(MEM_stage_inst_dmem_n17697), .A2(MEM_stage_inst_dmem_n17696), .ZN(MEM_stage_inst_dmem_n10518) );
NAND2_X1 MEM_stage_inst_dmem_U16032 ( .A1(EX_pipeline_reg_out_16), .A2(MEM_stage_inst_dmem_n17719), .ZN(MEM_stage_inst_dmem_n17696) );
NAND2_X1 MEM_stage_inst_dmem_U16031 ( .A1(MEM_stage_inst_dmem_ram_2267), .A2(MEM_stage_inst_dmem_n17718), .ZN(MEM_stage_inst_dmem_n17697) );
NAND2_X1 MEM_stage_inst_dmem_U16030 ( .A1(MEM_stage_inst_dmem_n17695), .A2(MEM_stage_inst_dmem_n17694), .ZN(MEM_stage_inst_dmem_n10519) );
NAND2_X1 MEM_stage_inst_dmem_U16029 ( .A1(EX_pipeline_reg_out_17), .A2(MEM_stage_inst_dmem_n17719), .ZN(MEM_stage_inst_dmem_n17694) );
NAND2_X1 MEM_stage_inst_dmem_U16028 ( .A1(MEM_stage_inst_dmem_ram_2268), .A2(MEM_stage_inst_dmem_n17718), .ZN(MEM_stage_inst_dmem_n17695) );
NAND2_X1 MEM_stage_inst_dmem_U16027 ( .A1(MEM_stage_inst_dmem_n17693), .A2(MEM_stage_inst_dmem_n17692), .ZN(MEM_stage_inst_dmem_n10520) );
NAND2_X1 MEM_stage_inst_dmem_U16026 ( .A1(EX_pipeline_reg_out_18), .A2(MEM_stage_inst_dmem_n17719), .ZN(MEM_stage_inst_dmem_n17692) );
NAND2_X1 MEM_stage_inst_dmem_U16025 ( .A1(MEM_stage_inst_dmem_ram_2269), .A2(MEM_stage_inst_dmem_n17718), .ZN(MEM_stage_inst_dmem_n17693) );
NAND2_X1 MEM_stage_inst_dmem_U16024 ( .A1(MEM_stage_inst_dmem_n17691), .A2(MEM_stage_inst_dmem_n17690), .ZN(MEM_stage_inst_dmem_n10521) );
NAND2_X1 MEM_stage_inst_dmem_U16023 ( .A1(EX_pipeline_reg_out_19), .A2(MEM_stage_inst_dmem_n17719), .ZN(MEM_stage_inst_dmem_n17690) );
NAND2_X1 MEM_stage_inst_dmem_U16022 ( .A1(MEM_stage_inst_dmem_ram_2270), .A2(MEM_stage_inst_dmem_n17718), .ZN(MEM_stage_inst_dmem_n17691) );
NAND2_X1 MEM_stage_inst_dmem_U16021 ( .A1(MEM_stage_inst_dmem_n17689), .A2(MEM_stage_inst_dmem_n17688), .ZN(MEM_stage_inst_dmem_n10522) );
NAND2_X1 MEM_stage_inst_dmem_U16020 ( .A1(EX_pipeline_reg_out_20), .A2(MEM_stage_inst_dmem_n17719), .ZN(MEM_stage_inst_dmem_n17688) );
INV_X1 MEM_stage_inst_dmem_U16019 ( .A(MEM_stage_inst_dmem_n17718), .ZN(MEM_stage_inst_dmem_n17719) );
NAND2_X1 MEM_stage_inst_dmem_U16018 ( .A1(MEM_stage_inst_dmem_ram_2271), .A2(MEM_stage_inst_dmem_n17718), .ZN(MEM_stage_inst_dmem_n17689) );
NAND2_X1 MEM_stage_inst_dmem_U16017 ( .A1(MEM_stage_inst_dmem_n21004), .A2(MEM_stage_inst_dmem_n18138), .ZN(MEM_stage_inst_dmem_n17718) );
NAND2_X1 MEM_stage_inst_dmem_U16016 ( .A1(MEM_stage_inst_dmem_n17687), .A2(MEM_stage_inst_dmem_n17686), .ZN(MEM_stage_inst_dmem_n10523) );
NAND2_X1 MEM_stage_inst_dmem_U16015 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n17685), .ZN(MEM_stage_inst_dmem_n17686) );
NAND2_X1 MEM_stage_inst_dmem_U16014 ( .A1(MEM_stage_inst_dmem_ram_2272), .A2(MEM_stage_inst_dmem_n17684), .ZN(MEM_stage_inst_dmem_n17687) );
NAND2_X1 MEM_stage_inst_dmem_U16013 ( .A1(MEM_stage_inst_dmem_n17683), .A2(MEM_stage_inst_dmem_n17682), .ZN(MEM_stage_inst_dmem_n10524) );
NAND2_X1 MEM_stage_inst_dmem_U16012 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n17685), .ZN(MEM_stage_inst_dmem_n17682) );
NAND2_X1 MEM_stage_inst_dmem_U16011 ( .A1(MEM_stage_inst_dmem_ram_2273), .A2(MEM_stage_inst_dmem_n17684), .ZN(MEM_stage_inst_dmem_n17683) );
NAND2_X1 MEM_stage_inst_dmem_U16010 ( .A1(MEM_stage_inst_dmem_n17681), .A2(MEM_stage_inst_dmem_n17680), .ZN(MEM_stage_inst_dmem_n10525) );
NAND2_X1 MEM_stage_inst_dmem_U16009 ( .A1(MEM_stage_inst_dmem_n18027), .A2(MEM_stage_inst_dmem_n17685), .ZN(MEM_stage_inst_dmem_n17680) );
NAND2_X1 MEM_stage_inst_dmem_U16008 ( .A1(MEM_stage_inst_dmem_ram_2274), .A2(MEM_stage_inst_dmem_n17684), .ZN(MEM_stage_inst_dmem_n17681) );
NAND2_X1 MEM_stage_inst_dmem_U16007 ( .A1(MEM_stage_inst_dmem_n17679), .A2(MEM_stage_inst_dmem_n17678), .ZN(MEM_stage_inst_dmem_n10526) );
NAND2_X1 MEM_stage_inst_dmem_U16006 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n17685), .ZN(MEM_stage_inst_dmem_n17678) );
NAND2_X1 MEM_stage_inst_dmem_U16005 ( .A1(MEM_stage_inst_dmem_ram_2275), .A2(MEM_stage_inst_dmem_n17684), .ZN(MEM_stage_inst_dmem_n17679) );
NAND2_X1 MEM_stage_inst_dmem_U16004 ( .A1(MEM_stage_inst_dmem_n17677), .A2(MEM_stage_inst_dmem_n17676), .ZN(MEM_stage_inst_dmem_n10527) );
NAND2_X1 MEM_stage_inst_dmem_U16003 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n17685), .ZN(MEM_stage_inst_dmem_n17676) );
NAND2_X1 MEM_stage_inst_dmem_U16002 ( .A1(MEM_stage_inst_dmem_ram_2276), .A2(MEM_stage_inst_dmem_n17684), .ZN(MEM_stage_inst_dmem_n17677) );
NAND2_X1 MEM_stage_inst_dmem_U16001 ( .A1(MEM_stage_inst_dmem_n17675), .A2(MEM_stage_inst_dmem_n17674), .ZN(MEM_stage_inst_dmem_n10528) );
NAND2_X1 MEM_stage_inst_dmem_U16000 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n17685), .ZN(MEM_stage_inst_dmem_n17674) );
NAND2_X1 MEM_stage_inst_dmem_U15999 ( .A1(MEM_stage_inst_dmem_ram_2277), .A2(MEM_stage_inst_dmem_n17684), .ZN(MEM_stage_inst_dmem_n17675) );
NAND2_X1 MEM_stage_inst_dmem_U15998 ( .A1(MEM_stage_inst_dmem_n17673), .A2(MEM_stage_inst_dmem_n17672), .ZN(MEM_stage_inst_dmem_n10529) );
NAND2_X1 MEM_stage_inst_dmem_U15997 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n17685), .ZN(MEM_stage_inst_dmem_n17672) );
NAND2_X1 MEM_stage_inst_dmem_U15996 ( .A1(MEM_stage_inst_dmem_ram_2278), .A2(MEM_stage_inst_dmem_n17684), .ZN(MEM_stage_inst_dmem_n17673) );
NAND2_X1 MEM_stage_inst_dmem_U15995 ( .A1(MEM_stage_inst_dmem_n17671), .A2(MEM_stage_inst_dmem_n17670), .ZN(MEM_stage_inst_dmem_n10530) );
NAND2_X1 MEM_stage_inst_dmem_U15994 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n17685), .ZN(MEM_stage_inst_dmem_n17670) );
NAND2_X1 MEM_stage_inst_dmem_U15993 ( .A1(MEM_stage_inst_dmem_ram_2279), .A2(MEM_stage_inst_dmem_n17684), .ZN(MEM_stage_inst_dmem_n17671) );
NAND2_X1 MEM_stage_inst_dmem_U15992 ( .A1(MEM_stage_inst_dmem_n17669), .A2(MEM_stage_inst_dmem_n17668), .ZN(MEM_stage_inst_dmem_n10531) );
NAND2_X1 MEM_stage_inst_dmem_U15991 ( .A1(MEM_stage_inst_dmem_n18013), .A2(MEM_stage_inst_dmem_n17685), .ZN(MEM_stage_inst_dmem_n17668) );
NAND2_X1 MEM_stage_inst_dmem_U15990 ( .A1(MEM_stage_inst_dmem_ram_2280), .A2(MEM_stage_inst_dmem_n17684), .ZN(MEM_stage_inst_dmem_n17669) );
NAND2_X1 MEM_stage_inst_dmem_U15989 ( .A1(MEM_stage_inst_dmem_n17667), .A2(MEM_stage_inst_dmem_n17666), .ZN(MEM_stage_inst_dmem_n10532) );
NAND2_X1 MEM_stage_inst_dmem_U15988 ( .A1(MEM_stage_inst_dmem_n96), .A2(MEM_stage_inst_dmem_n17685), .ZN(MEM_stage_inst_dmem_n17666) );
NAND2_X1 MEM_stage_inst_dmem_U15987 ( .A1(MEM_stage_inst_dmem_ram_2281), .A2(MEM_stage_inst_dmem_n17684), .ZN(MEM_stage_inst_dmem_n17667) );
NAND2_X1 MEM_stage_inst_dmem_U15986 ( .A1(MEM_stage_inst_dmem_n17665), .A2(MEM_stage_inst_dmem_n17664), .ZN(MEM_stage_inst_dmem_n10533) );
NAND2_X1 MEM_stage_inst_dmem_U15985 ( .A1(MEM_stage_inst_dmem_n18007), .A2(MEM_stage_inst_dmem_n17685), .ZN(MEM_stage_inst_dmem_n17664) );
NAND2_X1 MEM_stage_inst_dmem_U15984 ( .A1(MEM_stage_inst_dmem_ram_2282), .A2(MEM_stage_inst_dmem_n17684), .ZN(MEM_stage_inst_dmem_n17665) );
NAND2_X1 MEM_stage_inst_dmem_U15983 ( .A1(MEM_stage_inst_dmem_n17663), .A2(MEM_stage_inst_dmem_n17662), .ZN(MEM_stage_inst_dmem_n10534) );
NAND2_X1 MEM_stage_inst_dmem_U15982 ( .A1(MEM_stage_inst_dmem_n18004), .A2(MEM_stage_inst_dmem_n17685), .ZN(MEM_stage_inst_dmem_n17662) );
NAND2_X1 MEM_stage_inst_dmem_U15981 ( .A1(MEM_stage_inst_dmem_ram_2283), .A2(MEM_stage_inst_dmem_n17684), .ZN(MEM_stage_inst_dmem_n17663) );
NAND2_X1 MEM_stage_inst_dmem_U15980 ( .A1(MEM_stage_inst_dmem_n17661), .A2(MEM_stage_inst_dmem_n17660), .ZN(MEM_stage_inst_dmem_n10535) );
NAND2_X1 MEM_stage_inst_dmem_U15979 ( .A1(MEM_stage_inst_dmem_n18001), .A2(MEM_stage_inst_dmem_n17685), .ZN(MEM_stage_inst_dmem_n17660) );
NAND2_X1 MEM_stage_inst_dmem_U15978 ( .A1(MEM_stage_inst_dmem_ram_2284), .A2(MEM_stage_inst_dmem_n17684), .ZN(MEM_stage_inst_dmem_n17661) );
NAND2_X1 MEM_stage_inst_dmem_U15977 ( .A1(MEM_stage_inst_dmem_n17659), .A2(MEM_stage_inst_dmem_n17658), .ZN(MEM_stage_inst_dmem_n10536) );
NAND2_X1 MEM_stage_inst_dmem_U15976 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n17685), .ZN(MEM_stage_inst_dmem_n17658) );
NAND2_X1 MEM_stage_inst_dmem_U15975 ( .A1(MEM_stage_inst_dmem_ram_2285), .A2(MEM_stage_inst_dmem_n17684), .ZN(MEM_stage_inst_dmem_n17659) );
NAND2_X1 MEM_stage_inst_dmem_U15974 ( .A1(MEM_stage_inst_dmem_n17657), .A2(MEM_stage_inst_dmem_n17656), .ZN(MEM_stage_inst_dmem_n10537) );
NAND2_X1 MEM_stage_inst_dmem_U15973 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n17685), .ZN(MEM_stage_inst_dmem_n17656) );
NAND2_X1 MEM_stage_inst_dmem_U15972 ( .A1(MEM_stage_inst_dmem_ram_2286), .A2(MEM_stage_inst_dmem_n17684), .ZN(MEM_stage_inst_dmem_n17657) );
NAND2_X1 MEM_stage_inst_dmem_U15971 ( .A1(MEM_stage_inst_dmem_n17655), .A2(MEM_stage_inst_dmem_n17654), .ZN(MEM_stage_inst_dmem_n10538) );
NAND2_X1 MEM_stage_inst_dmem_U15970 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n17685), .ZN(MEM_stage_inst_dmem_n17654) );
INV_X1 MEM_stage_inst_dmem_U15969 ( .A(MEM_stage_inst_dmem_n17684), .ZN(MEM_stage_inst_dmem_n17685) );
NAND2_X1 MEM_stage_inst_dmem_U15968 ( .A1(MEM_stage_inst_dmem_ram_2287), .A2(MEM_stage_inst_dmem_n17684), .ZN(MEM_stage_inst_dmem_n17655) );
NAND2_X1 MEM_stage_inst_dmem_U15967 ( .A1(MEM_stage_inst_dmem_n20969), .A2(MEM_stage_inst_dmem_n18138), .ZN(MEM_stage_inst_dmem_n17684) );
NAND2_X1 MEM_stage_inst_dmem_U15966 ( .A1(MEM_stage_inst_dmem_n17653), .A2(MEM_stage_inst_dmem_n17652), .ZN(MEM_stage_inst_dmem_n10539) );
NAND2_X1 MEM_stage_inst_dmem_U15965 ( .A1(EX_pipeline_reg_out_5), .A2(MEM_stage_inst_dmem_n17651), .ZN(MEM_stage_inst_dmem_n17652) );
NAND2_X1 MEM_stage_inst_dmem_U15964 ( .A1(MEM_stage_inst_dmem_ram_2288), .A2(MEM_stage_inst_dmem_n17650), .ZN(MEM_stage_inst_dmem_n17653) );
NAND2_X1 MEM_stage_inst_dmem_U15963 ( .A1(MEM_stage_inst_dmem_n17649), .A2(MEM_stage_inst_dmem_n17648), .ZN(MEM_stage_inst_dmem_n10540) );
NAND2_X1 MEM_stage_inst_dmem_U15962 ( .A1(EX_pipeline_reg_out_6), .A2(MEM_stage_inst_dmem_n17651), .ZN(MEM_stage_inst_dmem_n17648) );
NAND2_X1 MEM_stage_inst_dmem_U15961 ( .A1(MEM_stage_inst_dmem_ram_2289), .A2(MEM_stage_inst_dmem_n17650), .ZN(MEM_stage_inst_dmem_n17649) );
NAND2_X1 MEM_stage_inst_dmem_U15960 ( .A1(MEM_stage_inst_dmem_n17647), .A2(MEM_stage_inst_dmem_n17646), .ZN(MEM_stage_inst_dmem_n10541) );
NAND2_X1 MEM_stage_inst_dmem_U15959 ( .A1(EX_pipeline_reg_out_7), .A2(MEM_stage_inst_dmem_n17651), .ZN(MEM_stage_inst_dmem_n17646) );
NAND2_X1 MEM_stage_inst_dmem_U15958 ( .A1(MEM_stage_inst_dmem_ram_2290), .A2(MEM_stage_inst_dmem_n17650), .ZN(MEM_stage_inst_dmem_n17647) );
NAND2_X1 MEM_stage_inst_dmem_U15957 ( .A1(MEM_stage_inst_dmem_n17645), .A2(MEM_stage_inst_dmem_n17644), .ZN(MEM_stage_inst_dmem_n10542) );
NAND2_X1 MEM_stage_inst_dmem_U15956 ( .A1(EX_pipeline_reg_out_8), .A2(MEM_stage_inst_dmem_n17651), .ZN(MEM_stage_inst_dmem_n17644) );
NAND2_X1 MEM_stage_inst_dmem_U15955 ( .A1(MEM_stage_inst_dmem_ram_2291), .A2(MEM_stage_inst_dmem_n17650), .ZN(MEM_stage_inst_dmem_n17645) );
NAND2_X1 MEM_stage_inst_dmem_U15954 ( .A1(MEM_stage_inst_dmem_n17643), .A2(MEM_stage_inst_dmem_n17642), .ZN(MEM_stage_inst_dmem_n10543) );
NAND2_X1 MEM_stage_inst_dmem_U15953 ( .A1(EX_pipeline_reg_out_9), .A2(MEM_stage_inst_dmem_n17651), .ZN(MEM_stage_inst_dmem_n17642) );
NAND2_X1 MEM_stage_inst_dmem_U15952 ( .A1(MEM_stage_inst_dmem_ram_2292), .A2(MEM_stage_inst_dmem_n17650), .ZN(MEM_stage_inst_dmem_n17643) );
NAND2_X1 MEM_stage_inst_dmem_U15951 ( .A1(MEM_stage_inst_dmem_n17641), .A2(MEM_stage_inst_dmem_n17640), .ZN(MEM_stage_inst_dmem_n10544) );
NAND2_X1 MEM_stage_inst_dmem_U15950 ( .A1(EX_pipeline_reg_out_10), .A2(MEM_stage_inst_dmem_n17651), .ZN(MEM_stage_inst_dmem_n17640) );
NAND2_X1 MEM_stage_inst_dmem_U15949 ( .A1(MEM_stage_inst_dmem_ram_2293), .A2(MEM_stage_inst_dmem_n17650), .ZN(MEM_stage_inst_dmem_n17641) );
NAND2_X1 MEM_stage_inst_dmem_U15948 ( .A1(MEM_stage_inst_dmem_n17639), .A2(MEM_stage_inst_dmem_n17638), .ZN(MEM_stage_inst_dmem_n10545) );
NAND2_X1 MEM_stage_inst_dmem_U15947 ( .A1(EX_pipeline_reg_out_11), .A2(MEM_stage_inst_dmem_n17651), .ZN(MEM_stage_inst_dmem_n17638) );
NAND2_X1 MEM_stage_inst_dmem_U15946 ( .A1(MEM_stage_inst_dmem_ram_2294), .A2(MEM_stage_inst_dmem_n17650), .ZN(MEM_stage_inst_dmem_n17639) );
NAND2_X1 MEM_stage_inst_dmem_U15945 ( .A1(MEM_stage_inst_dmem_n17637), .A2(MEM_stage_inst_dmem_n17636), .ZN(MEM_stage_inst_dmem_n10546) );
NAND2_X1 MEM_stage_inst_dmem_U15944 ( .A1(EX_pipeline_reg_out_12), .A2(MEM_stage_inst_dmem_n17651), .ZN(MEM_stage_inst_dmem_n17636) );
NAND2_X1 MEM_stage_inst_dmem_U15943 ( .A1(MEM_stage_inst_dmem_ram_2295), .A2(MEM_stage_inst_dmem_n17650), .ZN(MEM_stage_inst_dmem_n17637) );
NAND2_X1 MEM_stage_inst_dmem_U15942 ( .A1(MEM_stage_inst_dmem_n17635), .A2(MEM_stage_inst_dmem_n17634), .ZN(MEM_stage_inst_dmem_n10547) );
NAND2_X1 MEM_stage_inst_dmem_U15941 ( .A1(EX_pipeline_reg_out_13), .A2(MEM_stage_inst_dmem_n17651), .ZN(MEM_stage_inst_dmem_n17634) );
NAND2_X1 MEM_stage_inst_dmem_U15940 ( .A1(MEM_stage_inst_dmem_ram_2296), .A2(MEM_stage_inst_dmem_n17650), .ZN(MEM_stage_inst_dmem_n17635) );
NAND2_X1 MEM_stage_inst_dmem_U15939 ( .A1(MEM_stage_inst_dmem_n17633), .A2(MEM_stage_inst_dmem_n17632), .ZN(MEM_stage_inst_dmem_n10548) );
NAND2_X1 MEM_stage_inst_dmem_U15938 ( .A1(EX_pipeline_reg_out_14), .A2(MEM_stage_inst_dmem_n17651), .ZN(MEM_stage_inst_dmem_n17632) );
NAND2_X1 MEM_stage_inst_dmem_U15937 ( .A1(MEM_stage_inst_dmem_ram_2297), .A2(MEM_stage_inst_dmem_n17650), .ZN(MEM_stage_inst_dmem_n17633) );
NAND2_X1 MEM_stage_inst_dmem_U15936 ( .A1(MEM_stage_inst_dmem_n17631), .A2(MEM_stage_inst_dmem_n17630), .ZN(MEM_stage_inst_dmem_n10549) );
NAND2_X1 MEM_stage_inst_dmem_U15935 ( .A1(EX_pipeline_reg_out_15), .A2(MEM_stage_inst_dmem_n17651), .ZN(MEM_stage_inst_dmem_n17630) );
NAND2_X1 MEM_stage_inst_dmem_U15934 ( .A1(MEM_stage_inst_dmem_ram_2298), .A2(MEM_stage_inst_dmem_n17650), .ZN(MEM_stage_inst_dmem_n17631) );
NAND2_X1 MEM_stage_inst_dmem_U15933 ( .A1(MEM_stage_inst_dmem_n17629), .A2(MEM_stage_inst_dmem_n17628), .ZN(MEM_stage_inst_dmem_n10550) );
NAND2_X1 MEM_stage_inst_dmem_U15932 ( .A1(EX_pipeline_reg_out_16), .A2(MEM_stage_inst_dmem_n17651), .ZN(MEM_stage_inst_dmem_n17628) );
NAND2_X1 MEM_stage_inst_dmem_U15931 ( .A1(MEM_stage_inst_dmem_ram_2299), .A2(MEM_stage_inst_dmem_n17650), .ZN(MEM_stage_inst_dmem_n17629) );
NAND2_X1 MEM_stage_inst_dmem_U15930 ( .A1(MEM_stage_inst_dmem_n17627), .A2(MEM_stage_inst_dmem_n17626), .ZN(MEM_stage_inst_dmem_n10551) );
NAND2_X1 MEM_stage_inst_dmem_U15929 ( .A1(EX_pipeline_reg_out_17), .A2(MEM_stage_inst_dmem_n17651), .ZN(MEM_stage_inst_dmem_n17626) );
NAND2_X1 MEM_stage_inst_dmem_U15928 ( .A1(MEM_stage_inst_dmem_ram_2300), .A2(MEM_stage_inst_dmem_n17650), .ZN(MEM_stage_inst_dmem_n17627) );
NAND2_X1 MEM_stage_inst_dmem_U15927 ( .A1(MEM_stage_inst_dmem_n17625), .A2(MEM_stage_inst_dmem_n17624), .ZN(MEM_stage_inst_dmem_n10552) );
NAND2_X1 MEM_stage_inst_dmem_U15926 ( .A1(EX_pipeline_reg_out_18), .A2(MEM_stage_inst_dmem_n17651), .ZN(MEM_stage_inst_dmem_n17624) );
NAND2_X1 MEM_stage_inst_dmem_U15925 ( .A1(MEM_stage_inst_dmem_ram_2301), .A2(MEM_stage_inst_dmem_n17650), .ZN(MEM_stage_inst_dmem_n17625) );
NAND2_X1 MEM_stage_inst_dmem_U15924 ( .A1(MEM_stage_inst_dmem_n17623), .A2(MEM_stage_inst_dmem_n17622), .ZN(MEM_stage_inst_dmem_n10553) );
NAND2_X1 MEM_stage_inst_dmem_U15923 ( .A1(EX_pipeline_reg_out_19), .A2(MEM_stage_inst_dmem_n17651), .ZN(MEM_stage_inst_dmem_n17622) );
NAND2_X1 MEM_stage_inst_dmem_U15922 ( .A1(MEM_stage_inst_dmem_ram_2302), .A2(MEM_stage_inst_dmem_n17650), .ZN(MEM_stage_inst_dmem_n17623) );
NAND2_X1 MEM_stage_inst_dmem_U15921 ( .A1(MEM_stage_inst_dmem_n17621), .A2(MEM_stage_inst_dmem_n17620), .ZN(MEM_stage_inst_dmem_n10554) );
NAND2_X1 MEM_stage_inst_dmem_U15920 ( .A1(EX_pipeline_reg_out_20), .A2(MEM_stage_inst_dmem_n17651), .ZN(MEM_stage_inst_dmem_n17620) );
INV_X1 MEM_stage_inst_dmem_U15919 ( .A(MEM_stage_inst_dmem_n17650), .ZN(MEM_stage_inst_dmem_n17651) );
NAND2_X1 MEM_stage_inst_dmem_U15918 ( .A1(MEM_stage_inst_dmem_ram_2303), .A2(MEM_stage_inst_dmem_n17650), .ZN(MEM_stage_inst_dmem_n17621) );
NAND2_X1 MEM_stage_inst_dmem_U15917 ( .A1(MEM_stage_inst_dmem_n20934), .A2(MEM_stage_inst_dmem_n18138), .ZN(MEM_stage_inst_dmem_n17650) );
NOR2_X2 MEM_stage_inst_dmem_U15916 ( .A1(MEM_stage_inst_dmem_n17619), .A2(MEM_stage_inst_dmem_n20932), .ZN(MEM_stage_inst_dmem_n18138) );
NAND2_X1 MEM_stage_inst_dmem_U15915 ( .A1(MEM_stage_inst_dmem_n17618), .A2(MEM_stage_inst_dmem_n17617), .ZN(MEM_stage_inst_dmem_n20932) );
NAND2_X1 MEM_stage_inst_dmem_U15914 ( .A1(MEM_stage_inst_dmem_n17616), .A2(MEM_stage_inst_dmem_n17615), .ZN(MEM_stage_inst_dmem_n10555) );
NAND2_X1 MEM_stage_inst_dmem_U15913 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n17614), .ZN(MEM_stage_inst_dmem_n17615) );
NAND2_X1 MEM_stage_inst_dmem_U15912 ( .A1(MEM_stage_inst_dmem_ram_2304), .A2(MEM_stage_inst_dmem_n17613), .ZN(MEM_stage_inst_dmem_n17616) );
NAND2_X1 MEM_stage_inst_dmem_U15911 ( .A1(MEM_stage_inst_dmem_n17612), .A2(MEM_stage_inst_dmem_n17611), .ZN(MEM_stage_inst_dmem_n10556) );
NAND2_X1 MEM_stage_inst_dmem_U15910 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n17614), .ZN(MEM_stage_inst_dmem_n17611) );
NAND2_X1 MEM_stage_inst_dmem_U15909 ( .A1(MEM_stage_inst_dmem_ram_2305), .A2(MEM_stage_inst_dmem_n17613), .ZN(MEM_stage_inst_dmem_n17612) );
NAND2_X1 MEM_stage_inst_dmem_U15908 ( .A1(MEM_stage_inst_dmem_n17610), .A2(MEM_stage_inst_dmem_n17609), .ZN(MEM_stage_inst_dmem_n10557) );
NAND2_X1 MEM_stage_inst_dmem_U15907 ( .A1(MEM_stage_inst_dmem_n18027), .A2(MEM_stage_inst_dmem_n17614), .ZN(MEM_stage_inst_dmem_n17609) );
NAND2_X1 MEM_stage_inst_dmem_U15906 ( .A1(MEM_stage_inst_dmem_ram_2306), .A2(MEM_stage_inst_dmem_n17613), .ZN(MEM_stage_inst_dmem_n17610) );
NAND2_X1 MEM_stage_inst_dmem_U15905 ( .A1(MEM_stage_inst_dmem_n17608), .A2(MEM_stage_inst_dmem_n17607), .ZN(MEM_stage_inst_dmem_n10558) );
NAND2_X1 MEM_stage_inst_dmem_U15904 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n17614), .ZN(MEM_stage_inst_dmem_n17607) );
NAND2_X1 MEM_stage_inst_dmem_U15903 ( .A1(MEM_stage_inst_dmem_ram_2307), .A2(MEM_stage_inst_dmem_n17613), .ZN(MEM_stage_inst_dmem_n17608) );
NAND2_X1 MEM_stage_inst_dmem_U15902 ( .A1(MEM_stage_inst_dmem_n17606), .A2(MEM_stage_inst_dmem_n17605), .ZN(MEM_stage_inst_dmem_n10559) );
NAND2_X1 MEM_stage_inst_dmem_U15901 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n17614), .ZN(MEM_stage_inst_dmem_n17605) );
NAND2_X1 MEM_stage_inst_dmem_U15900 ( .A1(MEM_stage_inst_dmem_ram_2308), .A2(MEM_stage_inst_dmem_n17613), .ZN(MEM_stage_inst_dmem_n17606) );
NAND2_X1 MEM_stage_inst_dmem_U15899 ( .A1(MEM_stage_inst_dmem_n17604), .A2(MEM_stage_inst_dmem_n17603), .ZN(MEM_stage_inst_dmem_n10560) );
NAND2_X1 MEM_stage_inst_dmem_U15898 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n17614), .ZN(MEM_stage_inst_dmem_n17603) );
NAND2_X1 MEM_stage_inst_dmem_U15897 ( .A1(MEM_stage_inst_dmem_ram_2309), .A2(MEM_stage_inst_dmem_n17613), .ZN(MEM_stage_inst_dmem_n17604) );
NAND2_X1 MEM_stage_inst_dmem_U15896 ( .A1(MEM_stage_inst_dmem_n17602), .A2(MEM_stage_inst_dmem_n17601), .ZN(MEM_stage_inst_dmem_n10561) );
NAND2_X1 MEM_stage_inst_dmem_U15895 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n17614), .ZN(MEM_stage_inst_dmem_n17601) );
NAND2_X1 MEM_stage_inst_dmem_U15894 ( .A1(MEM_stage_inst_dmem_ram_2310), .A2(MEM_stage_inst_dmem_n17613), .ZN(MEM_stage_inst_dmem_n17602) );
NAND2_X1 MEM_stage_inst_dmem_U15893 ( .A1(MEM_stage_inst_dmem_n17600), .A2(MEM_stage_inst_dmem_n17599), .ZN(MEM_stage_inst_dmem_n10562) );
NAND2_X1 MEM_stage_inst_dmem_U15892 ( .A1(MEM_stage_inst_dmem_n112), .A2(MEM_stage_inst_dmem_n17614), .ZN(MEM_stage_inst_dmem_n17599) );
NAND2_X1 MEM_stage_inst_dmem_U15891 ( .A1(MEM_stage_inst_dmem_ram_2311), .A2(MEM_stage_inst_dmem_n17613), .ZN(MEM_stage_inst_dmem_n17600) );
NAND2_X1 MEM_stage_inst_dmem_U15890 ( .A1(MEM_stage_inst_dmem_n17598), .A2(MEM_stage_inst_dmem_n17597), .ZN(MEM_stage_inst_dmem_n10563) );
NAND2_X1 MEM_stage_inst_dmem_U15889 ( .A1(MEM_stage_inst_dmem_n18013), .A2(MEM_stage_inst_dmem_n17614), .ZN(MEM_stage_inst_dmem_n17597) );
NAND2_X1 MEM_stage_inst_dmem_U15888 ( .A1(MEM_stage_inst_dmem_ram_2312), .A2(MEM_stage_inst_dmem_n17613), .ZN(MEM_stage_inst_dmem_n17598) );
NAND2_X1 MEM_stage_inst_dmem_U15887 ( .A1(MEM_stage_inst_dmem_n17596), .A2(MEM_stage_inst_dmem_n17595), .ZN(MEM_stage_inst_dmem_n10564) );
NAND2_X1 MEM_stage_inst_dmem_U15886 ( .A1(MEM_stage_inst_dmem_n96), .A2(MEM_stage_inst_dmem_n17614), .ZN(MEM_stage_inst_dmem_n17595) );
NAND2_X1 MEM_stage_inst_dmem_U15885 ( .A1(MEM_stage_inst_dmem_ram_2313), .A2(MEM_stage_inst_dmem_n17613), .ZN(MEM_stage_inst_dmem_n17596) );
NAND2_X1 MEM_stage_inst_dmem_U15884 ( .A1(MEM_stage_inst_dmem_n17594), .A2(MEM_stage_inst_dmem_n17593), .ZN(MEM_stage_inst_dmem_n10565) );
NAND2_X1 MEM_stage_inst_dmem_U15883 ( .A1(MEM_stage_inst_dmem_n18007), .A2(MEM_stage_inst_dmem_n17614), .ZN(MEM_stage_inst_dmem_n17593) );
NAND2_X1 MEM_stage_inst_dmem_U15882 ( .A1(MEM_stage_inst_dmem_ram_2314), .A2(MEM_stage_inst_dmem_n17613), .ZN(MEM_stage_inst_dmem_n17594) );
NAND2_X1 MEM_stage_inst_dmem_U15881 ( .A1(MEM_stage_inst_dmem_n17592), .A2(MEM_stage_inst_dmem_n17591), .ZN(MEM_stage_inst_dmem_n10566) );
NAND2_X1 MEM_stage_inst_dmem_U15880 ( .A1(MEM_stage_inst_dmem_n18004), .A2(MEM_stage_inst_dmem_n17614), .ZN(MEM_stage_inst_dmem_n17591) );
NAND2_X1 MEM_stage_inst_dmem_U15879 ( .A1(MEM_stage_inst_dmem_ram_2315), .A2(MEM_stage_inst_dmem_n17613), .ZN(MEM_stage_inst_dmem_n17592) );
NAND2_X1 MEM_stage_inst_dmem_U15878 ( .A1(MEM_stage_inst_dmem_n17590), .A2(MEM_stage_inst_dmem_n17589), .ZN(MEM_stage_inst_dmem_n10567) );
NAND2_X1 MEM_stage_inst_dmem_U15877 ( .A1(MEM_stage_inst_dmem_n18001), .A2(MEM_stage_inst_dmem_n17614), .ZN(MEM_stage_inst_dmem_n17589) );
NAND2_X1 MEM_stage_inst_dmem_U15876 ( .A1(MEM_stage_inst_dmem_ram_2316), .A2(MEM_stage_inst_dmem_n17613), .ZN(MEM_stage_inst_dmem_n17590) );
NAND2_X1 MEM_stage_inst_dmem_U15875 ( .A1(MEM_stage_inst_dmem_n17588), .A2(MEM_stage_inst_dmem_n17587), .ZN(MEM_stage_inst_dmem_n10568) );
NAND2_X1 MEM_stage_inst_dmem_U15874 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n17614), .ZN(MEM_stage_inst_dmem_n17587) );
NAND2_X1 MEM_stage_inst_dmem_U15873 ( .A1(MEM_stage_inst_dmem_ram_2317), .A2(MEM_stage_inst_dmem_n17613), .ZN(MEM_stage_inst_dmem_n17588) );
NAND2_X1 MEM_stage_inst_dmem_U15872 ( .A1(MEM_stage_inst_dmem_n17586), .A2(MEM_stage_inst_dmem_n17585), .ZN(MEM_stage_inst_dmem_n10569) );
NAND2_X1 MEM_stage_inst_dmem_U15871 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n17614), .ZN(MEM_stage_inst_dmem_n17585) );
NAND2_X1 MEM_stage_inst_dmem_U15870 ( .A1(MEM_stage_inst_dmem_ram_2318), .A2(MEM_stage_inst_dmem_n17613), .ZN(MEM_stage_inst_dmem_n17586) );
NAND2_X1 MEM_stage_inst_dmem_U15869 ( .A1(MEM_stage_inst_dmem_n17584), .A2(MEM_stage_inst_dmem_n17583), .ZN(MEM_stage_inst_dmem_n10570) );
NAND2_X1 MEM_stage_inst_dmem_U15868 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n17614), .ZN(MEM_stage_inst_dmem_n17583) );
NAND2_X1 MEM_stage_inst_dmem_U15867 ( .A1(MEM_stage_inst_dmem_ram_2319), .A2(MEM_stage_inst_dmem_n17613), .ZN(MEM_stage_inst_dmem_n17584) );
NAND2_X1 MEM_stage_inst_dmem_U15866 ( .A1(MEM_stage_inst_dmem_n21465), .A2(MEM_stage_inst_dmem_n17582), .ZN(MEM_stage_inst_dmem_n17613) );
NAND2_X1 MEM_stage_inst_dmem_U15865 ( .A1(MEM_stage_inst_dmem_n17581), .A2(MEM_stage_inst_dmem_n17580), .ZN(MEM_stage_inst_dmem_n10571) );
NAND2_X1 MEM_stage_inst_dmem_U15864 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n17579), .ZN(MEM_stage_inst_dmem_n17580) );
NAND2_X1 MEM_stage_inst_dmem_U15863 ( .A1(MEM_stage_inst_dmem_ram_2320), .A2(MEM_stage_inst_dmem_n17578), .ZN(MEM_stage_inst_dmem_n17581) );
NAND2_X1 MEM_stage_inst_dmem_U15862 ( .A1(MEM_stage_inst_dmem_n17577), .A2(MEM_stage_inst_dmem_n17576), .ZN(MEM_stage_inst_dmem_n10572) );
NAND2_X1 MEM_stage_inst_dmem_U15861 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n17579), .ZN(MEM_stage_inst_dmem_n17576) );
NAND2_X1 MEM_stage_inst_dmem_U15860 ( .A1(MEM_stage_inst_dmem_ram_2321), .A2(MEM_stage_inst_dmem_n17578), .ZN(MEM_stage_inst_dmem_n17577) );
NAND2_X1 MEM_stage_inst_dmem_U15859 ( .A1(MEM_stage_inst_dmem_n17575), .A2(MEM_stage_inst_dmem_n17574), .ZN(MEM_stage_inst_dmem_n10573) );
NAND2_X1 MEM_stage_inst_dmem_U15858 ( .A1(MEM_stage_inst_dmem_n18027), .A2(MEM_stage_inst_dmem_n17579), .ZN(MEM_stage_inst_dmem_n17574) );
NAND2_X1 MEM_stage_inst_dmem_U15857 ( .A1(MEM_stage_inst_dmem_ram_2322), .A2(MEM_stage_inst_dmem_n17578), .ZN(MEM_stage_inst_dmem_n17575) );
NAND2_X1 MEM_stage_inst_dmem_U15856 ( .A1(MEM_stage_inst_dmem_n17573), .A2(MEM_stage_inst_dmem_n17572), .ZN(MEM_stage_inst_dmem_n10574) );
NAND2_X1 MEM_stage_inst_dmem_U15855 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n17579), .ZN(MEM_stage_inst_dmem_n17572) );
NAND2_X1 MEM_stage_inst_dmem_U15854 ( .A1(MEM_stage_inst_dmem_ram_2323), .A2(MEM_stage_inst_dmem_n17578), .ZN(MEM_stage_inst_dmem_n17573) );
NAND2_X1 MEM_stage_inst_dmem_U15853 ( .A1(MEM_stage_inst_dmem_n17571), .A2(MEM_stage_inst_dmem_n17570), .ZN(MEM_stage_inst_dmem_n10575) );
NAND2_X1 MEM_stage_inst_dmem_U15852 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n17579), .ZN(MEM_stage_inst_dmem_n17570) );
NAND2_X1 MEM_stage_inst_dmem_U15851 ( .A1(MEM_stage_inst_dmem_ram_2324), .A2(MEM_stage_inst_dmem_n17578), .ZN(MEM_stage_inst_dmem_n17571) );
NAND2_X1 MEM_stage_inst_dmem_U15850 ( .A1(MEM_stage_inst_dmem_n17569), .A2(MEM_stage_inst_dmem_n17568), .ZN(MEM_stage_inst_dmem_n10576) );
NAND2_X1 MEM_stage_inst_dmem_U15849 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n17579), .ZN(MEM_stage_inst_dmem_n17568) );
NAND2_X1 MEM_stage_inst_dmem_U15848 ( .A1(MEM_stage_inst_dmem_ram_2325), .A2(MEM_stage_inst_dmem_n17578), .ZN(MEM_stage_inst_dmem_n17569) );
NAND2_X1 MEM_stage_inst_dmem_U15847 ( .A1(MEM_stage_inst_dmem_n17567), .A2(MEM_stage_inst_dmem_n17566), .ZN(MEM_stage_inst_dmem_n10577) );
NAND2_X1 MEM_stage_inst_dmem_U15846 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n17579), .ZN(MEM_stage_inst_dmem_n17566) );
NAND2_X1 MEM_stage_inst_dmem_U15845 ( .A1(MEM_stage_inst_dmem_ram_2326), .A2(MEM_stage_inst_dmem_n17578), .ZN(MEM_stage_inst_dmem_n17567) );
NAND2_X1 MEM_stage_inst_dmem_U15844 ( .A1(MEM_stage_inst_dmem_n17565), .A2(MEM_stage_inst_dmem_n17564), .ZN(MEM_stage_inst_dmem_n10578) );
NAND2_X1 MEM_stage_inst_dmem_U15843 ( .A1(MEM_stage_inst_dmem_n16361), .A2(MEM_stage_inst_dmem_n17579), .ZN(MEM_stage_inst_dmem_n17564) );
NAND2_X1 MEM_stage_inst_dmem_U15842 ( .A1(MEM_stage_inst_dmem_ram_2327), .A2(MEM_stage_inst_dmem_n17578), .ZN(MEM_stage_inst_dmem_n17565) );
NAND2_X1 MEM_stage_inst_dmem_U15841 ( .A1(MEM_stage_inst_dmem_n17563), .A2(MEM_stage_inst_dmem_n17562), .ZN(MEM_stage_inst_dmem_n10579) );
NAND2_X1 MEM_stage_inst_dmem_U15840 ( .A1(MEM_stage_inst_dmem_n18013), .A2(MEM_stage_inst_dmem_n17579), .ZN(MEM_stage_inst_dmem_n17562) );
NAND2_X1 MEM_stage_inst_dmem_U15839 ( .A1(MEM_stage_inst_dmem_ram_2328), .A2(MEM_stage_inst_dmem_n17578), .ZN(MEM_stage_inst_dmem_n17563) );
NAND2_X1 MEM_stage_inst_dmem_U15838 ( .A1(MEM_stage_inst_dmem_n17561), .A2(MEM_stage_inst_dmem_n17560), .ZN(MEM_stage_inst_dmem_n10580) );
NAND2_X1 MEM_stage_inst_dmem_U15837 ( .A1(MEM_stage_inst_dmem_n96), .A2(MEM_stage_inst_dmem_n17579), .ZN(MEM_stage_inst_dmem_n17560) );
NAND2_X1 MEM_stage_inst_dmem_U15836 ( .A1(MEM_stage_inst_dmem_ram_2329), .A2(MEM_stage_inst_dmem_n17578), .ZN(MEM_stage_inst_dmem_n17561) );
NAND2_X1 MEM_stage_inst_dmem_U15835 ( .A1(MEM_stage_inst_dmem_n17559), .A2(MEM_stage_inst_dmem_n17558), .ZN(MEM_stage_inst_dmem_n10581) );
NAND2_X1 MEM_stage_inst_dmem_U15834 ( .A1(MEM_stage_inst_dmem_n18007), .A2(MEM_stage_inst_dmem_n17579), .ZN(MEM_stage_inst_dmem_n17558) );
NAND2_X1 MEM_stage_inst_dmem_U15833 ( .A1(MEM_stage_inst_dmem_ram_2330), .A2(MEM_stage_inst_dmem_n17578), .ZN(MEM_stage_inst_dmem_n17559) );
NAND2_X1 MEM_stage_inst_dmem_U15832 ( .A1(MEM_stage_inst_dmem_n17557), .A2(MEM_stage_inst_dmem_n17556), .ZN(MEM_stage_inst_dmem_n10582) );
NAND2_X1 MEM_stage_inst_dmem_U15831 ( .A1(MEM_stage_inst_dmem_n18004), .A2(MEM_stage_inst_dmem_n17579), .ZN(MEM_stage_inst_dmem_n17556) );
NAND2_X1 MEM_stage_inst_dmem_U15830 ( .A1(MEM_stage_inst_dmem_ram_2331), .A2(MEM_stage_inst_dmem_n17578), .ZN(MEM_stage_inst_dmem_n17557) );
NAND2_X1 MEM_stage_inst_dmem_U15829 ( .A1(MEM_stage_inst_dmem_n17555), .A2(MEM_stage_inst_dmem_n17554), .ZN(MEM_stage_inst_dmem_n10583) );
NAND2_X1 MEM_stage_inst_dmem_U15828 ( .A1(MEM_stage_inst_dmem_n18001), .A2(MEM_stage_inst_dmem_n17579), .ZN(MEM_stage_inst_dmem_n17554) );
NAND2_X1 MEM_stage_inst_dmem_U15827 ( .A1(MEM_stage_inst_dmem_ram_2332), .A2(MEM_stage_inst_dmem_n17578), .ZN(MEM_stage_inst_dmem_n17555) );
NAND2_X1 MEM_stage_inst_dmem_U15826 ( .A1(MEM_stage_inst_dmem_n17553), .A2(MEM_stage_inst_dmem_n17552), .ZN(MEM_stage_inst_dmem_n10584) );
NAND2_X1 MEM_stage_inst_dmem_U15825 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n17579), .ZN(MEM_stage_inst_dmem_n17552) );
NAND2_X1 MEM_stage_inst_dmem_U15824 ( .A1(MEM_stage_inst_dmem_ram_2333), .A2(MEM_stage_inst_dmem_n17578), .ZN(MEM_stage_inst_dmem_n17553) );
NAND2_X1 MEM_stage_inst_dmem_U15823 ( .A1(MEM_stage_inst_dmem_n17551), .A2(MEM_stage_inst_dmem_n17550), .ZN(MEM_stage_inst_dmem_n10585) );
NAND2_X1 MEM_stage_inst_dmem_U15822 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n17579), .ZN(MEM_stage_inst_dmem_n17550) );
NAND2_X1 MEM_stage_inst_dmem_U15821 ( .A1(MEM_stage_inst_dmem_ram_2334), .A2(MEM_stage_inst_dmem_n17578), .ZN(MEM_stage_inst_dmem_n17551) );
NAND2_X1 MEM_stage_inst_dmem_U15820 ( .A1(MEM_stage_inst_dmem_n17549), .A2(MEM_stage_inst_dmem_n17548), .ZN(MEM_stage_inst_dmem_n10586) );
NAND2_X1 MEM_stage_inst_dmem_U15819 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n17579), .ZN(MEM_stage_inst_dmem_n17548) );
INV_X1 MEM_stage_inst_dmem_U15818 ( .A(MEM_stage_inst_dmem_n17578), .ZN(MEM_stage_inst_dmem_n17579) );
NAND2_X1 MEM_stage_inst_dmem_U15817 ( .A1(MEM_stage_inst_dmem_ram_2335), .A2(MEM_stage_inst_dmem_n17578), .ZN(MEM_stage_inst_dmem_n17549) );
NAND2_X1 MEM_stage_inst_dmem_U15816 ( .A1(MEM_stage_inst_dmem_n21429), .A2(MEM_stage_inst_dmem_n17582), .ZN(MEM_stage_inst_dmem_n17578) );
NAND2_X1 MEM_stage_inst_dmem_U15815 ( .A1(MEM_stage_inst_dmem_n17547), .A2(MEM_stage_inst_dmem_n17546), .ZN(MEM_stage_inst_dmem_n10587) );
NAND2_X1 MEM_stage_inst_dmem_U15814 ( .A1(EX_pipeline_reg_out_5), .A2(MEM_stage_inst_dmem_n17545), .ZN(MEM_stage_inst_dmem_n17546) );
NAND2_X1 MEM_stage_inst_dmem_U15813 ( .A1(MEM_stage_inst_dmem_ram_2336), .A2(MEM_stage_inst_dmem_n17544), .ZN(MEM_stage_inst_dmem_n17547) );
NAND2_X1 MEM_stage_inst_dmem_U15812 ( .A1(MEM_stage_inst_dmem_n17543), .A2(MEM_stage_inst_dmem_n17542), .ZN(MEM_stage_inst_dmem_n10588) );
NAND2_X1 MEM_stage_inst_dmem_U15811 ( .A1(EX_pipeline_reg_out_6), .A2(MEM_stage_inst_dmem_n17545), .ZN(MEM_stage_inst_dmem_n17542) );
NAND2_X1 MEM_stage_inst_dmem_U15810 ( .A1(MEM_stage_inst_dmem_ram_2337), .A2(MEM_stage_inst_dmem_n17544), .ZN(MEM_stage_inst_dmem_n17543) );
NAND2_X1 MEM_stage_inst_dmem_U15809 ( .A1(MEM_stage_inst_dmem_n17541), .A2(MEM_stage_inst_dmem_n17540), .ZN(MEM_stage_inst_dmem_n10589) );
NAND2_X1 MEM_stage_inst_dmem_U15808 ( .A1(EX_pipeline_reg_out_7), .A2(MEM_stage_inst_dmem_n17545), .ZN(MEM_stage_inst_dmem_n17540) );
NAND2_X1 MEM_stage_inst_dmem_U15807 ( .A1(MEM_stage_inst_dmem_ram_2338), .A2(MEM_stage_inst_dmem_n17544), .ZN(MEM_stage_inst_dmem_n17541) );
NAND2_X1 MEM_stage_inst_dmem_U15806 ( .A1(MEM_stage_inst_dmem_n17539), .A2(MEM_stage_inst_dmem_n17538), .ZN(MEM_stage_inst_dmem_n10590) );
NAND2_X1 MEM_stage_inst_dmem_U15805 ( .A1(EX_pipeline_reg_out_8), .A2(MEM_stage_inst_dmem_n17545), .ZN(MEM_stage_inst_dmem_n17538) );
NAND2_X1 MEM_stage_inst_dmem_U15804 ( .A1(MEM_stage_inst_dmem_ram_2339), .A2(MEM_stage_inst_dmem_n17544), .ZN(MEM_stage_inst_dmem_n17539) );
NAND2_X1 MEM_stage_inst_dmem_U15803 ( .A1(MEM_stage_inst_dmem_n17537), .A2(MEM_stage_inst_dmem_n17536), .ZN(MEM_stage_inst_dmem_n10591) );
NAND2_X1 MEM_stage_inst_dmem_U15802 ( .A1(EX_pipeline_reg_out_9), .A2(MEM_stage_inst_dmem_n17545), .ZN(MEM_stage_inst_dmem_n17536) );
NAND2_X1 MEM_stage_inst_dmem_U15801 ( .A1(MEM_stage_inst_dmem_ram_2340), .A2(MEM_stage_inst_dmem_n17544), .ZN(MEM_stage_inst_dmem_n17537) );
NAND2_X1 MEM_stage_inst_dmem_U15800 ( .A1(MEM_stage_inst_dmem_n17535), .A2(MEM_stage_inst_dmem_n17534), .ZN(MEM_stage_inst_dmem_n10592) );
NAND2_X1 MEM_stage_inst_dmem_U15799 ( .A1(EX_pipeline_reg_out_10), .A2(MEM_stage_inst_dmem_n17545), .ZN(MEM_stage_inst_dmem_n17534) );
NAND2_X1 MEM_stage_inst_dmem_U15798 ( .A1(MEM_stage_inst_dmem_ram_2341), .A2(MEM_stage_inst_dmem_n17544), .ZN(MEM_stage_inst_dmem_n17535) );
NAND2_X1 MEM_stage_inst_dmem_U15797 ( .A1(MEM_stage_inst_dmem_n17533), .A2(MEM_stage_inst_dmem_n17532), .ZN(MEM_stage_inst_dmem_n10593) );
NAND2_X1 MEM_stage_inst_dmem_U15796 ( .A1(EX_pipeline_reg_out_11), .A2(MEM_stage_inst_dmem_n17545), .ZN(MEM_stage_inst_dmem_n17532) );
NAND2_X1 MEM_stage_inst_dmem_U15795 ( .A1(MEM_stage_inst_dmem_ram_2342), .A2(MEM_stage_inst_dmem_n17544), .ZN(MEM_stage_inst_dmem_n17533) );
NAND2_X1 MEM_stage_inst_dmem_U15794 ( .A1(MEM_stage_inst_dmem_n17531), .A2(MEM_stage_inst_dmem_n17530), .ZN(MEM_stage_inst_dmem_n10594) );
NAND2_X1 MEM_stage_inst_dmem_U15793 ( .A1(EX_pipeline_reg_out_12), .A2(MEM_stage_inst_dmem_n17545), .ZN(MEM_stage_inst_dmem_n17530) );
NAND2_X1 MEM_stage_inst_dmem_U15792 ( .A1(MEM_stage_inst_dmem_ram_2343), .A2(MEM_stage_inst_dmem_n17544), .ZN(MEM_stage_inst_dmem_n17531) );
NAND2_X1 MEM_stage_inst_dmem_U15791 ( .A1(MEM_stage_inst_dmem_n17529), .A2(MEM_stage_inst_dmem_n17528), .ZN(MEM_stage_inst_dmem_n10595) );
NAND2_X1 MEM_stage_inst_dmem_U15790 ( .A1(EX_pipeline_reg_out_13), .A2(MEM_stage_inst_dmem_n17545), .ZN(MEM_stage_inst_dmem_n17528) );
NAND2_X1 MEM_stage_inst_dmem_U15789 ( .A1(MEM_stage_inst_dmem_ram_2344), .A2(MEM_stage_inst_dmem_n17544), .ZN(MEM_stage_inst_dmem_n17529) );
NAND2_X1 MEM_stage_inst_dmem_U15788 ( .A1(MEM_stage_inst_dmem_n17527), .A2(MEM_stage_inst_dmem_n17526), .ZN(MEM_stage_inst_dmem_n10596) );
NAND2_X1 MEM_stage_inst_dmem_U15787 ( .A1(EX_pipeline_reg_out_14), .A2(MEM_stage_inst_dmem_n17545), .ZN(MEM_stage_inst_dmem_n17526) );
NAND2_X1 MEM_stage_inst_dmem_U15786 ( .A1(MEM_stage_inst_dmem_ram_2345), .A2(MEM_stage_inst_dmem_n17544), .ZN(MEM_stage_inst_dmem_n17527) );
NAND2_X1 MEM_stage_inst_dmem_U15785 ( .A1(MEM_stage_inst_dmem_n17525), .A2(MEM_stage_inst_dmem_n17524), .ZN(MEM_stage_inst_dmem_n10597) );
NAND2_X1 MEM_stage_inst_dmem_U15784 ( .A1(EX_pipeline_reg_out_15), .A2(MEM_stage_inst_dmem_n17545), .ZN(MEM_stage_inst_dmem_n17524) );
NAND2_X1 MEM_stage_inst_dmem_U15783 ( .A1(MEM_stage_inst_dmem_ram_2346), .A2(MEM_stage_inst_dmem_n17544), .ZN(MEM_stage_inst_dmem_n17525) );
NAND2_X1 MEM_stage_inst_dmem_U15782 ( .A1(MEM_stage_inst_dmem_n17523), .A2(MEM_stage_inst_dmem_n17522), .ZN(MEM_stage_inst_dmem_n10598) );
NAND2_X1 MEM_stage_inst_dmem_U15781 ( .A1(EX_pipeline_reg_out_16), .A2(MEM_stage_inst_dmem_n17545), .ZN(MEM_stage_inst_dmem_n17522) );
NAND2_X1 MEM_stage_inst_dmem_U15780 ( .A1(MEM_stage_inst_dmem_ram_2347), .A2(MEM_stage_inst_dmem_n17544), .ZN(MEM_stage_inst_dmem_n17523) );
NAND2_X1 MEM_stage_inst_dmem_U15779 ( .A1(MEM_stage_inst_dmem_n17521), .A2(MEM_stage_inst_dmem_n17520), .ZN(MEM_stage_inst_dmem_n10599) );
NAND2_X1 MEM_stage_inst_dmem_U15778 ( .A1(EX_pipeline_reg_out_17), .A2(MEM_stage_inst_dmem_n17545), .ZN(MEM_stage_inst_dmem_n17520) );
NAND2_X1 MEM_stage_inst_dmem_U15777 ( .A1(MEM_stage_inst_dmem_ram_2348), .A2(MEM_stage_inst_dmem_n17544), .ZN(MEM_stage_inst_dmem_n17521) );
NAND2_X1 MEM_stage_inst_dmem_U15776 ( .A1(MEM_stage_inst_dmem_n17519), .A2(MEM_stage_inst_dmem_n17518), .ZN(MEM_stage_inst_dmem_n10600) );
NAND2_X1 MEM_stage_inst_dmem_U15775 ( .A1(EX_pipeline_reg_out_18), .A2(MEM_stage_inst_dmem_n17545), .ZN(MEM_stage_inst_dmem_n17518) );
NAND2_X1 MEM_stage_inst_dmem_U15774 ( .A1(MEM_stage_inst_dmem_ram_2349), .A2(MEM_stage_inst_dmem_n17544), .ZN(MEM_stage_inst_dmem_n17519) );
NAND2_X1 MEM_stage_inst_dmem_U15773 ( .A1(MEM_stage_inst_dmem_n17517), .A2(MEM_stage_inst_dmem_n17516), .ZN(MEM_stage_inst_dmem_n10601) );
NAND2_X1 MEM_stage_inst_dmem_U15772 ( .A1(EX_pipeline_reg_out_19), .A2(MEM_stage_inst_dmem_n17545), .ZN(MEM_stage_inst_dmem_n17516) );
NAND2_X1 MEM_stage_inst_dmem_U15771 ( .A1(MEM_stage_inst_dmem_ram_2350), .A2(MEM_stage_inst_dmem_n17544), .ZN(MEM_stage_inst_dmem_n17517) );
NAND2_X1 MEM_stage_inst_dmem_U15770 ( .A1(MEM_stage_inst_dmem_n17515), .A2(MEM_stage_inst_dmem_n17514), .ZN(MEM_stage_inst_dmem_n10602) );
NAND2_X1 MEM_stage_inst_dmem_U15769 ( .A1(EX_pipeline_reg_out_20), .A2(MEM_stage_inst_dmem_n17545), .ZN(MEM_stage_inst_dmem_n17514) );
INV_X1 MEM_stage_inst_dmem_U15768 ( .A(MEM_stage_inst_dmem_n17544), .ZN(MEM_stage_inst_dmem_n17545) );
NAND2_X1 MEM_stage_inst_dmem_U15767 ( .A1(MEM_stage_inst_dmem_ram_2351), .A2(MEM_stage_inst_dmem_n17544), .ZN(MEM_stage_inst_dmem_n17515) );
NAND2_X1 MEM_stage_inst_dmem_U15766 ( .A1(MEM_stage_inst_dmem_n21394), .A2(MEM_stage_inst_dmem_n17582), .ZN(MEM_stage_inst_dmem_n17544) );
NAND2_X1 MEM_stage_inst_dmem_U15765 ( .A1(MEM_stage_inst_dmem_n17513), .A2(MEM_stage_inst_dmem_n17512), .ZN(MEM_stage_inst_dmem_n10603) );
NAND2_X1 MEM_stage_inst_dmem_U15764 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n17511), .ZN(MEM_stage_inst_dmem_n17512) );
NAND2_X1 MEM_stage_inst_dmem_U15763 ( .A1(MEM_stage_inst_dmem_ram_2352), .A2(MEM_stage_inst_dmem_n17510), .ZN(MEM_stage_inst_dmem_n17513) );
NAND2_X1 MEM_stage_inst_dmem_U15762 ( .A1(MEM_stage_inst_dmem_n17509), .A2(MEM_stage_inst_dmem_n17508), .ZN(MEM_stage_inst_dmem_n10604) );
NAND2_X1 MEM_stage_inst_dmem_U15761 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n17511), .ZN(MEM_stage_inst_dmem_n17508) );
NAND2_X1 MEM_stage_inst_dmem_U15760 ( .A1(MEM_stage_inst_dmem_ram_2353), .A2(MEM_stage_inst_dmem_n17510), .ZN(MEM_stage_inst_dmem_n17509) );
NAND2_X1 MEM_stage_inst_dmem_U15759 ( .A1(MEM_stage_inst_dmem_n17507), .A2(MEM_stage_inst_dmem_n17506), .ZN(MEM_stage_inst_dmem_n10605) );
NAND2_X1 MEM_stage_inst_dmem_U15758 ( .A1(MEM_stage_inst_dmem_n18027), .A2(MEM_stage_inst_dmem_n17511), .ZN(MEM_stage_inst_dmem_n17506) );
NAND2_X1 MEM_stage_inst_dmem_U15757 ( .A1(MEM_stage_inst_dmem_ram_2354), .A2(MEM_stage_inst_dmem_n17510), .ZN(MEM_stage_inst_dmem_n17507) );
NAND2_X1 MEM_stage_inst_dmem_U15756 ( .A1(MEM_stage_inst_dmem_n17505), .A2(MEM_stage_inst_dmem_n17504), .ZN(MEM_stage_inst_dmem_n10606) );
NAND2_X1 MEM_stage_inst_dmem_U15755 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n17511), .ZN(MEM_stage_inst_dmem_n17504) );
NAND2_X1 MEM_stage_inst_dmem_U15754 ( .A1(MEM_stage_inst_dmem_ram_2355), .A2(MEM_stage_inst_dmem_n17510), .ZN(MEM_stage_inst_dmem_n17505) );
NAND2_X1 MEM_stage_inst_dmem_U15753 ( .A1(MEM_stage_inst_dmem_n17503), .A2(MEM_stage_inst_dmem_n17502), .ZN(MEM_stage_inst_dmem_n10607) );
NAND2_X1 MEM_stage_inst_dmem_U15752 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n17511), .ZN(MEM_stage_inst_dmem_n17502) );
NAND2_X1 MEM_stage_inst_dmem_U15751 ( .A1(MEM_stage_inst_dmem_ram_2356), .A2(MEM_stage_inst_dmem_n17510), .ZN(MEM_stage_inst_dmem_n17503) );
NAND2_X1 MEM_stage_inst_dmem_U15750 ( .A1(MEM_stage_inst_dmem_n17501), .A2(MEM_stage_inst_dmem_n17500), .ZN(MEM_stage_inst_dmem_n10608) );
NAND2_X1 MEM_stage_inst_dmem_U15749 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n17511), .ZN(MEM_stage_inst_dmem_n17500) );
NAND2_X1 MEM_stage_inst_dmem_U15748 ( .A1(MEM_stage_inst_dmem_ram_2357), .A2(MEM_stage_inst_dmem_n17510), .ZN(MEM_stage_inst_dmem_n17501) );
NAND2_X1 MEM_stage_inst_dmem_U15747 ( .A1(MEM_stage_inst_dmem_n17499), .A2(MEM_stage_inst_dmem_n17498), .ZN(MEM_stage_inst_dmem_n10609) );
NAND2_X1 MEM_stage_inst_dmem_U15746 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n17511), .ZN(MEM_stage_inst_dmem_n17498) );
NAND2_X1 MEM_stage_inst_dmem_U15745 ( .A1(MEM_stage_inst_dmem_ram_2358), .A2(MEM_stage_inst_dmem_n17510), .ZN(MEM_stage_inst_dmem_n17499) );
NAND2_X1 MEM_stage_inst_dmem_U15744 ( .A1(MEM_stage_inst_dmem_n17497), .A2(MEM_stage_inst_dmem_n17496), .ZN(MEM_stage_inst_dmem_n10610) );
NAND2_X1 MEM_stage_inst_dmem_U15743 ( .A1(MEM_stage_inst_dmem_n112), .A2(MEM_stage_inst_dmem_n17511), .ZN(MEM_stage_inst_dmem_n17496) );
NAND2_X1 MEM_stage_inst_dmem_U15742 ( .A1(MEM_stage_inst_dmem_ram_2359), .A2(MEM_stage_inst_dmem_n17510), .ZN(MEM_stage_inst_dmem_n17497) );
NAND2_X1 MEM_stage_inst_dmem_U15741 ( .A1(MEM_stage_inst_dmem_n17495), .A2(MEM_stage_inst_dmem_n17494), .ZN(MEM_stage_inst_dmem_n10611) );
NAND2_X1 MEM_stage_inst_dmem_U15740 ( .A1(MEM_stage_inst_dmem_n18013), .A2(MEM_stage_inst_dmem_n17511), .ZN(MEM_stage_inst_dmem_n17494) );
NAND2_X1 MEM_stage_inst_dmem_U15739 ( .A1(MEM_stage_inst_dmem_ram_2360), .A2(MEM_stage_inst_dmem_n17510), .ZN(MEM_stage_inst_dmem_n17495) );
NAND2_X1 MEM_stage_inst_dmem_U15738 ( .A1(MEM_stage_inst_dmem_n17493), .A2(MEM_stage_inst_dmem_n17492), .ZN(MEM_stage_inst_dmem_n10612) );
NAND2_X1 MEM_stage_inst_dmem_U15737 ( .A1(MEM_stage_inst_dmem_n96), .A2(MEM_stage_inst_dmem_n17511), .ZN(MEM_stage_inst_dmem_n17492) );
NAND2_X1 MEM_stage_inst_dmem_U15736 ( .A1(MEM_stage_inst_dmem_ram_2361), .A2(MEM_stage_inst_dmem_n17510), .ZN(MEM_stage_inst_dmem_n17493) );
NAND2_X1 MEM_stage_inst_dmem_U15735 ( .A1(MEM_stage_inst_dmem_n17491), .A2(MEM_stage_inst_dmem_n17490), .ZN(MEM_stage_inst_dmem_n10613) );
NAND2_X1 MEM_stage_inst_dmem_U15734 ( .A1(MEM_stage_inst_dmem_n18007), .A2(MEM_stage_inst_dmem_n17511), .ZN(MEM_stage_inst_dmem_n17490) );
NAND2_X1 MEM_stage_inst_dmem_U15733 ( .A1(MEM_stage_inst_dmem_ram_2362), .A2(MEM_stage_inst_dmem_n17510), .ZN(MEM_stage_inst_dmem_n17491) );
NAND2_X1 MEM_stage_inst_dmem_U15732 ( .A1(MEM_stage_inst_dmem_n17489), .A2(MEM_stage_inst_dmem_n17488), .ZN(MEM_stage_inst_dmem_n10614) );
NAND2_X1 MEM_stage_inst_dmem_U15731 ( .A1(MEM_stage_inst_dmem_n18004), .A2(MEM_stage_inst_dmem_n17511), .ZN(MEM_stage_inst_dmem_n17488) );
NAND2_X1 MEM_stage_inst_dmem_U15730 ( .A1(MEM_stage_inst_dmem_ram_2363), .A2(MEM_stage_inst_dmem_n17510), .ZN(MEM_stage_inst_dmem_n17489) );
NAND2_X1 MEM_stage_inst_dmem_U15729 ( .A1(MEM_stage_inst_dmem_n17487), .A2(MEM_stage_inst_dmem_n17486), .ZN(MEM_stage_inst_dmem_n10615) );
NAND2_X1 MEM_stage_inst_dmem_U15728 ( .A1(MEM_stage_inst_dmem_n18001), .A2(MEM_stage_inst_dmem_n17511), .ZN(MEM_stage_inst_dmem_n17486) );
NAND2_X1 MEM_stage_inst_dmem_U15727 ( .A1(MEM_stage_inst_dmem_ram_2364), .A2(MEM_stage_inst_dmem_n17510), .ZN(MEM_stage_inst_dmem_n17487) );
NAND2_X1 MEM_stage_inst_dmem_U15726 ( .A1(MEM_stage_inst_dmem_n17485), .A2(MEM_stage_inst_dmem_n17484), .ZN(MEM_stage_inst_dmem_n10616) );
NAND2_X1 MEM_stage_inst_dmem_U15725 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n17511), .ZN(MEM_stage_inst_dmem_n17484) );
NAND2_X1 MEM_stage_inst_dmem_U15724 ( .A1(MEM_stage_inst_dmem_ram_2365), .A2(MEM_stage_inst_dmem_n17510), .ZN(MEM_stage_inst_dmem_n17485) );
NAND2_X1 MEM_stage_inst_dmem_U15723 ( .A1(MEM_stage_inst_dmem_n17483), .A2(MEM_stage_inst_dmem_n17482), .ZN(MEM_stage_inst_dmem_n10617) );
NAND2_X1 MEM_stage_inst_dmem_U15722 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n17511), .ZN(MEM_stage_inst_dmem_n17482) );
NAND2_X1 MEM_stage_inst_dmem_U15721 ( .A1(MEM_stage_inst_dmem_ram_2366), .A2(MEM_stage_inst_dmem_n17510), .ZN(MEM_stage_inst_dmem_n17483) );
NAND2_X1 MEM_stage_inst_dmem_U15720 ( .A1(MEM_stage_inst_dmem_n17481), .A2(MEM_stage_inst_dmem_n17480), .ZN(MEM_stage_inst_dmem_n10618) );
NAND2_X1 MEM_stage_inst_dmem_U15719 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n17511), .ZN(MEM_stage_inst_dmem_n17480) );
INV_X1 MEM_stage_inst_dmem_U15718 ( .A(MEM_stage_inst_dmem_n17510), .ZN(MEM_stage_inst_dmem_n17511) );
NAND2_X1 MEM_stage_inst_dmem_U15717 ( .A1(MEM_stage_inst_dmem_ram_2367), .A2(MEM_stage_inst_dmem_n17510), .ZN(MEM_stage_inst_dmem_n17481) );
NAND2_X1 MEM_stage_inst_dmem_U15716 ( .A1(MEM_stage_inst_dmem_n21359), .A2(MEM_stage_inst_dmem_n17582), .ZN(MEM_stage_inst_dmem_n17510) );
NAND2_X1 MEM_stage_inst_dmem_U15715 ( .A1(MEM_stage_inst_dmem_n17479), .A2(MEM_stage_inst_dmem_n17478), .ZN(MEM_stage_inst_dmem_n10619) );
NAND2_X1 MEM_stage_inst_dmem_U15714 ( .A1(EX_pipeline_reg_out_5), .A2(MEM_stage_inst_dmem_n17477), .ZN(MEM_stage_inst_dmem_n17478) );
NAND2_X1 MEM_stage_inst_dmem_U15713 ( .A1(MEM_stage_inst_dmem_ram_2368), .A2(MEM_stage_inst_dmem_n17476), .ZN(MEM_stage_inst_dmem_n17479) );
NAND2_X1 MEM_stage_inst_dmem_U15712 ( .A1(MEM_stage_inst_dmem_n17475), .A2(MEM_stage_inst_dmem_n17474), .ZN(MEM_stage_inst_dmem_n10620) );
NAND2_X1 MEM_stage_inst_dmem_U15711 ( .A1(EX_pipeline_reg_out_6), .A2(MEM_stage_inst_dmem_n17477), .ZN(MEM_stage_inst_dmem_n17474) );
NAND2_X1 MEM_stage_inst_dmem_U15710 ( .A1(MEM_stage_inst_dmem_ram_2369), .A2(MEM_stage_inst_dmem_n17476), .ZN(MEM_stage_inst_dmem_n17475) );
NAND2_X1 MEM_stage_inst_dmem_U15709 ( .A1(MEM_stage_inst_dmem_n17473), .A2(MEM_stage_inst_dmem_n17472), .ZN(MEM_stage_inst_dmem_n10621) );
NAND2_X1 MEM_stage_inst_dmem_U15708 ( .A1(EX_pipeline_reg_out_7), .A2(MEM_stage_inst_dmem_n17477), .ZN(MEM_stage_inst_dmem_n17472) );
NAND2_X1 MEM_stage_inst_dmem_U15707 ( .A1(MEM_stage_inst_dmem_ram_2370), .A2(MEM_stage_inst_dmem_n17476), .ZN(MEM_stage_inst_dmem_n17473) );
NAND2_X1 MEM_stage_inst_dmem_U15706 ( .A1(MEM_stage_inst_dmem_n17471), .A2(MEM_stage_inst_dmem_n17470), .ZN(MEM_stage_inst_dmem_n10622) );
NAND2_X1 MEM_stage_inst_dmem_U15705 ( .A1(EX_pipeline_reg_out_8), .A2(MEM_stage_inst_dmem_n17477), .ZN(MEM_stage_inst_dmem_n17470) );
NAND2_X1 MEM_stage_inst_dmem_U15704 ( .A1(MEM_stage_inst_dmem_ram_2371), .A2(MEM_stage_inst_dmem_n17476), .ZN(MEM_stage_inst_dmem_n17471) );
NAND2_X1 MEM_stage_inst_dmem_U15703 ( .A1(MEM_stage_inst_dmem_n17469), .A2(MEM_stage_inst_dmem_n17468), .ZN(MEM_stage_inst_dmem_n10623) );
NAND2_X1 MEM_stage_inst_dmem_U15702 ( .A1(EX_pipeline_reg_out_9), .A2(MEM_stage_inst_dmem_n17477), .ZN(MEM_stage_inst_dmem_n17468) );
NAND2_X1 MEM_stage_inst_dmem_U15701 ( .A1(MEM_stage_inst_dmem_ram_2372), .A2(MEM_stage_inst_dmem_n17476), .ZN(MEM_stage_inst_dmem_n17469) );
NAND2_X1 MEM_stage_inst_dmem_U15700 ( .A1(MEM_stage_inst_dmem_n17467), .A2(MEM_stage_inst_dmem_n17466), .ZN(MEM_stage_inst_dmem_n10624) );
NAND2_X1 MEM_stage_inst_dmem_U15699 ( .A1(EX_pipeline_reg_out_10), .A2(MEM_stage_inst_dmem_n17477), .ZN(MEM_stage_inst_dmem_n17466) );
NAND2_X1 MEM_stage_inst_dmem_U15698 ( .A1(MEM_stage_inst_dmem_ram_2373), .A2(MEM_stage_inst_dmem_n17476), .ZN(MEM_stage_inst_dmem_n17467) );
NAND2_X1 MEM_stage_inst_dmem_U15697 ( .A1(MEM_stage_inst_dmem_n17465), .A2(MEM_stage_inst_dmem_n17464), .ZN(MEM_stage_inst_dmem_n10625) );
NAND2_X1 MEM_stage_inst_dmem_U15696 ( .A1(EX_pipeline_reg_out_11), .A2(MEM_stage_inst_dmem_n17477), .ZN(MEM_stage_inst_dmem_n17464) );
NAND2_X1 MEM_stage_inst_dmem_U15695 ( .A1(MEM_stage_inst_dmem_ram_2374), .A2(MEM_stage_inst_dmem_n17476), .ZN(MEM_stage_inst_dmem_n17465) );
NAND2_X1 MEM_stage_inst_dmem_U15694 ( .A1(MEM_stage_inst_dmem_n17463), .A2(MEM_stage_inst_dmem_n17462), .ZN(MEM_stage_inst_dmem_n10626) );
NAND2_X1 MEM_stage_inst_dmem_U15693 ( .A1(EX_pipeline_reg_out_12), .A2(MEM_stage_inst_dmem_n17477), .ZN(MEM_stage_inst_dmem_n17462) );
NAND2_X1 MEM_stage_inst_dmem_U15692 ( .A1(MEM_stage_inst_dmem_ram_2375), .A2(MEM_stage_inst_dmem_n17476), .ZN(MEM_stage_inst_dmem_n17463) );
NAND2_X1 MEM_stage_inst_dmem_U15691 ( .A1(MEM_stage_inst_dmem_n17461), .A2(MEM_stage_inst_dmem_n17460), .ZN(MEM_stage_inst_dmem_n10627) );
NAND2_X1 MEM_stage_inst_dmem_U15690 ( .A1(EX_pipeline_reg_out_13), .A2(MEM_stage_inst_dmem_n17477), .ZN(MEM_stage_inst_dmem_n17460) );
NAND2_X1 MEM_stage_inst_dmem_U15689 ( .A1(MEM_stage_inst_dmem_ram_2376), .A2(MEM_stage_inst_dmem_n17476), .ZN(MEM_stage_inst_dmem_n17461) );
NAND2_X1 MEM_stage_inst_dmem_U15688 ( .A1(MEM_stage_inst_dmem_n17459), .A2(MEM_stage_inst_dmem_n17458), .ZN(MEM_stage_inst_dmem_n10628) );
NAND2_X1 MEM_stage_inst_dmem_U15687 ( .A1(EX_pipeline_reg_out_14), .A2(MEM_stage_inst_dmem_n17477), .ZN(MEM_stage_inst_dmem_n17458) );
NAND2_X1 MEM_stage_inst_dmem_U15686 ( .A1(MEM_stage_inst_dmem_ram_2377), .A2(MEM_stage_inst_dmem_n17476), .ZN(MEM_stage_inst_dmem_n17459) );
NAND2_X1 MEM_stage_inst_dmem_U15685 ( .A1(MEM_stage_inst_dmem_n17457), .A2(MEM_stage_inst_dmem_n17456), .ZN(MEM_stage_inst_dmem_n10629) );
NAND2_X1 MEM_stage_inst_dmem_U15684 ( .A1(EX_pipeline_reg_out_15), .A2(MEM_stage_inst_dmem_n17477), .ZN(MEM_stage_inst_dmem_n17456) );
NAND2_X1 MEM_stage_inst_dmem_U15683 ( .A1(MEM_stage_inst_dmem_ram_2378), .A2(MEM_stage_inst_dmem_n17476), .ZN(MEM_stage_inst_dmem_n17457) );
NAND2_X1 MEM_stage_inst_dmem_U15682 ( .A1(MEM_stage_inst_dmem_n17455), .A2(MEM_stage_inst_dmem_n17454), .ZN(MEM_stage_inst_dmem_n10630) );
NAND2_X1 MEM_stage_inst_dmem_U15681 ( .A1(EX_pipeline_reg_out_16), .A2(MEM_stage_inst_dmem_n17477), .ZN(MEM_stage_inst_dmem_n17454) );
NAND2_X1 MEM_stage_inst_dmem_U15680 ( .A1(MEM_stage_inst_dmem_ram_2379), .A2(MEM_stage_inst_dmem_n17476), .ZN(MEM_stage_inst_dmem_n17455) );
NAND2_X1 MEM_stage_inst_dmem_U15679 ( .A1(MEM_stage_inst_dmem_n17453), .A2(MEM_stage_inst_dmem_n17452), .ZN(MEM_stage_inst_dmem_n10631) );
NAND2_X1 MEM_stage_inst_dmem_U15678 ( .A1(EX_pipeline_reg_out_17), .A2(MEM_stage_inst_dmem_n17477), .ZN(MEM_stage_inst_dmem_n17452) );
NAND2_X1 MEM_stage_inst_dmem_U15677 ( .A1(MEM_stage_inst_dmem_ram_2380), .A2(MEM_stage_inst_dmem_n17476), .ZN(MEM_stage_inst_dmem_n17453) );
NAND2_X1 MEM_stage_inst_dmem_U15676 ( .A1(MEM_stage_inst_dmem_n17451), .A2(MEM_stage_inst_dmem_n17450), .ZN(MEM_stage_inst_dmem_n10632) );
NAND2_X1 MEM_stage_inst_dmem_U15675 ( .A1(EX_pipeline_reg_out_18), .A2(MEM_stage_inst_dmem_n17477), .ZN(MEM_stage_inst_dmem_n17450) );
NAND2_X1 MEM_stage_inst_dmem_U15674 ( .A1(MEM_stage_inst_dmem_ram_2381), .A2(MEM_stage_inst_dmem_n17476), .ZN(MEM_stage_inst_dmem_n17451) );
NAND2_X1 MEM_stage_inst_dmem_U15673 ( .A1(MEM_stage_inst_dmem_n17449), .A2(MEM_stage_inst_dmem_n17448), .ZN(MEM_stage_inst_dmem_n10633) );
NAND2_X1 MEM_stage_inst_dmem_U15672 ( .A1(EX_pipeline_reg_out_19), .A2(MEM_stage_inst_dmem_n17477), .ZN(MEM_stage_inst_dmem_n17448) );
NAND2_X1 MEM_stage_inst_dmem_U15671 ( .A1(MEM_stage_inst_dmem_ram_2382), .A2(MEM_stage_inst_dmem_n17476), .ZN(MEM_stage_inst_dmem_n17449) );
NAND2_X1 MEM_stage_inst_dmem_U15670 ( .A1(MEM_stage_inst_dmem_n17447), .A2(MEM_stage_inst_dmem_n17446), .ZN(MEM_stage_inst_dmem_n10634) );
NAND2_X1 MEM_stage_inst_dmem_U15669 ( .A1(EX_pipeline_reg_out_20), .A2(MEM_stage_inst_dmem_n17477), .ZN(MEM_stage_inst_dmem_n17446) );
INV_X1 MEM_stage_inst_dmem_U15668 ( .A(MEM_stage_inst_dmem_n17476), .ZN(MEM_stage_inst_dmem_n17477) );
NAND2_X1 MEM_stage_inst_dmem_U15667 ( .A1(MEM_stage_inst_dmem_ram_2383), .A2(MEM_stage_inst_dmem_n17476), .ZN(MEM_stage_inst_dmem_n17447) );
NAND2_X1 MEM_stage_inst_dmem_U15666 ( .A1(MEM_stage_inst_dmem_n21319), .A2(MEM_stage_inst_dmem_n17582), .ZN(MEM_stage_inst_dmem_n17476) );
NAND2_X1 MEM_stage_inst_dmem_U15665 ( .A1(MEM_stage_inst_dmem_n17445), .A2(MEM_stage_inst_dmem_n17444), .ZN(MEM_stage_inst_dmem_n10635) );
NAND2_X1 MEM_stage_inst_dmem_U15664 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n17443), .ZN(MEM_stage_inst_dmem_n17444) );
NAND2_X1 MEM_stage_inst_dmem_U15663 ( .A1(MEM_stage_inst_dmem_ram_2384), .A2(MEM_stage_inst_dmem_n17442), .ZN(MEM_stage_inst_dmem_n17445) );
NAND2_X1 MEM_stage_inst_dmem_U15662 ( .A1(MEM_stage_inst_dmem_n17441), .A2(MEM_stage_inst_dmem_n17440), .ZN(MEM_stage_inst_dmem_n10636) );
NAND2_X1 MEM_stage_inst_dmem_U15661 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n17443), .ZN(MEM_stage_inst_dmem_n17440) );
NAND2_X1 MEM_stage_inst_dmem_U15660 ( .A1(MEM_stage_inst_dmem_ram_2385), .A2(MEM_stage_inst_dmem_n17442), .ZN(MEM_stage_inst_dmem_n17441) );
NAND2_X1 MEM_stage_inst_dmem_U15659 ( .A1(MEM_stage_inst_dmem_n17439), .A2(MEM_stage_inst_dmem_n17438), .ZN(MEM_stage_inst_dmem_n10637) );
NAND2_X1 MEM_stage_inst_dmem_U15658 ( .A1(MEM_stage_inst_dmem_n18027), .A2(MEM_stage_inst_dmem_n17443), .ZN(MEM_stage_inst_dmem_n17438) );
NAND2_X1 MEM_stage_inst_dmem_U15657 ( .A1(MEM_stage_inst_dmem_ram_2386), .A2(MEM_stage_inst_dmem_n17442), .ZN(MEM_stage_inst_dmem_n17439) );
NAND2_X1 MEM_stage_inst_dmem_U15656 ( .A1(MEM_stage_inst_dmem_n17437), .A2(MEM_stage_inst_dmem_n17436), .ZN(MEM_stage_inst_dmem_n10638) );
NAND2_X1 MEM_stage_inst_dmem_U15655 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n17443), .ZN(MEM_stage_inst_dmem_n17436) );
NAND2_X1 MEM_stage_inst_dmem_U15654 ( .A1(MEM_stage_inst_dmem_ram_2387), .A2(MEM_stage_inst_dmem_n17442), .ZN(MEM_stage_inst_dmem_n17437) );
NAND2_X1 MEM_stage_inst_dmem_U15653 ( .A1(MEM_stage_inst_dmem_n17435), .A2(MEM_stage_inst_dmem_n17434), .ZN(MEM_stage_inst_dmem_n10639) );
NAND2_X1 MEM_stage_inst_dmem_U15652 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n17443), .ZN(MEM_stage_inst_dmem_n17434) );
NAND2_X1 MEM_stage_inst_dmem_U15651 ( .A1(MEM_stage_inst_dmem_ram_2388), .A2(MEM_stage_inst_dmem_n17442), .ZN(MEM_stage_inst_dmem_n17435) );
NAND2_X1 MEM_stage_inst_dmem_U15650 ( .A1(MEM_stage_inst_dmem_n17433), .A2(MEM_stage_inst_dmem_n17432), .ZN(MEM_stage_inst_dmem_n10640) );
NAND2_X1 MEM_stage_inst_dmem_U15649 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n17443), .ZN(MEM_stage_inst_dmem_n17432) );
NAND2_X1 MEM_stage_inst_dmem_U15648 ( .A1(MEM_stage_inst_dmem_ram_2389), .A2(MEM_stage_inst_dmem_n17442), .ZN(MEM_stage_inst_dmem_n17433) );
NAND2_X1 MEM_stage_inst_dmem_U15647 ( .A1(MEM_stage_inst_dmem_n17431), .A2(MEM_stage_inst_dmem_n17430), .ZN(MEM_stage_inst_dmem_n10641) );
NAND2_X1 MEM_stage_inst_dmem_U15646 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n17443), .ZN(MEM_stage_inst_dmem_n17430) );
NAND2_X1 MEM_stage_inst_dmem_U15645 ( .A1(MEM_stage_inst_dmem_ram_2390), .A2(MEM_stage_inst_dmem_n17442), .ZN(MEM_stage_inst_dmem_n17431) );
NAND2_X1 MEM_stage_inst_dmem_U15644 ( .A1(MEM_stage_inst_dmem_n17429), .A2(MEM_stage_inst_dmem_n17428), .ZN(MEM_stage_inst_dmem_n10642) );
NAND2_X1 MEM_stage_inst_dmem_U15643 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n17443), .ZN(MEM_stage_inst_dmem_n17428) );
NAND2_X1 MEM_stage_inst_dmem_U15642 ( .A1(MEM_stage_inst_dmem_ram_2391), .A2(MEM_stage_inst_dmem_n17442), .ZN(MEM_stage_inst_dmem_n17429) );
NAND2_X1 MEM_stage_inst_dmem_U15641 ( .A1(MEM_stage_inst_dmem_n17427), .A2(MEM_stage_inst_dmem_n17426), .ZN(MEM_stage_inst_dmem_n10643) );
NAND2_X1 MEM_stage_inst_dmem_U15640 ( .A1(MEM_stage_inst_dmem_n18013), .A2(MEM_stage_inst_dmem_n17443), .ZN(MEM_stage_inst_dmem_n17426) );
NAND2_X1 MEM_stage_inst_dmem_U15639 ( .A1(MEM_stage_inst_dmem_ram_2392), .A2(MEM_stage_inst_dmem_n17442), .ZN(MEM_stage_inst_dmem_n17427) );
NAND2_X1 MEM_stage_inst_dmem_U15638 ( .A1(MEM_stage_inst_dmem_n17425), .A2(MEM_stage_inst_dmem_n17424), .ZN(MEM_stage_inst_dmem_n10644) );
NAND2_X1 MEM_stage_inst_dmem_U15637 ( .A1(MEM_stage_inst_dmem_n96), .A2(MEM_stage_inst_dmem_n17443), .ZN(MEM_stage_inst_dmem_n17424) );
NAND2_X1 MEM_stage_inst_dmem_U15636 ( .A1(MEM_stage_inst_dmem_ram_2393), .A2(MEM_stage_inst_dmem_n17442), .ZN(MEM_stage_inst_dmem_n17425) );
NAND2_X1 MEM_stage_inst_dmem_U15635 ( .A1(MEM_stage_inst_dmem_n17423), .A2(MEM_stage_inst_dmem_n17422), .ZN(MEM_stage_inst_dmem_n10645) );
NAND2_X1 MEM_stage_inst_dmem_U15634 ( .A1(MEM_stage_inst_dmem_n18007), .A2(MEM_stage_inst_dmem_n17443), .ZN(MEM_stage_inst_dmem_n17422) );
NAND2_X1 MEM_stage_inst_dmem_U15633 ( .A1(MEM_stage_inst_dmem_ram_2394), .A2(MEM_stage_inst_dmem_n17442), .ZN(MEM_stage_inst_dmem_n17423) );
NAND2_X1 MEM_stage_inst_dmem_U15632 ( .A1(MEM_stage_inst_dmem_n17421), .A2(MEM_stage_inst_dmem_n17420), .ZN(MEM_stage_inst_dmem_n10646) );
NAND2_X1 MEM_stage_inst_dmem_U15631 ( .A1(MEM_stage_inst_dmem_n18004), .A2(MEM_stage_inst_dmem_n17443), .ZN(MEM_stage_inst_dmem_n17420) );
NAND2_X1 MEM_stage_inst_dmem_U15630 ( .A1(MEM_stage_inst_dmem_ram_2395), .A2(MEM_stage_inst_dmem_n17442), .ZN(MEM_stage_inst_dmem_n17421) );
NAND2_X1 MEM_stage_inst_dmem_U15629 ( .A1(MEM_stage_inst_dmem_n17419), .A2(MEM_stage_inst_dmem_n17418), .ZN(MEM_stage_inst_dmem_n10647) );
NAND2_X1 MEM_stage_inst_dmem_U15628 ( .A1(MEM_stage_inst_dmem_n18001), .A2(MEM_stage_inst_dmem_n17443), .ZN(MEM_stage_inst_dmem_n17418) );
NAND2_X1 MEM_stage_inst_dmem_U15627 ( .A1(MEM_stage_inst_dmem_ram_2396), .A2(MEM_stage_inst_dmem_n17442), .ZN(MEM_stage_inst_dmem_n17419) );
NAND2_X1 MEM_stage_inst_dmem_U15626 ( .A1(MEM_stage_inst_dmem_n17417), .A2(MEM_stage_inst_dmem_n17416), .ZN(MEM_stage_inst_dmem_n10648) );
NAND2_X1 MEM_stage_inst_dmem_U15625 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n17443), .ZN(MEM_stage_inst_dmem_n17416) );
NAND2_X1 MEM_stage_inst_dmem_U15624 ( .A1(MEM_stage_inst_dmem_ram_2397), .A2(MEM_stage_inst_dmem_n17442), .ZN(MEM_stage_inst_dmem_n17417) );
NAND2_X1 MEM_stage_inst_dmem_U15623 ( .A1(MEM_stage_inst_dmem_n17415), .A2(MEM_stage_inst_dmem_n17414), .ZN(MEM_stage_inst_dmem_n10649) );
NAND2_X1 MEM_stage_inst_dmem_U15622 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n17443), .ZN(MEM_stage_inst_dmem_n17414) );
NAND2_X1 MEM_stage_inst_dmem_U15621 ( .A1(MEM_stage_inst_dmem_ram_2398), .A2(MEM_stage_inst_dmem_n17442), .ZN(MEM_stage_inst_dmem_n17415) );
NAND2_X1 MEM_stage_inst_dmem_U15620 ( .A1(MEM_stage_inst_dmem_n17413), .A2(MEM_stage_inst_dmem_n17412), .ZN(MEM_stage_inst_dmem_n10650) );
NAND2_X1 MEM_stage_inst_dmem_U15619 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n17443), .ZN(MEM_stage_inst_dmem_n17412) );
INV_X1 MEM_stage_inst_dmem_U15618 ( .A(MEM_stage_inst_dmem_n17442), .ZN(MEM_stage_inst_dmem_n17443) );
NAND2_X1 MEM_stage_inst_dmem_U15617 ( .A1(MEM_stage_inst_dmem_ram_2399), .A2(MEM_stage_inst_dmem_n17442), .ZN(MEM_stage_inst_dmem_n17413) );
NAND2_X1 MEM_stage_inst_dmem_U15616 ( .A1(MEM_stage_inst_dmem_n21284), .A2(MEM_stage_inst_dmem_n17582), .ZN(MEM_stage_inst_dmem_n17442) );
NAND2_X1 MEM_stage_inst_dmem_U15615 ( .A1(MEM_stage_inst_dmem_n17411), .A2(MEM_stage_inst_dmem_n17410), .ZN(MEM_stage_inst_dmem_n10651) );
NAND2_X1 MEM_stage_inst_dmem_U15614 ( .A1(EX_pipeline_reg_out_5), .A2(MEM_stage_inst_dmem_n17409), .ZN(MEM_stage_inst_dmem_n17410) );
NAND2_X1 MEM_stage_inst_dmem_U15613 ( .A1(MEM_stage_inst_dmem_ram_2400), .A2(MEM_stage_inst_dmem_n17408), .ZN(MEM_stage_inst_dmem_n17411) );
NAND2_X1 MEM_stage_inst_dmem_U15612 ( .A1(MEM_stage_inst_dmem_n17407), .A2(MEM_stage_inst_dmem_n17406), .ZN(MEM_stage_inst_dmem_n10652) );
NAND2_X1 MEM_stage_inst_dmem_U15611 ( .A1(EX_pipeline_reg_out_6), .A2(MEM_stage_inst_dmem_n17409), .ZN(MEM_stage_inst_dmem_n17406) );
NAND2_X1 MEM_stage_inst_dmem_U15610 ( .A1(MEM_stage_inst_dmem_ram_2401), .A2(MEM_stage_inst_dmem_n17408), .ZN(MEM_stage_inst_dmem_n17407) );
NAND2_X1 MEM_stage_inst_dmem_U15609 ( .A1(MEM_stage_inst_dmem_n17405), .A2(MEM_stage_inst_dmem_n17404), .ZN(MEM_stage_inst_dmem_n10653) );
NAND2_X1 MEM_stage_inst_dmem_U15608 ( .A1(EX_pipeline_reg_out_7), .A2(MEM_stage_inst_dmem_n17409), .ZN(MEM_stage_inst_dmem_n17404) );
NAND2_X1 MEM_stage_inst_dmem_U15607 ( .A1(MEM_stage_inst_dmem_ram_2402), .A2(MEM_stage_inst_dmem_n17408), .ZN(MEM_stage_inst_dmem_n17405) );
NAND2_X1 MEM_stage_inst_dmem_U15606 ( .A1(MEM_stage_inst_dmem_n17403), .A2(MEM_stage_inst_dmem_n17402), .ZN(MEM_stage_inst_dmem_n10654) );
NAND2_X1 MEM_stage_inst_dmem_U15605 ( .A1(EX_pipeline_reg_out_8), .A2(MEM_stage_inst_dmem_n17409), .ZN(MEM_stage_inst_dmem_n17402) );
NAND2_X1 MEM_stage_inst_dmem_U15604 ( .A1(MEM_stage_inst_dmem_ram_2403), .A2(MEM_stage_inst_dmem_n17408), .ZN(MEM_stage_inst_dmem_n17403) );
NAND2_X1 MEM_stage_inst_dmem_U15603 ( .A1(MEM_stage_inst_dmem_n17401), .A2(MEM_stage_inst_dmem_n17400), .ZN(MEM_stage_inst_dmem_n10655) );
NAND2_X1 MEM_stage_inst_dmem_U15602 ( .A1(EX_pipeline_reg_out_9), .A2(MEM_stage_inst_dmem_n17409), .ZN(MEM_stage_inst_dmem_n17400) );
NAND2_X1 MEM_stage_inst_dmem_U15601 ( .A1(MEM_stage_inst_dmem_ram_2404), .A2(MEM_stage_inst_dmem_n17408), .ZN(MEM_stage_inst_dmem_n17401) );
NAND2_X1 MEM_stage_inst_dmem_U15600 ( .A1(MEM_stage_inst_dmem_n17399), .A2(MEM_stage_inst_dmem_n17398), .ZN(MEM_stage_inst_dmem_n10656) );
NAND2_X1 MEM_stage_inst_dmem_U15599 ( .A1(EX_pipeline_reg_out_10), .A2(MEM_stage_inst_dmem_n17409), .ZN(MEM_stage_inst_dmem_n17398) );
NAND2_X1 MEM_stage_inst_dmem_U15598 ( .A1(MEM_stage_inst_dmem_ram_2405), .A2(MEM_stage_inst_dmem_n17408), .ZN(MEM_stage_inst_dmem_n17399) );
NAND2_X1 MEM_stage_inst_dmem_U15597 ( .A1(MEM_stage_inst_dmem_n17397), .A2(MEM_stage_inst_dmem_n17396), .ZN(MEM_stage_inst_dmem_n10657) );
NAND2_X1 MEM_stage_inst_dmem_U15596 ( .A1(EX_pipeline_reg_out_11), .A2(MEM_stage_inst_dmem_n17409), .ZN(MEM_stage_inst_dmem_n17396) );
NAND2_X1 MEM_stage_inst_dmem_U15595 ( .A1(MEM_stage_inst_dmem_ram_2406), .A2(MEM_stage_inst_dmem_n17408), .ZN(MEM_stage_inst_dmem_n17397) );
NAND2_X1 MEM_stage_inst_dmem_U15594 ( .A1(MEM_stage_inst_dmem_n17395), .A2(MEM_stage_inst_dmem_n17394), .ZN(MEM_stage_inst_dmem_n10658) );
NAND2_X1 MEM_stage_inst_dmem_U15593 ( .A1(EX_pipeline_reg_out_12), .A2(MEM_stage_inst_dmem_n17409), .ZN(MEM_stage_inst_dmem_n17394) );
NAND2_X1 MEM_stage_inst_dmem_U15592 ( .A1(MEM_stage_inst_dmem_ram_2407), .A2(MEM_stage_inst_dmem_n17408), .ZN(MEM_stage_inst_dmem_n17395) );
NAND2_X1 MEM_stage_inst_dmem_U15591 ( .A1(MEM_stage_inst_dmem_n17393), .A2(MEM_stage_inst_dmem_n17392), .ZN(MEM_stage_inst_dmem_n10659) );
NAND2_X1 MEM_stage_inst_dmem_U15590 ( .A1(EX_pipeline_reg_out_13), .A2(MEM_stage_inst_dmem_n17409), .ZN(MEM_stage_inst_dmem_n17392) );
NAND2_X1 MEM_stage_inst_dmem_U15589 ( .A1(MEM_stage_inst_dmem_ram_2408), .A2(MEM_stage_inst_dmem_n17408), .ZN(MEM_stage_inst_dmem_n17393) );
NAND2_X1 MEM_stage_inst_dmem_U15588 ( .A1(MEM_stage_inst_dmem_n17391), .A2(MEM_stage_inst_dmem_n17390), .ZN(MEM_stage_inst_dmem_n10660) );
NAND2_X1 MEM_stage_inst_dmem_U15587 ( .A1(EX_pipeline_reg_out_14), .A2(MEM_stage_inst_dmem_n17409), .ZN(MEM_stage_inst_dmem_n17390) );
NAND2_X1 MEM_stage_inst_dmem_U15586 ( .A1(MEM_stage_inst_dmem_ram_2409), .A2(MEM_stage_inst_dmem_n17408), .ZN(MEM_stage_inst_dmem_n17391) );
NAND2_X1 MEM_stage_inst_dmem_U15585 ( .A1(MEM_stage_inst_dmem_n17389), .A2(MEM_stage_inst_dmem_n17388), .ZN(MEM_stage_inst_dmem_n10661) );
NAND2_X1 MEM_stage_inst_dmem_U15584 ( .A1(EX_pipeline_reg_out_15), .A2(MEM_stage_inst_dmem_n17409), .ZN(MEM_stage_inst_dmem_n17388) );
NAND2_X1 MEM_stage_inst_dmem_U15583 ( .A1(MEM_stage_inst_dmem_ram_2410), .A2(MEM_stage_inst_dmem_n17408), .ZN(MEM_stage_inst_dmem_n17389) );
NAND2_X1 MEM_stage_inst_dmem_U15582 ( .A1(MEM_stage_inst_dmem_n17387), .A2(MEM_stage_inst_dmem_n17386), .ZN(MEM_stage_inst_dmem_n10662) );
NAND2_X1 MEM_stage_inst_dmem_U15581 ( .A1(EX_pipeline_reg_out_16), .A2(MEM_stage_inst_dmem_n17409), .ZN(MEM_stage_inst_dmem_n17386) );
NAND2_X1 MEM_stage_inst_dmem_U15580 ( .A1(MEM_stage_inst_dmem_ram_2411), .A2(MEM_stage_inst_dmem_n17408), .ZN(MEM_stage_inst_dmem_n17387) );
NAND2_X1 MEM_stage_inst_dmem_U15579 ( .A1(MEM_stage_inst_dmem_n17385), .A2(MEM_stage_inst_dmem_n17384), .ZN(MEM_stage_inst_dmem_n10663) );
NAND2_X1 MEM_stage_inst_dmem_U15578 ( .A1(EX_pipeline_reg_out_17), .A2(MEM_stage_inst_dmem_n17409), .ZN(MEM_stage_inst_dmem_n17384) );
NAND2_X1 MEM_stage_inst_dmem_U15577 ( .A1(MEM_stage_inst_dmem_ram_2412), .A2(MEM_stage_inst_dmem_n17408), .ZN(MEM_stage_inst_dmem_n17385) );
NAND2_X1 MEM_stage_inst_dmem_U15576 ( .A1(MEM_stage_inst_dmem_n17383), .A2(MEM_stage_inst_dmem_n17382), .ZN(MEM_stage_inst_dmem_n10664) );
NAND2_X1 MEM_stage_inst_dmem_U15575 ( .A1(EX_pipeline_reg_out_18), .A2(MEM_stage_inst_dmem_n17409), .ZN(MEM_stage_inst_dmem_n17382) );
NAND2_X1 MEM_stage_inst_dmem_U15574 ( .A1(MEM_stage_inst_dmem_ram_2413), .A2(MEM_stage_inst_dmem_n17408), .ZN(MEM_stage_inst_dmem_n17383) );
NAND2_X1 MEM_stage_inst_dmem_U15573 ( .A1(MEM_stage_inst_dmem_n17381), .A2(MEM_stage_inst_dmem_n17380), .ZN(MEM_stage_inst_dmem_n10665) );
NAND2_X1 MEM_stage_inst_dmem_U15572 ( .A1(EX_pipeline_reg_out_19), .A2(MEM_stage_inst_dmem_n17409), .ZN(MEM_stage_inst_dmem_n17380) );
NAND2_X1 MEM_stage_inst_dmem_U15571 ( .A1(MEM_stage_inst_dmem_ram_2414), .A2(MEM_stage_inst_dmem_n17408), .ZN(MEM_stage_inst_dmem_n17381) );
NAND2_X1 MEM_stage_inst_dmem_U15570 ( .A1(MEM_stage_inst_dmem_n17379), .A2(MEM_stage_inst_dmem_n17378), .ZN(MEM_stage_inst_dmem_n10666) );
NAND2_X1 MEM_stage_inst_dmem_U15569 ( .A1(EX_pipeline_reg_out_20), .A2(MEM_stage_inst_dmem_n17409), .ZN(MEM_stage_inst_dmem_n17378) );
INV_X1 MEM_stage_inst_dmem_U15568 ( .A(MEM_stage_inst_dmem_n17408), .ZN(MEM_stage_inst_dmem_n17409) );
NAND2_X1 MEM_stage_inst_dmem_U15567 ( .A1(MEM_stage_inst_dmem_ram_2415), .A2(MEM_stage_inst_dmem_n17408), .ZN(MEM_stage_inst_dmem_n17379) );
NAND2_X1 MEM_stage_inst_dmem_U15566 ( .A1(MEM_stage_inst_dmem_n21249), .A2(MEM_stage_inst_dmem_n17582), .ZN(MEM_stage_inst_dmem_n17408) );
NAND2_X1 MEM_stage_inst_dmem_U15565 ( .A1(MEM_stage_inst_dmem_n17377), .A2(MEM_stage_inst_dmem_n17376), .ZN(MEM_stage_inst_dmem_n10667) );
NAND2_X1 MEM_stage_inst_dmem_U15564 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n17375), .ZN(MEM_stage_inst_dmem_n17376) );
NAND2_X1 MEM_stage_inst_dmem_U15563 ( .A1(MEM_stage_inst_dmem_ram_2416), .A2(MEM_stage_inst_dmem_n17374), .ZN(MEM_stage_inst_dmem_n17377) );
NAND2_X1 MEM_stage_inst_dmem_U15562 ( .A1(MEM_stage_inst_dmem_n17373), .A2(MEM_stage_inst_dmem_n17372), .ZN(MEM_stage_inst_dmem_n10668) );
NAND2_X1 MEM_stage_inst_dmem_U15561 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n17375), .ZN(MEM_stage_inst_dmem_n17372) );
NAND2_X1 MEM_stage_inst_dmem_U15560 ( .A1(MEM_stage_inst_dmem_ram_2417), .A2(MEM_stage_inst_dmem_n17374), .ZN(MEM_stage_inst_dmem_n17373) );
NAND2_X1 MEM_stage_inst_dmem_U15559 ( .A1(MEM_stage_inst_dmem_n17371), .A2(MEM_stage_inst_dmem_n17370), .ZN(MEM_stage_inst_dmem_n10669) );
NAND2_X1 MEM_stage_inst_dmem_U15558 ( .A1(MEM_stage_inst_dmem_n18027), .A2(MEM_stage_inst_dmem_n17375), .ZN(MEM_stage_inst_dmem_n17370) );
NAND2_X1 MEM_stage_inst_dmem_U15557 ( .A1(MEM_stage_inst_dmem_ram_2418), .A2(MEM_stage_inst_dmem_n17374), .ZN(MEM_stage_inst_dmem_n17371) );
NAND2_X1 MEM_stage_inst_dmem_U15556 ( .A1(MEM_stage_inst_dmem_n17369), .A2(MEM_stage_inst_dmem_n17368), .ZN(MEM_stage_inst_dmem_n10670) );
NAND2_X1 MEM_stage_inst_dmem_U15555 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n17375), .ZN(MEM_stage_inst_dmem_n17368) );
NAND2_X1 MEM_stage_inst_dmem_U15554 ( .A1(MEM_stage_inst_dmem_ram_2419), .A2(MEM_stage_inst_dmem_n17374), .ZN(MEM_stage_inst_dmem_n17369) );
NAND2_X1 MEM_stage_inst_dmem_U15553 ( .A1(MEM_stage_inst_dmem_n17367), .A2(MEM_stage_inst_dmem_n17366), .ZN(MEM_stage_inst_dmem_n10671) );
NAND2_X1 MEM_stage_inst_dmem_U15552 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n17375), .ZN(MEM_stage_inst_dmem_n17366) );
NAND2_X1 MEM_stage_inst_dmem_U15551 ( .A1(MEM_stage_inst_dmem_ram_2420), .A2(MEM_stage_inst_dmem_n17374), .ZN(MEM_stage_inst_dmem_n17367) );
NAND2_X1 MEM_stage_inst_dmem_U15550 ( .A1(MEM_stage_inst_dmem_n17365), .A2(MEM_stage_inst_dmem_n17364), .ZN(MEM_stage_inst_dmem_n10672) );
NAND2_X1 MEM_stage_inst_dmem_U15549 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n17375), .ZN(MEM_stage_inst_dmem_n17364) );
NAND2_X1 MEM_stage_inst_dmem_U15548 ( .A1(MEM_stage_inst_dmem_ram_2421), .A2(MEM_stage_inst_dmem_n17374), .ZN(MEM_stage_inst_dmem_n17365) );
NAND2_X1 MEM_stage_inst_dmem_U15547 ( .A1(MEM_stage_inst_dmem_n17363), .A2(MEM_stage_inst_dmem_n17362), .ZN(MEM_stage_inst_dmem_n10673) );
NAND2_X1 MEM_stage_inst_dmem_U15546 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n17375), .ZN(MEM_stage_inst_dmem_n17362) );
NAND2_X1 MEM_stage_inst_dmem_U15545 ( .A1(MEM_stage_inst_dmem_ram_2422), .A2(MEM_stage_inst_dmem_n17374), .ZN(MEM_stage_inst_dmem_n17363) );
NAND2_X1 MEM_stage_inst_dmem_U15544 ( .A1(MEM_stage_inst_dmem_n17361), .A2(MEM_stage_inst_dmem_n17360), .ZN(MEM_stage_inst_dmem_n10674) );
NAND2_X1 MEM_stage_inst_dmem_U15543 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n17375), .ZN(MEM_stage_inst_dmem_n17360) );
NAND2_X1 MEM_stage_inst_dmem_U15542 ( .A1(MEM_stage_inst_dmem_ram_2423), .A2(MEM_stage_inst_dmem_n17374), .ZN(MEM_stage_inst_dmem_n17361) );
NAND2_X1 MEM_stage_inst_dmem_U15541 ( .A1(MEM_stage_inst_dmem_n17359), .A2(MEM_stage_inst_dmem_n17358), .ZN(MEM_stage_inst_dmem_n10675) );
NAND2_X1 MEM_stage_inst_dmem_U15540 ( .A1(MEM_stage_inst_dmem_n18013), .A2(MEM_stage_inst_dmem_n17375), .ZN(MEM_stage_inst_dmem_n17358) );
NAND2_X1 MEM_stage_inst_dmem_U15539 ( .A1(MEM_stage_inst_dmem_ram_2424), .A2(MEM_stage_inst_dmem_n17374), .ZN(MEM_stage_inst_dmem_n17359) );
NAND2_X1 MEM_stage_inst_dmem_U15538 ( .A1(MEM_stage_inst_dmem_n17357), .A2(MEM_stage_inst_dmem_n17356), .ZN(MEM_stage_inst_dmem_n10676) );
NAND2_X1 MEM_stage_inst_dmem_U15537 ( .A1(MEM_stage_inst_dmem_n96), .A2(MEM_stage_inst_dmem_n17375), .ZN(MEM_stage_inst_dmem_n17356) );
NAND2_X1 MEM_stage_inst_dmem_U15536 ( .A1(MEM_stage_inst_dmem_ram_2425), .A2(MEM_stage_inst_dmem_n17374), .ZN(MEM_stage_inst_dmem_n17357) );
NAND2_X1 MEM_stage_inst_dmem_U15535 ( .A1(MEM_stage_inst_dmem_n17355), .A2(MEM_stage_inst_dmem_n17354), .ZN(MEM_stage_inst_dmem_n10677) );
NAND2_X1 MEM_stage_inst_dmem_U15534 ( .A1(MEM_stage_inst_dmem_n18007), .A2(MEM_stage_inst_dmem_n17375), .ZN(MEM_stage_inst_dmem_n17354) );
NAND2_X1 MEM_stage_inst_dmem_U15533 ( .A1(MEM_stage_inst_dmem_ram_2426), .A2(MEM_stage_inst_dmem_n17374), .ZN(MEM_stage_inst_dmem_n17355) );
NAND2_X1 MEM_stage_inst_dmem_U15532 ( .A1(MEM_stage_inst_dmem_n17353), .A2(MEM_stage_inst_dmem_n17352), .ZN(MEM_stage_inst_dmem_n10678) );
NAND2_X1 MEM_stage_inst_dmem_U15531 ( .A1(MEM_stage_inst_dmem_n18004), .A2(MEM_stage_inst_dmem_n17375), .ZN(MEM_stage_inst_dmem_n17352) );
NAND2_X1 MEM_stage_inst_dmem_U15530 ( .A1(MEM_stage_inst_dmem_ram_2427), .A2(MEM_stage_inst_dmem_n17374), .ZN(MEM_stage_inst_dmem_n17353) );
NAND2_X1 MEM_stage_inst_dmem_U15529 ( .A1(MEM_stage_inst_dmem_n17351), .A2(MEM_stage_inst_dmem_n17350), .ZN(MEM_stage_inst_dmem_n10679) );
NAND2_X1 MEM_stage_inst_dmem_U15528 ( .A1(MEM_stage_inst_dmem_n18001), .A2(MEM_stage_inst_dmem_n17375), .ZN(MEM_stage_inst_dmem_n17350) );
NAND2_X1 MEM_stage_inst_dmem_U15527 ( .A1(MEM_stage_inst_dmem_ram_2428), .A2(MEM_stage_inst_dmem_n17374), .ZN(MEM_stage_inst_dmem_n17351) );
NAND2_X1 MEM_stage_inst_dmem_U15526 ( .A1(MEM_stage_inst_dmem_n17349), .A2(MEM_stage_inst_dmem_n17348), .ZN(MEM_stage_inst_dmem_n10680) );
NAND2_X1 MEM_stage_inst_dmem_U15525 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n17375), .ZN(MEM_stage_inst_dmem_n17348) );
NAND2_X1 MEM_stage_inst_dmem_U15524 ( .A1(MEM_stage_inst_dmem_ram_2429), .A2(MEM_stage_inst_dmem_n17374), .ZN(MEM_stage_inst_dmem_n17349) );
NAND2_X1 MEM_stage_inst_dmem_U15523 ( .A1(MEM_stage_inst_dmem_n17347), .A2(MEM_stage_inst_dmem_n17346), .ZN(MEM_stage_inst_dmem_n10681) );
NAND2_X1 MEM_stage_inst_dmem_U15522 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n17375), .ZN(MEM_stage_inst_dmem_n17346) );
NAND2_X1 MEM_stage_inst_dmem_U15521 ( .A1(MEM_stage_inst_dmem_ram_2430), .A2(MEM_stage_inst_dmem_n17374), .ZN(MEM_stage_inst_dmem_n17347) );
NAND2_X1 MEM_stage_inst_dmem_U15520 ( .A1(MEM_stage_inst_dmem_n17345), .A2(MEM_stage_inst_dmem_n17344), .ZN(MEM_stage_inst_dmem_n10682) );
NAND2_X1 MEM_stage_inst_dmem_U15519 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n17375), .ZN(MEM_stage_inst_dmem_n17344) );
NAND2_X1 MEM_stage_inst_dmem_U15518 ( .A1(MEM_stage_inst_dmem_ram_2431), .A2(MEM_stage_inst_dmem_n17374), .ZN(MEM_stage_inst_dmem_n17345) );
NAND2_X1 MEM_stage_inst_dmem_U15517 ( .A1(MEM_stage_inst_dmem_n21214), .A2(MEM_stage_inst_dmem_n17582), .ZN(MEM_stage_inst_dmem_n17374) );
NAND2_X1 MEM_stage_inst_dmem_U15516 ( .A1(MEM_stage_inst_dmem_n17343), .A2(MEM_stage_inst_dmem_n17342), .ZN(MEM_stage_inst_dmem_n10683) );
NAND2_X1 MEM_stage_inst_dmem_U15515 ( .A1(EX_pipeline_reg_out_5), .A2(MEM_stage_inst_dmem_n17341), .ZN(MEM_stage_inst_dmem_n17342) );
NAND2_X1 MEM_stage_inst_dmem_U15514 ( .A1(MEM_stage_inst_dmem_ram_2432), .A2(MEM_stage_inst_dmem_n17340), .ZN(MEM_stage_inst_dmem_n17343) );
NAND2_X1 MEM_stage_inst_dmem_U15513 ( .A1(MEM_stage_inst_dmem_n17339), .A2(MEM_stage_inst_dmem_n17338), .ZN(MEM_stage_inst_dmem_n10684) );
NAND2_X1 MEM_stage_inst_dmem_U15512 ( .A1(EX_pipeline_reg_out_6), .A2(MEM_stage_inst_dmem_n17341), .ZN(MEM_stage_inst_dmem_n17338) );
NAND2_X1 MEM_stage_inst_dmem_U15511 ( .A1(MEM_stage_inst_dmem_ram_2433), .A2(MEM_stage_inst_dmem_n17340), .ZN(MEM_stage_inst_dmem_n17339) );
NAND2_X1 MEM_stage_inst_dmem_U15510 ( .A1(MEM_stage_inst_dmem_n17337), .A2(MEM_stage_inst_dmem_n17336), .ZN(MEM_stage_inst_dmem_n10685) );
NAND2_X1 MEM_stage_inst_dmem_U15509 ( .A1(EX_pipeline_reg_out_7), .A2(MEM_stage_inst_dmem_n17341), .ZN(MEM_stage_inst_dmem_n17336) );
NAND2_X1 MEM_stage_inst_dmem_U15508 ( .A1(MEM_stage_inst_dmem_ram_2434), .A2(MEM_stage_inst_dmem_n17340), .ZN(MEM_stage_inst_dmem_n17337) );
NAND2_X1 MEM_stage_inst_dmem_U15507 ( .A1(MEM_stage_inst_dmem_n17335), .A2(MEM_stage_inst_dmem_n17334), .ZN(MEM_stage_inst_dmem_n10686) );
NAND2_X1 MEM_stage_inst_dmem_U15506 ( .A1(EX_pipeline_reg_out_8), .A2(MEM_stage_inst_dmem_n17341), .ZN(MEM_stage_inst_dmem_n17334) );
NAND2_X1 MEM_stage_inst_dmem_U15505 ( .A1(MEM_stage_inst_dmem_ram_2435), .A2(MEM_stage_inst_dmem_n17340), .ZN(MEM_stage_inst_dmem_n17335) );
NAND2_X1 MEM_stage_inst_dmem_U15504 ( .A1(MEM_stage_inst_dmem_n17333), .A2(MEM_stage_inst_dmem_n17332), .ZN(MEM_stage_inst_dmem_n10687) );
NAND2_X1 MEM_stage_inst_dmem_U15503 ( .A1(EX_pipeline_reg_out_9), .A2(MEM_stage_inst_dmem_n17341), .ZN(MEM_stage_inst_dmem_n17332) );
NAND2_X1 MEM_stage_inst_dmem_U15502 ( .A1(MEM_stage_inst_dmem_ram_2436), .A2(MEM_stage_inst_dmem_n17340), .ZN(MEM_stage_inst_dmem_n17333) );
NAND2_X1 MEM_stage_inst_dmem_U15501 ( .A1(MEM_stage_inst_dmem_n17331), .A2(MEM_stage_inst_dmem_n17330), .ZN(MEM_stage_inst_dmem_n10688) );
NAND2_X1 MEM_stage_inst_dmem_U15500 ( .A1(EX_pipeline_reg_out_10), .A2(MEM_stage_inst_dmem_n17341), .ZN(MEM_stage_inst_dmem_n17330) );
NAND2_X1 MEM_stage_inst_dmem_U15499 ( .A1(MEM_stage_inst_dmem_ram_2437), .A2(MEM_stage_inst_dmem_n17340), .ZN(MEM_stage_inst_dmem_n17331) );
NAND2_X1 MEM_stage_inst_dmem_U15498 ( .A1(MEM_stage_inst_dmem_n17329), .A2(MEM_stage_inst_dmem_n17328), .ZN(MEM_stage_inst_dmem_n10689) );
NAND2_X1 MEM_stage_inst_dmem_U15497 ( .A1(EX_pipeline_reg_out_11), .A2(MEM_stage_inst_dmem_n17341), .ZN(MEM_stage_inst_dmem_n17328) );
NAND2_X1 MEM_stage_inst_dmem_U15496 ( .A1(MEM_stage_inst_dmem_ram_2438), .A2(MEM_stage_inst_dmem_n17340), .ZN(MEM_stage_inst_dmem_n17329) );
NAND2_X1 MEM_stage_inst_dmem_U15495 ( .A1(MEM_stage_inst_dmem_n17327), .A2(MEM_stage_inst_dmem_n17326), .ZN(MEM_stage_inst_dmem_n10690) );
NAND2_X1 MEM_stage_inst_dmem_U15494 ( .A1(EX_pipeline_reg_out_12), .A2(MEM_stage_inst_dmem_n17341), .ZN(MEM_stage_inst_dmem_n17326) );
NAND2_X1 MEM_stage_inst_dmem_U15493 ( .A1(MEM_stage_inst_dmem_ram_2439), .A2(MEM_stage_inst_dmem_n17340), .ZN(MEM_stage_inst_dmem_n17327) );
NAND2_X1 MEM_stage_inst_dmem_U15492 ( .A1(MEM_stage_inst_dmem_n17325), .A2(MEM_stage_inst_dmem_n17324), .ZN(MEM_stage_inst_dmem_n10691) );
NAND2_X1 MEM_stage_inst_dmem_U15491 ( .A1(EX_pipeline_reg_out_13), .A2(MEM_stage_inst_dmem_n17341), .ZN(MEM_stage_inst_dmem_n17324) );
NAND2_X1 MEM_stage_inst_dmem_U15490 ( .A1(MEM_stage_inst_dmem_ram_2440), .A2(MEM_stage_inst_dmem_n17340), .ZN(MEM_stage_inst_dmem_n17325) );
NAND2_X1 MEM_stage_inst_dmem_U15489 ( .A1(MEM_stage_inst_dmem_n17323), .A2(MEM_stage_inst_dmem_n17322), .ZN(MEM_stage_inst_dmem_n10692) );
NAND2_X1 MEM_stage_inst_dmem_U15488 ( .A1(EX_pipeline_reg_out_14), .A2(MEM_stage_inst_dmem_n17341), .ZN(MEM_stage_inst_dmem_n17322) );
NAND2_X1 MEM_stage_inst_dmem_U15487 ( .A1(MEM_stage_inst_dmem_ram_2441), .A2(MEM_stage_inst_dmem_n17340), .ZN(MEM_stage_inst_dmem_n17323) );
NAND2_X1 MEM_stage_inst_dmem_U15486 ( .A1(MEM_stage_inst_dmem_n17321), .A2(MEM_stage_inst_dmem_n17320), .ZN(MEM_stage_inst_dmem_n10693) );
NAND2_X1 MEM_stage_inst_dmem_U15485 ( .A1(EX_pipeline_reg_out_15), .A2(MEM_stage_inst_dmem_n17341), .ZN(MEM_stage_inst_dmem_n17320) );
NAND2_X1 MEM_stage_inst_dmem_U15484 ( .A1(MEM_stage_inst_dmem_ram_2442), .A2(MEM_stage_inst_dmem_n17340), .ZN(MEM_stage_inst_dmem_n17321) );
NAND2_X1 MEM_stage_inst_dmem_U15483 ( .A1(MEM_stage_inst_dmem_n17319), .A2(MEM_stage_inst_dmem_n17318), .ZN(MEM_stage_inst_dmem_n10694) );
NAND2_X1 MEM_stage_inst_dmem_U15482 ( .A1(EX_pipeline_reg_out_16), .A2(MEM_stage_inst_dmem_n17341), .ZN(MEM_stage_inst_dmem_n17318) );
NAND2_X1 MEM_stage_inst_dmem_U15481 ( .A1(MEM_stage_inst_dmem_ram_2443), .A2(MEM_stage_inst_dmem_n17340), .ZN(MEM_stage_inst_dmem_n17319) );
NAND2_X1 MEM_stage_inst_dmem_U15480 ( .A1(MEM_stage_inst_dmem_n17317), .A2(MEM_stage_inst_dmem_n17316), .ZN(MEM_stage_inst_dmem_n10695) );
NAND2_X1 MEM_stage_inst_dmem_U15479 ( .A1(EX_pipeline_reg_out_17), .A2(MEM_stage_inst_dmem_n17341), .ZN(MEM_stage_inst_dmem_n17316) );
NAND2_X1 MEM_stage_inst_dmem_U15478 ( .A1(MEM_stage_inst_dmem_ram_2444), .A2(MEM_stage_inst_dmem_n17340), .ZN(MEM_stage_inst_dmem_n17317) );
NAND2_X1 MEM_stage_inst_dmem_U15477 ( .A1(MEM_stage_inst_dmem_n17315), .A2(MEM_stage_inst_dmem_n17314), .ZN(MEM_stage_inst_dmem_n10696) );
NAND2_X1 MEM_stage_inst_dmem_U15476 ( .A1(EX_pipeline_reg_out_18), .A2(MEM_stage_inst_dmem_n17341), .ZN(MEM_stage_inst_dmem_n17314) );
NAND2_X1 MEM_stage_inst_dmem_U15475 ( .A1(MEM_stage_inst_dmem_ram_2445), .A2(MEM_stage_inst_dmem_n17340), .ZN(MEM_stage_inst_dmem_n17315) );
NAND2_X1 MEM_stage_inst_dmem_U15474 ( .A1(MEM_stage_inst_dmem_n17313), .A2(MEM_stage_inst_dmem_n17312), .ZN(MEM_stage_inst_dmem_n10697) );
NAND2_X1 MEM_stage_inst_dmem_U15473 ( .A1(EX_pipeline_reg_out_19), .A2(MEM_stage_inst_dmem_n17341), .ZN(MEM_stage_inst_dmem_n17312) );
NAND2_X1 MEM_stage_inst_dmem_U15472 ( .A1(MEM_stage_inst_dmem_ram_2446), .A2(MEM_stage_inst_dmem_n17340), .ZN(MEM_stage_inst_dmem_n17313) );
NAND2_X1 MEM_stage_inst_dmem_U15471 ( .A1(MEM_stage_inst_dmem_n17311), .A2(MEM_stage_inst_dmem_n17310), .ZN(MEM_stage_inst_dmem_n10698) );
NAND2_X1 MEM_stage_inst_dmem_U15470 ( .A1(EX_pipeline_reg_out_20), .A2(MEM_stage_inst_dmem_n17341), .ZN(MEM_stage_inst_dmem_n17310) );
INV_X1 MEM_stage_inst_dmem_U15469 ( .A(MEM_stage_inst_dmem_n17340), .ZN(MEM_stage_inst_dmem_n17341) );
NAND2_X1 MEM_stage_inst_dmem_U15468 ( .A1(MEM_stage_inst_dmem_ram_2447), .A2(MEM_stage_inst_dmem_n17340), .ZN(MEM_stage_inst_dmem_n17311) );
NAND2_X1 MEM_stage_inst_dmem_U15467 ( .A1(MEM_stage_inst_dmem_n21179), .A2(MEM_stage_inst_dmem_n17582), .ZN(MEM_stage_inst_dmem_n17340) );
NAND2_X1 MEM_stage_inst_dmem_U15466 ( .A1(MEM_stage_inst_dmem_n17309), .A2(MEM_stage_inst_dmem_n17308), .ZN(MEM_stage_inst_dmem_n10699) );
NAND2_X1 MEM_stage_inst_dmem_U15465 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n17307), .ZN(MEM_stage_inst_dmem_n17308) );
NAND2_X1 MEM_stage_inst_dmem_U15464 ( .A1(MEM_stage_inst_dmem_ram_2448), .A2(MEM_stage_inst_dmem_n17306), .ZN(MEM_stage_inst_dmem_n17309) );
NAND2_X1 MEM_stage_inst_dmem_U15463 ( .A1(MEM_stage_inst_dmem_n17305), .A2(MEM_stage_inst_dmem_n17304), .ZN(MEM_stage_inst_dmem_n10700) );
NAND2_X1 MEM_stage_inst_dmem_U15462 ( .A1(EX_pipeline_reg_out_6), .A2(MEM_stage_inst_dmem_n17307), .ZN(MEM_stage_inst_dmem_n17304) );
NAND2_X1 MEM_stage_inst_dmem_U15461 ( .A1(MEM_stage_inst_dmem_ram_2449), .A2(MEM_stage_inst_dmem_n17306), .ZN(MEM_stage_inst_dmem_n17305) );
NAND2_X1 MEM_stage_inst_dmem_U15460 ( .A1(MEM_stage_inst_dmem_n17303), .A2(MEM_stage_inst_dmem_n17302), .ZN(MEM_stage_inst_dmem_n10701) );
NAND2_X1 MEM_stage_inst_dmem_U15459 ( .A1(MEM_stage_inst_dmem_n18027), .A2(MEM_stage_inst_dmem_n17307), .ZN(MEM_stage_inst_dmem_n17302) );
NAND2_X1 MEM_stage_inst_dmem_U15458 ( .A1(MEM_stage_inst_dmem_ram_2450), .A2(MEM_stage_inst_dmem_n17306), .ZN(MEM_stage_inst_dmem_n17303) );
NAND2_X1 MEM_stage_inst_dmem_U15457 ( .A1(MEM_stage_inst_dmem_n17301), .A2(MEM_stage_inst_dmem_n17300), .ZN(MEM_stage_inst_dmem_n10702) );
NAND2_X1 MEM_stage_inst_dmem_U15456 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n17307), .ZN(MEM_stage_inst_dmem_n17300) );
NAND2_X1 MEM_stage_inst_dmem_U15455 ( .A1(MEM_stage_inst_dmem_ram_2451), .A2(MEM_stage_inst_dmem_n17306), .ZN(MEM_stage_inst_dmem_n17301) );
NAND2_X1 MEM_stage_inst_dmem_U15454 ( .A1(MEM_stage_inst_dmem_n17299), .A2(MEM_stage_inst_dmem_n17298), .ZN(MEM_stage_inst_dmem_n10703) );
NAND2_X1 MEM_stage_inst_dmem_U15453 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n17307), .ZN(MEM_stage_inst_dmem_n17298) );
NAND2_X1 MEM_stage_inst_dmem_U15452 ( .A1(MEM_stage_inst_dmem_ram_2452), .A2(MEM_stage_inst_dmem_n17306), .ZN(MEM_stage_inst_dmem_n17299) );
NAND2_X1 MEM_stage_inst_dmem_U15451 ( .A1(MEM_stage_inst_dmem_n17297), .A2(MEM_stage_inst_dmem_n17296), .ZN(MEM_stage_inst_dmem_n10704) );
NAND2_X1 MEM_stage_inst_dmem_U15450 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n17307), .ZN(MEM_stage_inst_dmem_n17296) );
NAND2_X1 MEM_stage_inst_dmem_U15449 ( .A1(MEM_stage_inst_dmem_ram_2453), .A2(MEM_stage_inst_dmem_n17306), .ZN(MEM_stage_inst_dmem_n17297) );
NAND2_X1 MEM_stage_inst_dmem_U15448 ( .A1(MEM_stage_inst_dmem_n17295), .A2(MEM_stage_inst_dmem_n17294), .ZN(MEM_stage_inst_dmem_n10705) );
NAND2_X1 MEM_stage_inst_dmem_U15447 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n17307), .ZN(MEM_stage_inst_dmem_n17294) );
NAND2_X1 MEM_stage_inst_dmem_U15446 ( .A1(MEM_stage_inst_dmem_ram_2454), .A2(MEM_stage_inst_dmem_n17306), .ZN(MEM_stage_inst_dmem_n17295) );
NAND2_X1 MEM_stage_inst_dmem_U15445 ( .A1(MEM_stage_inst_dmem_n17293), .A2(MEM_stage_inst_dmem_n17292), .ZN(MEM_stage_inst_dmem_n10706) );
NAND2_X1 MEM_stage_inst_dmem_U15444 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n17307), .ZN(MEM_stage_inst_dmem_n17292) );
NAND2_X1 MEM_stage_inst_dmem_U15443 ( .A1(MEM_stage_inst_dmem_ram_2455), .A2(MEM_stage_inst_dmem_n17306), .ZN(MEM_stage_inst_dmem_n17293) );
NAND2_X1 MEM_stage_inst_dmem_U15442 ( .A1(MEM_stage_inst_dmem_n17291), .A2(MEM_stage_inst_dmem_n17290), .ZN(MEM_stage_inst_dmem_n10707) );
NAND2_X1 MEM_stage_inst_dmem_U15441 ( .A1(MEM_stage_inst_dmem_n18013), .A2(MEM_stage_inst_dmem_n17307), .ZN(MEM_stage_inst_dmem_n17290) );
NAND2_X1 MEM_stage_inst_dmem_U15440 ( .A1(MEM_stage_inst_dmem_ram_2456), .A2(MEM_stage_inst_dmem_n17306), .ZN(MEM_stage_inst_dmem_n17291) );
NAND2_X1 MEM_stage_inst_dmem_U15439 ( .A1(MEM_stage_inst_dmem_n17289), .A2(MEM_stage_inst_dmem_n17288), .ZN(MEM_stage_inst_dmem_n10708) );
NAND2_X1 MEM_stage_inst_dmem_U15438 ( .A1(MEM_stage_inst_dmem_n96), .A2(MEM_stage_inst_dmem_n17307), .ZN(MEM_stage_inst_dmem_n17288) );
NAND2_X1 MEM_stage_inst_dmem_U15437 ( .A1(MEM_stage_inst_dmem_ram_2457), .A2(MEM_stage_inst_dmem_n17306), .ZN(MEM_stage_inst_dmem_n17289) );
NAND2_X1 MEM_stage_inst_dmem_U15436 ( .A1(MEM_stage_inst_dmem_n17287), .A2(MEM_stage_inst_dmem_n17286), .ZN(MEM_stage_inst_dmem_n10709) );
NAND2_X1 MEM_stage_inst_dmem_U15435 ( .A1(MEM_stage_inst_dmem_n18007), .A2(MEM_stage_inst_dmem_n17307), .ZN(MEM_stage_inst_dmem_n17286) );
NAND2_X1 MEM_stage_inst_dmem_U15434 ( .A1(MEM_stage_inst_dmem_ram_2458), .A2(MEM_stage_inst_dmem_n17306), .ZN(MEM_stage_inst_dmem_n17287) );
NAND2_X1 MEM_stage_inst_dmem_U15433 ( .A1(MEM_stage_inst_dmem_n17285), .A2(MEM_stage_inst_dmem_n17284), .ZN(MEM_stage_inst_dmem_n10710) );
NAND2_X1 MEM_stage_inst_dmem_U15432 ( .A1(MEM_stage_inst_dmem_n18004), .A2(MEM_stage_inst_dmem_n17307), .ZN(MEM_stage_inst_dmem_n17284) );
NAND2_X1 MEM_stage_inst_dmem_U15431 ( .A1(MEM_stage_inst_dmem_ram_2459), .A2(MEM_stage_inst_dmem_n17306), .ZN(MEM_stage_inst_dmem_n17285) );
NAND2_X1 MEM_stage_inst_dmem_U15430 ( .A1(MEM_stage_inst_dmem_n17283), .A2(MEM_stage_inst_dmem_n17282), .ZN(MEM_stage_inst_dmem_n10711) );
NAND2_X1 MEM_stage_inst_dmem_U15429 ( .A1(MEM_stage_inst_dmem_n18001), .A2(MEM_stage_inst_dmem_n17307), .ZN(MEM_stage_inst_dmem_n17282) );
NAND2_X1 MEM_stage_inst_dmem_U15428 ( .A1(MEM_stage_inst_dmem_ram_2460), .A2(MEM_stage_inst_dmem_n17306), .ZN(MEM_stage_inst_dmem_n17283) );
NAND2_X1 MEM_stage_inst_dmem_U15427 ( .A1(MEM_stage_inst_dmem_n17281), .A2(MEM_stage_inst_dmem_n17280), .ZN(MEM_stage_inst_dmem_n10712) );
NAND2_X1 MEM_stage_inst_dmem_U15426 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n17307), .ZN(MEM_stage_inst_dmem_n17280) );
NAND2_X1 MEM_stage_inst_dmem_U15425 ( .A1(MEM_stage_inst_dmem_ram_2461), .A2(MEM_stage_inst_dmem_n17306), .ZN(MEM_stage_inst_dmem_n17281) );
NAND2_X1 MEM_stage_inst_dmem_U15424 ( .A1(MEM_stage_inst_dmem_n17279), .A2(MEM_stage_inst_dmem_n17278), .ZN(MEM_stage_inst_dmem_n10713) );
NAND2_X1 MEM_stage_inst_dmem_U15423 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n17307), .ZN(MEM_stage_inst_dmem_n17278) );
NAND2_X1 MEM_stage_inst_dmem_U15422 ( .A1(MEM_stage_inst_dmem_ram_2462), .A2(MEM_stage_inst_dmem_n17306), .ZN(MEM_stage_inst_dmem_n17279) );
NAND2_X1 MEM_stage_inst_dmem_U15421 ( .A1(MEM_stage_inst_dmem_n17277), .A2(MEM_stage_inst_dmem_n17276), .ZN(MEM_stage_inst_dmem_n10714) );
NAND2_X1 MEM_stage_inst_dmem_U15420 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n17307), .ZN(MEM_stage_inst_dmem_n17276) );
INV_X1 MEM_stage_inst_dmem_U15419 ( .A(MEM_stage_inst_dmem_n17306), .ZN(MEM_stage_inst_dmem_n17307) );
NAND2_X1 MEM_stage_inst_dmem_U15418 ( .A1(MEM_stage_inst_dmem_ram_2463), .A2(MEM_stage_inst_dmem_n17306), .ZN(MEM_stage_inst_dmem_n17277) );
NAND2_X1 MEM_stage_inst_dmem_U15417 ( .A1(MEM_stage_inst_dmem_n21144), .A2(MEM_stage_inst_dmem_n17582), .ZN(MEM_stage_inst_dmem_n17306) );
NAND2_X1 MEM_stage_inst_dmem_U15416 ( .A1(MEM_stage_inst_dmem_n17275), .A2(MEM_stage_inst_dmem_n17274), .ZN(MEM_stage_inst_dmem_n10715) );
NAND2_X1 MEM_stage_inst_dmem_U15415 ( .A1(EX_pipeline_reg_out_5), .A2(MEM_stage_inst_dmem_n17273), .ZN(MEM_stage_inst_dmem_n17274) );
NAND2_X1 MEM_stage_inst_dmem_U15414 ( .A1(MEM_stage_inst_dmem_ram_2464), .A2(MEM_stage_inst_dmem_n17272), .ZN(MEM_stage_inst_dmem_n17275) );
NAND2_X1 MEM_stage_inst_dmem_U15413 ( .A1(MEM_stage_inst_dmem_n17271), .A2(MEM_stage_inst_dmem_n17270), .ZN(MEM_stage_inst_dmem_n10716) );
NAND2_X1 MEM_stage_inst_dmem_U15412 ( .A1(EX_pipeline_reg_out_6), .A2(MEM_stage_inst_dmem_n17273), .ZN(MEM_stage_inst_dmem_n17270) );
NAND2_X1 MEM_stage_inst_dmem_U15411 ( .A1(MEM_stage_inst_dmem_ram_2465), .A2(MEM_stage_inst_dmem_n17272), .ZN(MEM_stage_inst_dmem_n17271) );
NAND2_X1 MEM_stage_inst_dmem_U15410 ( .A1(MEM_stage_inst_dmem_n17269), .A2(MEM_stage_inst_dmem_n17268), .ZN(MEM_stage_inst_dmem_n10717) );
NAND2_X1 MEM_stage_inst_dmem_U15409 ( .A1(EX_pipeline_reg_out_7), .A2(MEM_stage_inst_dmem_n17273), .ZN(MEM_stage_inst_dmem_n17268) );
NAND2_X1 MEM_stage_inst_dmem_U15408 ( .A1(MEM_stage_inst_dmem_ram_2466), .A2(MEM_stage_inst_dmem_n17272), .ZN(MEM_stage_inst_dmem_n17269) );
NAND2_X1 MEM_stage_inst_dmem_U15407 ( .A1(MEM_stage_inst_dmem_n17267), .A2(MEM_stage_inst_dmem_n17266), .ZN(MEM_stage_inst_dmem_n10718) );
NAND2_X1 MEM_stage_inst_dmem_U15406 ( .A1(EX_pipeline_reg_out_8), .A2(MEM_stage_inst_dmem_n17273), .ZN(MEM_stage_inst_dmem_n17266) );
NAND2_X1 MEM_stage_inst_dmem_U15405 ( .A1(MEM_stage_inst_dmem_ram_2467), .A2(MEM_stage_inst_dmem_n17272), .ZN(MEM_stage_inst_dmem_n17267) );
NAND2_X1 MEM_stage_inst_dmem_U15404 ( .A1(MEM_stage_inst_dmem_n17265), .A2(MEM_stage_inst_dmem_n17264), .ZN(MEM_stage_inst_dmem_n10719) );
NAND2_X1 MEM_stage_inst_dmem_U15403 ( .A1(EX_pipeline_reg_out_9), .A2(MEM_stage_inst_dmem_n17273), .ZN(MEM_stage_inst_dmem_n17264) );
NAND2_X1 MEM_stage_inst_dmem_U15402 ( .A1(MEM_stage_inst_dmem_ram_2468), .A2(MEM_stage_inst_dmem_n17272), .ZN(MEM_stage_inst_dmem_n17265) );
NAND2_X1 MEM_stage_inst_dmem_U15401 ( .A1(MEM_stage_inst_dmem_n17263), .A2(MEM_stage_inst_dmem_n17262), .ZN(MEM_stage_inst_dmem_n10720) );
NAND2_X1 MEM_stage_inst_dmem_U15400 ( .A1(EX_pipeline_reg_out_10), .A2(MEM_stage_inst_dmem_n17273), .ZN(MEM_stage_inst_dmem_n17262) );
NAND2_X1 MEM_stage_inst_dmem_U15399 ( .A1(MEM_stage_inst_dmem_ram_2469), .A2(MEM_stage_inst_dmem_n17272), .ZN(MEM_stage_inst_dmem_n17263) );
NAND2_X1 MEM_stage_inst_dmem_U15398 ( .A1(MEM_stage_inst_dmem_n17261), .A2(MEM_stage_inst_dmem_n17260), .ZN(MEM_stage_inst_dmem_n10721) );
NAND2_X1 MEM_stage_inst_dmem_U15397 ( .A1(EX_pipeline_reg_out_11), .A2(MEM_stage_inst_dmem_n17273), .ZN(MEM_stage_inst_dmem_n17260) );
NAND2_X1 MEM_stage_inst_dmem_U15396 ( .A1(MEM_stage_inst_dmem_ram_2470), .A2(MEM_stage_inst_dmem_n17272), .ZN(MEM_stage_inst_dmem_n17261) );
NAND2_X1 MEM_stage_inst_dmem_U15395 ( .A1(MEM_stage_inst_dmem_n17259), .A2(MEM_stage_inst_dmem_n17258), .ZN(MEM_stage_inst_dmem_n10722) );
NAND2_X1 MEM_stage_inst_dmem_U15394 ( .A1(EX_pipeline_reg_out_12), .A2(MEM_stage_inst_dmem_n17273), .ZN(MEM_stage_inst_dmem_n17258) );
NAND2_X1 MEM_stage_inst_dmem_U15393 ( .A1(MEM_stage_inst_dmem_ram_2471), .A2(MEM_stage_inst_dmem_n17272), .ZN(MEM_stage_inst_dmem_n17259) );
NAND2_X1 MEM_stage_inst_dmem_U15392 ( .A1(MEM_stage_inst_dmem_n17257), .A2(MEM_stage_inst_dmem_n17256), .ZN(MEM_stage_inst_dmem_n10723) );
NAND2_X1 MEM_stage_inst_dmem_U15391 ( .A1(EX_pipeline_reg_out_13), .A2(MEM_stage_inst_dmem_n17273), .ZN(MEM_stage_inst_dmem_n17256) );
NAND2_X1 MEM_stage_inst_dmem_U15390 ( .A1(MEM_stage_inst_dmem_ram_2472), .A2(MEM_stage_inst_dmem_n17272), .ZN(MEM_stage_inst_dmem_n17257) );
NAND2_X1 MEM_stage_inst_dmem_U15389 ( .A1(MEM_stage_inst_dmem_n17255), .A2(MEM_stage_inst_dmem_n17254), .ZN(MEM_stage_inst_dmem_n10724) );
NAND2_X1 MEM_stage_inst_dmem_U15388 ( .A1(EX_pipeline_reg_out_14), .A2(MEM_stage_inst_dmem_n17273), .ZN(MEM_stage_inst_dmem_n17254) );
NAND2_X1 MEM_stage_inst_dmem_U15387 ( .A1(MEM_stage_inst_dmem_ram_2473), .A2(MEM_stage_inst_dmem_n17272), .ZN(MEM_stage_inst_dmem_n17255) );
NAND2_X1 MEM_stage_inst_dmem_U15386 ( .A1(MEM_stage_inst_dmem_n17253), .A2(MEM_stage_inst_dmem_n17252), .ZN(MEM_stage_inst_dmem_n10725) );
NAND2_X1 MEM_stage_inst_dmem_U15385 ( .A1(EX_pipeline_reg_out_15), .A2(MEM_stage_inst_dmem_n17273), .ZN(MEM_stage_inst_dmem_n17252) );
NAND2_X1 MEM_stage_inst_dmem_U15384 ( .A1(MEM_stage_inst_dmem_ram_2474), .A2(MEM_stage_inst_dmem_n17272), .ZN(MEM_stage_inst_dmem_n17253) );
NAND2_X1 MEM_stage_inst_dmem_U15383 ( .A1(MEM_stage_inst_dmem_n17251), .A2(MEM_stage_inst_dmem_n17250), .ZN(MEM_stage_inst_dmem_n10726) );
NAND2_X1 MEM_stage_inst_dmem_U15382 ( .A1(EX_pipeline_reg_out_16), .A2(MEM_stage_inst_dmem_n17273), .ZN(MEM_stage_inst_dmem_n17250) );
NAND2_X1 MEM_stage_inst_dmem_U15381 ( .A1(MEM_stage_inst_dmem_ram_2475), .A2(MEM_stage_inst_dmem_n17272), .ZN(MEM_stage_inst_dmem_n17251) );
NAND2_X1 MEM_stage_inst_dmem_U15380 ( .A1(MEM_stage_inst_dmem_n17249), .A2(MEM_stage_inst_dmem_n17248), .ZN(MEM_stage_inst_dmem_n10727) );
NAND2_X1 MEM_stage_inst_dmem_U15379 ( .A1(EX_pipeline_reg_out_17), .A2(MEM_stage_inst_dmem_n17273), .ZN(MEM_stage_inst_dmem_n17248) );
NAND2_X1 MEM_stage_inst_dmem_U15378 ( .A1(MEM_stage_inst_dmem_ram_2476), .A2(MEM_stage_inst_dmem_n17272), .ZN(MEM_stage_inst_dmem_n17249) );
NAND2_X1 MEM_stage_inst_dmem_U15377 ( .A1(MEM_stage_inst_dmem_n17247), .A2(MEM_stage_inst_dmem_n17246), .ZN(MEM_stage_inst_dmem_n10728) );
NAND2_X1 MEM_stage_inst_dmem_U15376 ( .A1(EX_pipeline_reg_out_18), .A2(MEM_stage_inst_dmem_n17273), .ZN(MEM_stage_inst_dmem_n17246) );
NAND2_X1 MEM_stage_inst_dmem_U15375 ( .A1(MEM_stage_inst_dmem_ram_2477), .A2(MEM_stage_inst_dmem_n17272), .ZN(MEM_stage_inst_dmem_n17247) );
NAND2_X1 MEM_stage_inst_dmem_U15374 ( .A1(MEM_stage_inst_dmem_n17245), .A2(MEM_stage_inst_dmem_n17244), .ZN(MEM_stage_inst_dmem_n10729) );
NAND2_X1 MEM_stage_inst_dmem_U15373 ( .A1(EX_pipeline_reg_out_19), .A2(MEM_stage_inst_dmem_n17273), .ZN(MEM_stage_inst_dmem_n17244) );
NAND2_X1 MEM_stage_inst_dmem_U15372 ( .A1(MEM_stage_inst_dmem_ram_2478), .A2(MEM_stage_inst_dmem_n17272), .ZN(MEM_stage_inst_dmem_n17245) );
NAND2_X1 MEM_stage_inst_dmem_U15371 ( .A1(MEM_stage_inst_dmem_n17243), .A2(MEM_stage_inst_dmem_n17242), .ZN(MEM_stage_inst_dmem_n10730) );
NAND2_X1 MEM_stage_inst_dmem_U15370 ( .A1(EX_pipeline_reg_out_20), .A2(MEM_stage_inst_dmem_n17273), .ZN(MEM_stage_inst_dmem_n17242) );
INV_X1 MEM_stage_inst_dmem_U15369 ( .A(MEM_stage_inst_dmem_n17272), .ZN(MEM_stage_inst_dmem_n17273) );
NAND2_X1 MEM_stage_inst_dmem_U15368 ( .A1(MEM_stage_inst_dmem_ram_2479), .A2(MEM_stage_inst_dmem_n17272), .ZN(MEM_stage_inst_dmem_n17243) );
NAND2_X1 MEM_stage_inst_dmem_U15367 ( .A1(MEM_stage_inst_dmem_n21109), .A2(MEM_stage_inst_dmem_n17582), .ZN(MEM_stage_inst_dmem_n17272) );
NAND2_X1 MEM_stage_inst_dmem_U15366 ( .A1(MEM_stage_inst_dmem_n17241), .A2(MEM_stage_inst_dmem_n17240), .ZN(MEM_stage_inst_dmem_n10731) );
NAND2_X1 MEM_stage_inst_dmem_U15365 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n17239), .ZN(MEM_stage_inst_dmem_n17240) );
NAND2_X1 MEM_stage_inst_dmem_U15364 ( .A1(MEM_stage_inst_dmem_ram_2480), .A2(MEM_stage_inst_dmem_n17238), .ZN(MEM_stage_inst_dmem_n17241) );
NAND2_X1 MEM_stage_inst_dmem_U15363 ( .A1(MEM_stage_inst_dmem_n17237), .A2(MEM_stage_inst_dmem_n17236), .ZN(MEM_stage_inst_dmem_n10732) );
NAND2_X1 MEM_stage_inst_dmem_U15362 ( .A1(MEM_stage_inst_dmem_n20547), .A2(MEM_stage_inst_dmem_n17239), .ZN(MEM_stage_inst_dmem_n17236) );
NAND2_X1 MEM_stage_inst_dmem_U15361 ( .A1(MEM_stage_inst_dmem_ram_2481), .A2(MEM_stage_inst_dmem_n17238), .ZN(MEM_stage_inst_dmem_n17237) );
NAND2_X1 MEM_stage_inst_dmem_U15360 ( .A1(MEM_stage_inst_dmem_n17235), .A2(MEM_stage_inst_dmem_n17234), .ZN(MEM_stage_inst_dmem_n10733) );
NAND2_X1 MEM_stage_inst_dmem_U15359 ( .A1(MEM_stage_inst_dmem_n18027), .A2(MEM_stage_inst_dmem_n17239), .ZN(MEM_stage_inst_dmem_n17234) );
NAND2_X1 MEM_stage_inst_dmem_U15358 ( .A1(MEM_stage_inst_dmem_ram_2482), .A2(MEM_stage_inst_dmem_n17238), .ZN(MEM_stage_inst_dmem_n17235) );
NAND2_X1 MEM_stage_inst_dmem_U15357 ( .A1(MEM_stage_inst_dmem_n17233), .A2(MEM_stage_inst_dmem_n17232), .ZN(MEM_stage_inst_dmem_n10734) );
NAND2_X1 MEM_stage_inst_dmem_U15356 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n17239), .ZN(MEM_stage_inst_dmem_n17232) );
NAND2_X1 MEM_stage_inst_dmem_U15355 ( .A1(MEM_stage_inst_dmem_ram_2483), .A2(MEM_stage_inst_dmem_n17238), .ZN(MEM_stage_inst_dmem_n17233) );
NAND2_X1 MEM_stage_inst_dmem_U15354 ( .A1(MEM_stage_inst_dmem_n17231), .A2(MEM_stage_inst_dmem_n17230), .ZN(MEM_stage_inst_dmem_n10735) );
NAND2_X1 MEM_stage_inst_dmem_U15353 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n17239), .ZN(MEM_stage_inst_dmem_n17230) );
NAND2_X1 MEM_stage_inst_dmem_U15352 ( .A1(MEM_stage_inst_dmem_ram_2484), .A2(MEM_stage_inst_dmem_n17238), .ZN(MEM_stage_inst_dmem_n17231) );
NAND2_X1 MEM_stage_inst_dmem_U15351 ( .A1(MEM_stage_inst_dmem_n17229), .A2(MEM_stage_inst_dmem_n17228), .ZN(MEM_stage_inst_dmem_n10736) );
NAND2_X1 MEM_stage_inst_dmem_U15350 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n17239), .ZN(MEM_stage_inst_dmem_n17228) );
NAND2_X1 MEM_stage_inst_dmem_U15349 ( .A1(MEM_stage_inst_dmem_ram_2485), .A2(MEM_stage_inst_dmem_n17238), .ZN(MEM_stage_inst_dmem_n17229) );
NAND2_X1 MEM_stage_inst_dmem_U15348 ( .A1(MEM_stage_inst_dmem_n17227), .A2(MEM_stage_inst_dmem_n17226), .ZN(MEM_stage_inst_dmem_n10737) );
NAND2_X1 MEM_stage_inst_dmem_U15347 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n17239), .ZN(MEM_stage_inst_dmem_n17226) );
NAND2_X1 MEM_stage_inst_dmem_U15346 ( .A1(MEM_stage_inst_dmem_ram_2486), .A2(MEM_stage_inst_dmem_n17238), .ZN(MEM_stage_inst_dmem_n17227) );
NAND2_X1 MEM_stage_inst_dmem_U15345 ( .A1(MEM_stage_inst_dmem_n17225), .A2(MEM_stage_inst_dmem_n17224), .ZN(MEM_stage_inst_dmem_n10738) );
NAND2_X1 MEM_stage_inst_dmem_U15344 ( .A1(MEM_stage_inst_dmem_n112), .A2(MEM_stage_inst_dmem_n17239), .ZN(MEM_stage_inst_dmem_n17224) );
NAND2_X1 MEM_stage_inst_dmem_U15343 ( .A1(MEM_stage_inst_dmem_ram_2487), .A2(MEM_stage_inst_dmem_n17238), .ZN(MEM_stage_inst_dmem_n17225) );
NAND2_X1 MEM_stage_inst_dmem_U15342 ( .A1(MEM_stage_inst_dmem_n17223), .A2(MEM_stage_inst_dmem_n17222), .ZN(MEM_stage_inst_dmem_n10739) );
NAND2_X1 MEM_stage_inst_dmem_U15341 ( .A1(MEM_stage_inst_dmem_n18013), .A2(MEM_stage_inst_dmem_n17239), .ZN(MEM_stage_inst_dmem_n17222) );
NAND2_X1 MEM_stage_inst_dmem_U15340 ( .A1(MEM_stage_inst_dmem_ram_2488), .A2(MEM_stage_inst_dmem_n17238), .ZN(MEM_stage_inst_dmem_n17223) );
NAND2_X1 MEM_stage_inst_dmem_U15339 ( .A1(MEM_stage_inst_dmem_n17221), .A2(MEM_stage_inst_dmem_n17220), .ZN(MEM_stage_inst_dmem_n10740) );
NAND2_X1 MEM_stage_inst_dmem_U15338 ( .A1(MEM_stage_inst_dmem_n96), .A2(MEM_stage_inst_dmem_n17239), .ZN(MEM_stage_inst_dmem_n17220) );
NAND2_X1 MEM_stage_inst_dmem_U15337 ( .A1(MEM_stage_inst_dmem_ram_2489), .A2(MEM_stage_inst_dmem_n17238), .ZN(MEM_stage_inst_dmem_n17221) );
NAND2_X1 MEM_stage_inst_dmem_U15336 ( .A1(MEM_stage_inst_dmem_n17219), .A2(MEM_stage_inst_dmem_n17218), .ZN(MEM_stage_inst_dmem_n10741) );
NAND2_X1 MEM_stage_inst_dmem_U15335 ( .A1(MEM_stage_inst_dmem_n18007), .A2(MEM_stage_inst_dmem_n17239), .ZN(MEM_stage_inst_dmem_n17218) );
NAND2_X1 MEM_stage_inst_dmem_U15334 ( .A1(MEM_stage_inst_dmem_ram_2490), .A2(MEM_stage_inst_dmem_n17238), .ZN(MEM_stage_inst_dmem_n17219) );
NAND2_X1 MEM_stage_inst_dmem_U15333 ( .A1(MEM_stage_inst_dmem_n17217), .A2(MEM_stage_inst_dmem_n17216), .ZN(MEM_stage_inst_dmem_n10742) );
NAND2_X1 MEM_stage_inst_dmem_U15332 ( .A1(MEM_stage_inst_dmem_n18004), .A2(MEM_stage_inst_dmem_n17239), .ZN(MEM_stage_inst_dmem_n17216) );
NAND2_X1 MEM_stage_inst_dmem_U15331 ( .A1(MEM_stage_inst_dmem_ram_2491), .A2(MEM_stage_inst_dmem_n17238), .ZN(MEM_stage_inst_dmem_n17217) );
NAND2_X1 MEM_stage_inst_dmem_U15330 ( .A1(MEM_stage_inst_dmem_n17215), .A2(MEM_stage_inst_dmem_n17214), .ZN(MEM_stage_inst_dmem_n10743) );
NAND2_X1 MEM_stage_inst_dmem_U15329 ( .A1(MEM_stage_inst_dmem_n18001), .A2(MEM_stage_inst_dmem_n17239), .ZN(MEM_stage_inst_dmem_n17214) );
NAND2_X1 MEM_stage_inst_dmem_U15328 ( .A1(MEM_stage_inst_dmem_ram_2492), .A2(MEM_stage_inst_dmem_n17238), .ZN(MEM_stage_inst_dmem_n17215) );
NAND2_X1 MEM_stage_inst_dmem_U15327 ( .A1(MEM_stage_inst_dmem_n17213), .A2(MEM_stage_inst_dmem_n17212), .ZN(MEM_stage_inst_dmem_n10744) );
NAND2_X1 MEM_stage_inst_dmem_U15326 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n17239), .ZN(MEM_stage_inst_dmem_n17212) );
NAND2_X1 MEM_stage_inst_dmem_U15325 ( .A1(MEM_stage_inst_dmem_ram_2493), .A2(MEM_stage_inst_dmem_n17238), .ZN(MEM_stage_inst_dmem_n17213) );
NAND2_X1 MEM_stage_inst_dmem_U15324 ( .A1(MEM_stage_inst_dmem_n17211), .A2(MEM_stage_inst_dmem_n17210), .ZN(MEM_stage_inst_dmem_n10745) );
NAND2_X1 MEM_stage_inst_dmem_U15323 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n17239), .ZN(MEM_stage_inst_dmem_n17210) );
NAND2_X1 MEM_stage_inst_dmem_U15322 ( .A1(MEM_stage_inst_dmem_ram_2494), .A2(MEM_stage_inst_dmem_n17238), .ZN(MEM_stage_inst_dmem_n17211) );
NAND2_X1 MEM_stage_inst_dmem_U15321 ( .A1(MEM_stage_inst_dmem_n17209), .A2(MEM_stage_inst_dmem_n17208), .ZN(MEM_stage_inst_dmem_n10746) );
NAND2_X1 MEM_stage_inst_dmem_U15320 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n17239), .ZN(MEM_stage_inst_dmem_n17208) );
INV_X1 MEM_stage_inst_dmem_U15319 ( .A(MEM_stage_inst_dmem_n17238), .ZN(MEM_stage_inst_dmem_n17239) );
NAND2_X1 MEM_stage_inst_dmem_U15318 ( .A1(MEM_stage_inst_dmem_ram_2495), .A2(MEM_stage_inst_dmem_n17238), .ZN(MEM_stage_inst_dmem_n17209) );
NAND2_X1 MEM_stage_inst_dmem_U15317 ( .A1(MEM_stage_inst_dmem_n21074), .A2(MEM_stage_inst_dmem_n17582), .ZN(MEM_stage_inst_dmem_n17238) );
NAND2_X1 MEM_stage_inst_dmem_U15316 ( .A1(MEM_stage_inst_dmem_n17207), .A2(MEM_stage_inst_dmem_n17206), .ZN(MEM_stage_inst_dmem_n10747) );
NAND2_X1 MEM_stage_inst_dmem_U15315 ( .A1(EX_pipeline_reg_out_5), .A2(MEM_stage_inst_dmem_n17205), .ZN(MEM_stage_inst_dmem_n17206) );
NAND2_X1 MEM_stage_inst_dmem_U15314 ( .A1(MEM_stage_inst_dmem_ram_2496), .A2(MEM_stage_inst_dmem_n17204), .ZN(MEM_stage_inst_dmem_n17207) );
NAND2_X1 MEM_stage_inst_dmem_U15313 ( .A1(MEM_stage_inst_dmem_n17203), .A2(MEM_stage_inst_dmem_n17202), .ZN(MEM_stage_inst_dmem_n10748) );
NAND2_X1 MEM_stage_inst_dmem_U15312 ( .A1(EX_pipeline_reg_out_6), .A2(MEM_stage_inst_dmem_n17205), .ZN(MEM_stage_inst_dmem_n17202) );
NAND2_X1 MEM_stage_inst_dmem_U15311 ( .A1(MEM_stage_inst_dmem_ram_2497), .A2(MEM_stage_inst_dmem_n17204), .ZN(MEM_stage_inst_dmem_n17203) );
NAND2_X1 MEM_stage_inst_dmem_U15310 ( .A1(MEM_stage_inst_dmem_n17201), .A2(MEM_stage_inst_dmem_n17200), .ZN(MEM_stage_inst_dmem_n10749) );
NAND2_X1 MEM_stage_inst_dmem_U15309 ( .A1(EX_pipeline_reg_out_7), .A2(MEM_stage_inst_dmem_n17205), .ZN(MEM_stage_inst_dmem_n17200) );
NAND2_X1 MEM_stage_inst_dmem_U15308 ( .A1(MEM_stage_inst_dmem_ram_2498), .A2(MEM_stage_inst_dmem_n17204), .ZN(MEM_stage_inst_dmem_n17201) );
NAND2_X1 MEM_stage_inst_dmem_U15307 ( .A1(MEM_stage_inst_dmem_n17199), .A2(MEM_stage_inst_dmem_n17198), .ZN(MEM_stage_inst_dmem_n10750) );
NAND2_X1 MEM_stage_inst_dmem_U15306 ( .A1(EX_pipeline_reg_out_8), .A2(MEM_stage_inst_dmem_n17205), .ZN(MEM_stage_inst_dmem_n17198) );
NAND2_X1 MEM_stage_inst_dmem_U15305 ( .A1(MEM_stage_inst_dmem_ram_2499), .A2(MEM_stage_inst_dmem_n17204), .ZN(MEM_stage_inst_dmem_n17199) );
NAND2_X1 MEM_stage_inst_dmem_U15304 ( .A1(MEM_stage_inst_dmem_n17197), .A2(MEM_stage_inst_dmem_n17196), .ZN(MEM_stage_inst_dmem_n10751) );
NAND2_X1 MEM_stage_inst_dmem_U15303 ( .A1(EX_pipeline_reg_out_9), .A2(MEM_stage_inst_dmem_n17205), .ZN(MEM_stage_inst_dmem_n17196) );
NAND2_X1 MEM_stage_inst_dmem_U15302 ( .A1(MEM_stage_inst_dmem_ram_2500), .A2(MEM_stage_inst_dmem_n17204), .ZN(MEM_stage_inst_dmem_n17197) );
NAND2_X1 MEM_stage_inst_dmem_U15301 ( .A1(MEM_stage_inst_dmem_n17195), .A2(MEM_stage_inst_dmem_n17194), .ZN(MEM_stage_inst_dmem_n10752) );
NAND2_X1 MEM_stage_inst_dmem_U15300 ( .A1(EX_pipeline_reg_out_10), .A2(MEM_stage_inst_dmem_n17205), .ZN(MEM_stage_inst_dmem_n17194) );
NAND2_X1 MEM_stage_inst_dmem_U15299 ( .A1(MEM_stage_inst_dmem_ram_2501), .A2(MEM_stage_inst_dmem_n17204), .ZN(MEM_stage_inst_dmem_n17195) );
NAND2_X1 MEM_stage_inst_dmem_U15298 ( .A1(MEM_stage_inst_dmem_n17193), .A2(MEM_stage_inst_dmem_n17192), .ZN(MEM_stage_inst_dmem_n10753) );
NAND2_X1 MEM_stage_inst_dmem_U15297 ( .A1(EX_pipeline_reg_out_11), .A2(MEM_stage_inst_dmem_n17205), .ZN(MEM_stage_inst_dmem_n17192) );
NAND2_X1 MEM_stage_inst_dmem_U15296 ( .A1(MEM_stage_inst_dmem_ram_2502), .A2(MEM_stage_inst_dmem_n17204), .ZN(MEM_stage_inst_dmem_n17193) );
NAND2_X1 MEM_stage_inst_dmem_U15295 ( .A1(MEM_stage_inst_dmem_n17191), .A2(MEM_stage_inst_dmem_n17190), .ZN(MEM_stage_inst_dmem_n10754) );
NAND2_X1 MEM_stage_inst_dmem_U15294 ( .A1(EX_pipeline_reg_out_12), .A2(MEM_stage_inst_dmem_n17205), .ZN(MEM_stage_inst_dmem_n17190) );
NAND2_X1 MEM_stage_inst_dmem_U15293 ( .A1(MEM_stage_inst_dmem_ram_2503), .A2(MEM_stage_inst_dmem_n17204), .ZN(MEM_stage_inst_dmem_n17191) );
NAND2_X1 MEM_stage_inst_dmem_U15292 ( .A1(MEM_stage_inst_dmem_n17189), .A2(MEM_stage_inst_dmem_n17188), .ZN(MEM_stage_inst_dmem_n10755) );
NAND2_X1 MEM_stage_inst_dmem_U15291 ( .A1(EX_pipeline_reg_out_13), .A2(MEM_stage_inst_dmem_n17205), .ZN(MEM_stage_inst_dmem_n17188) );
NAND2_X1 MEM_stage_inst_dmem_U15290 ( .A1(MEM_stage_inst_dmem_ram_2504), .A2(MEM_stage_inst_dmem_n17204), .ZN(MEM_stage_inst_dmem_n17189) );
NAND2_X1 MEM_stage_inst_dmem_U15289 ( .A1(MEM_stage_inst_dmem_n17187), .A2(MEM_stage_inst_dmem_n17186), .ZN(MEM_stage_inst_dmem_n10756) );
NAND2_X1 MEM_stage_inst_dmem_U15288 ( .A1(EX_pipeline_reg_out_14), .A2(MEM_stage_inst_dmem_n17205), .ZN(MEM_stage_inst_dmem_n17186) );
NAND2_X1 MEM_stage_inst_dmem_U15287 ( .A1(MEM_stage_inst_dmem_ram_2505), .A2(MEM_stage_inst_dmem_n17204), .ZN(MEM_stage_inst_dmem_n17187) );
NAND2_X1 MEM_stage_inst_dmem_U15286 ( .A1(MEM_stage_inst_dmem_n17185), .A2(MEM_stage_inst_dmem_n17184), .ZN(MEM_stage_inst_dmem_n10757) );
NAND2_X1 MEM_stage_inst_dmem_U15285 ( .A1(EX_pipeline_reg_out_15), .A2(MEM_stage_inst_dmem_n17205), .ZN(MEM_stage_inst_dmem_n17184) );
NAND2_X1 MEM_stage_inst_dmem_U15284 ( .A1(MEM_stage_inst_dmem_ram_2506), .A2(MEM_stage_inst_dmem_n17204), .ZN(MEM_stage_inst_dmem_n17185) );
NAND2_X1 MEM_stage_inst_dmem_U15283 ( .A1(MEM_stage_inst_dmem_n17183), .A2(MEM_stage_inst_dmem_n17182), .ZN(MEM_stage_inst_dmem_n10758) );
NAND2_X1 MEM_stage_inst_dmem_U15282 ( .A1(EX_pipeline_reg_out_16), .A2(MEM_stage_inst_dmem_n17205), .ZN(MEM_stage_inst_dmem_n17182) );
NAND2_X1 MEM_stage_inst_dmem_U15281 ( .A1(MEM_stage_inst_dmem_ram_2507), .A2(MEM_stage_inst_dmem_n17204), .ZN(MEM_stage_inst_dmem_n17183) );
NAND2_X1 MEM_stage_inst_dmem_U15280 ( .A1(MEM_stage_inst_dmem_n17181), .A2(MEM_stage_inst_dmem_n17180), .ZN(MEM_stage_inst_dmem_n10759) );
NAND2_X1 MEM_stage_inst_dmem_U15279 ( .A1(EX_pipeline_reg_out_17), .A2(MEM_stage_inst_dmem_n17205), .ZN(MEM_stage_inst_dmem_n17180) );
NAND2_X1 MEM_stage_inst_dmem_U15278 ( .A1(MEM_stage_inst_dmem_ram_2508), .A2(MEM_stage_inst_dmem_n17204), .ZN(MEM_stage_inst_dmem_n17181) );
NAND2_X1 MEM_stage_inst_dmem_U15277 ( .A1(MEM_stage_inst_dmem_n17179), .A2(MEM_stage_inst_dmem_n17178), .ZN(MEM_stage_inst_dmem_n10760) );
NAND2_X1 MEM_stage_inst_dmem_U15276 ( .A1(EX_pipeline_reg_out_18), .A2(MEM_stage_inst_dmem_n17205), .ZN(MEM_stage_inst_dmem_n17178) );
NAND2_X1 MEM_stage_inst_dmem_U15275 ( .A1(MEM_stage_inst_dmem_ram_2509), .A2(MEM_stage_inst_dmem_n17204), .ZN(MEM_stage_inst_dmem_n17179) );
NAND2_X1 MEM_stage_inst_dmem_U15274 ( .A1(MEM_stage_inst_dmem_n17177), .A2(MEM_stage_inst_dmem_n17176), .ZN(MEM_stage_inst_dmem_n10761) );
NAND2_X1 MEM_stage_inst_dmem_U15273 ( .A1(EX_pipeline_reg_out_19), .A2(MEM_stage_inst_dmem_n17205), .ZN(MEM_stage_inst_dmem_n17176) );
NAND2_X1 MEM_stage_inst_dmem_U15272 ( .A1(MEM_stage_inst_dmem_ram_2510), .A2(MEM_stage_inst_dmem_n17204), .ZN(MEM_stage_inst_dmem_n17177) );
NAND2_X1 MEM_stage_inst_dmem_U15271 ( .A1(MEM_stage_inst_dmem_n17175), .A2(MEM_stage_inst_dmem_n17174), .ZN(MEM_stage_inst_dmem_n10762) );
NAND2_X1 MEM_stage_inst_dmem_U15270 ( .A1(EX_pipeline_reg_out_20), .A2(MEM_stage_inst_dmem_n17205), .ZN(MEM_stage_inst_dmem_n17174) );
INV_X1 MEM_stage_inst_dmem_U15269 ( .A(MEM_stage_inst_dmem_n17204), .ZN(MEM_stage_inst_dmem_n17205) );
NAND2_X1 MEM_stage_inst_dmem_U15268 ( .A1(MEM_stage_inst_dmem_ram_2511), .A2(MEM_stage_inst_dmem_n17204), .ZN(MEM_stage_inst_dmem_n17175) );
NAND2_X1 MEM_stage_inst_dmem_U15267 ( .A1(MEM_stage_inst_dmem_n21039), .A2(MEM_stage_inst_dmem_n17582), .ZN(MEM_stage_inst_dmem_n17204) );
NAND2_X1 MEM_stage_inst_dmem_U15266 ( .A1(MEM_stage_inst_dmem_n17173), .A2(MEM_stage_inst_dmem_n17172), .ZN(MEM_stage_inst_dmem_n10763) );
NAND2_X1 MEM_stage_inst_dmem_U15265 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n17171), .ZN(MEM_stage_inst_dmem_n17172) );
NAND2_X1 MEM_stage_inst_dmem_U15264 ( .A1(MEM_stage_inst_dmem_ram_2512), .A2(MEM_stage_inst_dmem_n17170), .ZN(MEM_stage_inst_dmem_n17173) );
NAND2_X1 MEM_stage_inst_dmem_U15263 ( .A1(MEM_stage_inst_dmem_n17169), .A2(MEM_stage_inst_dmem_n17168), .ZN(MEM_stage_inst_dmem_n10764) );
NAND2_X1 MEM_stage_inst_dmem_U15262 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n17171), .ZN(MEM_stage_inst_dmem_n17168) );
NAND2_X1 MEM_stage_inst_dmem_U15261 ( .A1(MEM_stage_inst_dmem_ram_2513), .A2(MEM_stage_inst_dmem_n17170), .ZN(MEM_stage_inst_dmem_n17169) );
NAND2_X1 MEM_stage_inst_dmem_U15260 ( .A1(MEM_stage_inst_dmem_n17167), .A2(MEM_stage_inst_dmem_n17166), .ZN(MEM_stage_inst_dmem_n10765) );
NAND2_X1 MEM_stage_inst_dmem_U15259 ( .A1(MEM_stage_inst_dmem_n18027), .A2(MEM_stage_inst_dmem_n17171), .ZN(MEM_stage_inst_dmem_n17166) );
NAND2_X1 MEM_stage_inst_dmem_U15258 ( .A1(MEM_stage_inst_dmem_ram_2514), .A2(MEM_stage_inst_dmem_n17170), .ZN(MEM_stage_inst_dmem_n17167) );
NAND2_X1 MEM_stage_inst_dmem_U15257 ( .A1(MEM_stage_inst_dmem_n17165), .A2(MEM_stage_inst_dmem_n17164), .ZN(MEM_stage_inst_dmem_n10766) );
NAND2_X1 MEM_stage_inst_dmem_U15256 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n17171), .ZN(MEM_stage_inst_dmem_n17164) );
NAND2_X1 MEM_stage_inst_dmem_U15255 ( .A1(MEM_stage_inst_dmem_ram_2515), .A2(MEM_stage_inst_dmem_n17170), .ZN(MEM_stage_inst_dmem_n17165) );
NAND2_X1 MEM_stage_inst_dmem_U15254 ( .A1(MEM_stage_inst_dmem_n17163), .A2(MEM_stage_inst_dmem_n17162), .ZN(MEM_stage_inst_dmem_n10767) );
NAND2_X1 MEM_stage_inst_dmem_U15253 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n17171), .ZN(MEM_stage_inst_dmem_n17162) );
NAND2_X1 MEM_stage_inst_dmem_U15252 ( .A1(MEM_stage_inst_dmem_ram_2516), .A2(MEM_stage_inst_dmem_n17170), .ZN(MEM_stage_inst_dmem_n17163) );
NAND2_X1 MEM_stage_inst_dmem_U15251 ( .A1(MEM_stage_inst_dmem_n17161), .A2(MEM_stage_inst_dmem_n17160), .ZN(MEM_stage_inst_dmem_n10768) );
NAND2_X1 MEM_stage_inst_dmem_U15250 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n17171), .ZN(MEM_stage_inst_dmem_n17160) );
NAND2_X1 MEM_stage_inst_dmem_U15249 ( .A1(MEM_stage_inst_dmem_ram_2517), .A2(MEM_stage_inst_dmem_n17170), .ZN(MEM_stage_inst_dmem_n17161) );
NAND2_X1 MEM_stage_inst_dmem_U15248 ( .A1(MEM_stage_inst_dmem_n17159), .A2(MEM_stage_inst_dmem_n17158), .ZN(MEM_stage_inst_dmem_n10769) );
NAND2_X1 MEM_stage_inst_dmem_U15247 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n17171), .ZN(MEM_stage_inst_dmem_n17158) );
NAND2_X1 MEM_stage_inst_dmem_U15246 ( .A1(MEM_stage_inst_dmem_ram_2518), .A2(MEM_stage_inst_dmem_n17170), .ZN(MEM_stage_inst_dmem_n17159) );
NAND2_X1 MEM_stage_inst_dmem_U15245 ( .A1(MEM_stage_inst_dmem_n17157), .A2(MEM_stage_inst_dmem_n17156), .ZN(MEM_stage_inst_dmem_n10770) );
NAND2_X1 MEM_stage_inst_dmem_U15244 ( .A1(MEM_stage_inst_dmem_n112), .A2(MEM_stage_inst_dmem_n17171), .ZN(MEM_stage_inst_dmem_n17156) );
NAND2_X1 MEM_stage_inst_dmem_U15243 ( .A1(MEM_stage_inst_dmem_ram_2519), .A2(MEM_stage_inst_dmem_n17170), .ZN(MEM_stage_inst_dmem_n17157) );
NAND2_X1 MEM_stage_inst_dmem_U15242 ( .A1(MEM_stage_inst_dmem_n17155), .A2(MEM_stage_inst_dmem_n17154), .ZN(MEM_stage_inst_dmem_n10771) );
NAND2_X1 MEM_stage_inst_dmem_U15241 ( .A1(MEM_stage_inst_dmem_n18013), .A2(MEM_stage_inst_dmem_n17171), .ZN(MEM_stage_inst_dmem_n17154) );
NAND2_X1 MEM_stage_inst_dmem_U15240 ( .A1(MEM_stage_inst_dmem_ram_2520), .A2(MEM_stage_inst_dmem_n17170), .ZN(MEM_stage_inst_dmem_n17155) );
NAND2_X1 MEM_stage_inst_dmem_U15239 ( .A1(MEM_stage_inst_dmem_n17153), .A2(MEM_stage_inst_dmem_n17152), .ZN(MEM_stage_inst_dmem_n10772) );
NAND2_X1 MEM_stage_inst_dmem_U15238 ( .A1(MEM_stage_inst_dmem_n96), .A2(MEM_stage_inst_dmem_n17171), .ZN(MEM_stage_inst_dmem_n17152) );
NAND2_X1 MEM_stage_inst_dmem_U15237 ( .A1(MEM_stage_inst_dmem_ram_2521), .A2(MEM_stage_inst_dmem_n17170), .ZN(MEM_stage_inst_dmem_n17153) );
NAND2_X1 MEM_stage_inst_dmem_U15236 ( .A1(MEM_stage_inst_dmem_n17151), .A2(MEM_stage_inst_dmem_n17150), .ZN(MEM_stage_inst_dmem_n10773) );
NAND2_X1 MEM_stage_inst_dmem_U15235 ( .A1(MEM_stage_inst_dmem_n18007), .A2(MEM_stage_inst_dmem_n17171), .ZN(MEM_stage_inst_dmem_n17150) );
NAND2_X1 MEM_stage_inst_dmem_U15234 ( .A1(MEM_stage_inst_dmem_ram_2522), .A2(MEM_stage_inst_dmem_n17170), .ZN(MEM_stage_inst_dmem_n17151) );
NAND2_X1 MEM_stage_inst_dmem_U15233 ( .A1(MEM_stage_inst_dmem_n17149), .A2(MEM_stage_inst_dmem_n17148), .ZN(MEM_stage_inst_dmem_n10774) );
NAND2_X1 MEM_stage_inst_dmem_U15232 ( .A1(MEM_stage_inst_dmem_n18004), .A2(MEM_stage_inst_dmem_n17171), .ZN(MEM_stage_inst_dmem_n17148) );
NAND2_X1 MEM_stage_inst_dmem_U15231 ( .A1(MEM_stage_inst_dmem_ram_2523), .A2(MEM_stage_inst_dmem_n17170), .ZN(MEM_stage_inst_dmem_n17149) );
NAND2_X1 MEM_stage_inst_dmem_U15230 ( .A1(MEM_stage_inst_dmem_n17147), .A2(MEM_stage_inst_dmem_n17146), .ZN(MEM_stage_inst_dmem_n10775) );
NAND2_X1 MEM_stage_inst_dmem_U15229 ( .A1(MEM_stage_inst_dmem_n18001), .A2(MEM_stage_inst_dmem_n17171), .ZN(MEM_stage_inst_dmem_n17146) );
NAND2_X1 MEM_stage_inst_dmem_U15228 ( .A1(MEM_stage_inst_dmem_ram_2524), .A2(MEM_stage_inst_dmem_n17170), .ZN(MEM_stage_inst_dmem_n17147) );
NAND2_X1 MEM_stage_inst_dmem_U15227 ( .A1(MEM_stage_inst_dmem_n17145), .A2(MEM_stage_inst_dmem_n17144), .ZN(MEM_stage_inst_dmem_n10776) );
NAND2_X1 MEM_stage_inst_dmem_U15226 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n17171), .ZN(MEM_stage_inst_dmem_n17144) );
NAND2_X1 MEM_stage_inst_dmem_U15225 ( .A1(MEM_stage_inst_dmem_ram_2525), .A2(MEM_stage_inst_dmem_n17170), .ZN(MEM_stage_inst_dmem_n17145) );
NAND2_X1 MEM_stage_inst_dmem_U15224 ( .A1(MEM_stage_inst_dmem_n17143), .A2(MEM_stage_inst_dmem_n17142), .ZN(MEM_stage_inst_dmem_n10777) );
NAND2_X1 MEM_stage_inst_dmem_U15223 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n17171), .ZN(MEM_stage_inst_dmem_n17142) );
NAND2_X1 MEM_stage_inst_dmem_U15222 ( .A1(MEM_stage_inst_dmem_ram_2526), .A2(MEM_stage_inst_dmem_n17170), .ZN(MEM_stage_inst_dmem_n17143) );
NAND2_X1 MEM_stage_inst_dmem_U15221 ( .A1(MEM_stage_inst_dmem_n17141), .A2(MEM_stage_inst_dmem_n17140), .ZN(MEM_stage_inst_dmem_n10778) );
NAND2_X1 MEM_stage_inst_dmem_U15220 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n17171), .ZN(MEM_stage_inst_dmem_n17140) );
INV_X1 MEM_stage_inst_dmem_U15219 ( .A(MEM_stage_inst_dmem_n17170), .ZN(MEM_stage_inst_dmem_n17171) );
NAND2_X1 MEM_stage_inst_dmem_U15218 ( .A1(MEM_stage_inst_dmem_ram_2527), .A2(MEM_stage_inst_dmem_n17170), .ZN(MEM_stage_inst_dmem_n17141) );
NAND2_X1 MEM_stage_inst_dmem_U15217 ( .A1(MEM_stage_inst_dmem_n21004), .A2(MEM_stage_inst_dmem_n17582), .ZN(MEM_stage_inst_dmem_n17170) );
NAND2_X1 MEM_stage_inst_dmem_U15216 ( .A1(MEM_stage_inst_dmem_n17139), .A2(MEM_stage_inst_dmem_n17138), .ZN(MEM_stage_inst_dmem_n10779) );
NAND2_X1 MEM_stage_inst_dmem_U15215 ( .A1(EX_pipeline_reg_out_5), .A2(MEM_stage_inst_dmem_n17137), .ZN(MEM_stage_inst_dmem_n17138) );
NAND2_X1 MEM_stage_inst_dmem_U15214 ( .A1(MEM_stage_inst_dmem_ram_2528), .A2(MEM_stage_inst_dmem_n17136), .ZN(MEM_stage_inst_dmem_n17139) );
NAND2_X1 MEM_stage_inst_dmem_U15213 ( .A1(MEM_stage_inst_dmem_n17135), .A2(MEM_stage_inst_dmem_n17134), .ZN(MEM_stage_inst_dmem_n10780) );
NAND2_X1 MEM_stage_inst_dmem_U15212 ( .A1(EX_pipeline_reg_out_6), .A2(MEM_stage_inst_dmem_n17137), .ZN(MEM_stage_inst_dmem_n17134) );
NAND2_X1 MEM_stage_inst_dmem_U15211 ( .A1(MEM_stage_inst_dmem_ram_2529), .A2(MEM_stage_inst_dmem_n17136), .ZN(MEM_stage_inst_dmem_n17135) );
NAND2_X1 MEM_stage_inst_dmem_U15210 ( .A1(MEM_stage_inst_dmem_n17133), .A2(MEM_stage_inst_dmem_n17132), .ZN(MEM_stage_inst_dmem_n10781) );
NAND2_X1 MEM_stage_inst_dmem_U15209 ( .A1(EX_pipeline_reg_out_7), .A2(MEM_stage_inst_dmem_n17137), .ZN(MEM_stage_inst_dmem_n17132) );
NAND2_X1 MEM_stage_inst_dmem_U15208 ( .A1(MEM_stage_inst_dmem_ram_2530), .A2(MEM_stage_inst_dmem_n17136), .ZN(MEM_stage_inst_dmem_n17133) );
NAND2_X1 MEM_stage_inst_dmem_U15207 ( .A1(MEM_stage_inst_dmem_n17131), .A2(MEM_stage_inst_dmem_n17130), .ZN(MEM_stage_inst_dmem_n10782) );
NAND2_X1 MEM_stage_inst_dmem_U15206 ( .A1(EX_pipeline_reg_out_8), .A2(MEM_stage_inst_dmem_n17137), .ZN(MEM_stage_inst_dmem_n17130) );
NAND2_X1 MEM_stage_inst_dmem_U15205 ( .A1(MEM_stage_inst_dmem_ram_2531), .A2(MEM_stage_inst_dmem_n17136), .ZN(MEM_stage_inst_dmem_n17131) );
NAND2_X1 MEM_stage_inst_dmem_U15204 ( .A1(MEM_stage_inst_dmem_n17129), .A2(MEM_stage_inst_dmem_n17128), .ZN(MEM_stage_inst_dmem_n10783) );
NAND2_X1 MEM_stage_inst_dmem_U15203 ( .A1(EX_pipeline_reg_out_9), .A2(MEM_stage_inst_dmem_n17137), .ZN(MEM_stage_inst_dmem_n17128) );
NAND2_X1 MEM_stage_inst_dmem_U15202 ( .A1(MEM_stage_inst_dmem_ram_2532), .A2(MEM_stage_inst_dmem_n17136), .ZN(MEM_stage_inst_dmem_n17129) );
NAND2_X1 MEM_stage_inst_dmem_U15201 ( .A1(MEM_stage_inst_dmem_n17127), .A2(MEM_stage_inst_dmem_n17126), .ZN(MEM_stage_inst_dmem_n10784) );
NAND2_X1 MEM_stage_inst_dmem_U15200 ( .A1(EX_pipeline_reg_out_10), .A2(MEM_stage_inst_dmem_n17137), .ZN(MEM_stage_inst_dmem_n17126) );
NAND2_X1 MEM_stage_inst_dmem_U15199 ( .A1(MEM_stage_inst_dmem_ram_2533), .A2(MEM_stage_inst_dmem_n17136), .ZN(MEM_stage_inst_dmem_n17127) );
NAND2_X1 MEM_stage_inst_dmem_U15198 ( .A1(MEM_stage_inst_dmem_n17125), .A2(MEM_stage_inst_dmem_n17124), .ZN(MEM_stage_inst_dmem_n10785) );
NAND2_X1 MEM_stage_inst_dmem_U15197 ( .A1(EX_pipeline_reg_out_11), .A2(MEM_stage_inst_dmem_n17137), .ZN(MEM_stage_inst_dmem_n17124) );
NAND2_X1 MEM_stage_inst_dmem_U15196 ( .A1(MEM_stage_inst_dmem_ram_2534), .A2(MEM_stage_inst_dmem_n17136), .ZN(MEM_stage_inst_dmem_n17125) );
NAND2_X1 MEM_stage_inst_dmem_U15195 ( .A1(MEM_stage_inst_dmem_n17123), .A2(MEM_stage_inst_dmem_n17122), .ZN(MEM_stage_inst_dmem_n10786) );
NAND2_X1 MEM_stage_inst_dmem_U15194 ( .A1(EX_pipeline_reg_out_12), .A2(MEM_stage_inst_dmem_n17137), .ZN(MEM_stage_inst_dmem_n17122) );
NAND2_X1 MEM_stage_inst_dmem_U15193 ( .A1(MEM_stage_inst_dmem_ram_2535), .A2(MEM_stage_inst_dmem_n17136), .ZN(MEM_stage_inst_dmem_n17123) );
NAND2_X1 MEM_stage_inst_dmem_U15192 ( .A1(MEM_stage_inst_dmem_n17121), .A2(MEM_stage_inst_dmem_n17120), .ZN(MEM_stage_inst_dmem_n10787) );
NAND2_X1 MEM_stage_inst_dmem_U15191 ( .A1(EX_pipeline_reg_out_13), .A2(MEM_stage_inst_dmem_n17137), .ZN(MEM_stage_inst_dmem_n17120) );
NAND2_X1 MEM_stage_inst_dmem_U15190 ( .A1(MEM_stage_inst_dmem_ram_2536), .A2(MEM_stage_inst_dmem_n17136), .ZN(MEM_stage_inst_dmem_n17121) );
NAND2_X1 MEM_stage_inst_dmem_U15189 ( .A1(MEM_stage_inst_dmem_n17119), .A2(MEM_stage_inst_dmem_n17118), .ZN(MEM_stage_inst_dmem_n10788) );
NAND2_X1 MEM_stage_inst_dmem_U15188 ( .A1(EX_pipeline_reg_out_14), .A2(MEM_stage_inst_dmem_n17137), .ZN(MEM_stage_inst_dmem_n17118) );
NAND2_X1 MEM_stage_inst_dmem_U15187 ( .A1(MEM_stage_inst_dmem_ram_2537), .A2(MEM_stage_inst_dmem_n17136), .ZN(MEM_stage_inst_dmem_n17119) );
NAND2_X1 MEM_stage_inst_dmem_U15186 ( .A1(MEM_stage_inst_dmem_n17117), .A2(MEM_stage_inst_dmem_n17116), .ZN(MEM_stage_inst_dmem_n10789) );
NAND2_X1 MEM_stage_inst_dmem_U15185 ( .A1(EX_pipeline_reg_out_15), .A2(MEM_stage_inst_dmem_n17137), .ZN(MEM_stage_inst_dmem_n17116) );
NAND2_X1 MEM_stage_inst_dmem_U15184 ( .A1(MEM_stage_inst_dmem_ram_2538), .A2(MEM_stage_inst_dmem_n17136), .ZN(MEM_stage_inst_dmem_n17117) );
NAND2_X1 MEM_stage_inst_dmem_U15183 ( .A1(MEM_stage_inst_dmem_n17115), .A2(MEM_stage_inst_dmem_n17114), .ZN(MEM_stage_inst_dmem_n10790) );
NAND2_X1 MEM_stage_inst_dmem_U15182 ( .A1(EX_pipeline_reg_out_16), .A2(MEM_stage_inst_dmem_n17137), .ZN(MEM_stage_inst_dmem_n17114) );
NAND2_X1 MEM_stage_inst_dmem_U15181 ( .A1(MEM_stage_inst_dmem_ram_2539), .A2(MEM_stage_inst_dmem_n17136), .ZN(MEM_stage_inst_dmem_n17115) );
NAND2_X1 MEM_stage_inst_dmem_U15180 ( .A1(MEM_stage_inst_dmem_n17113), .A2(MEM_stage_inst_dmem_n17112), .ZN(MEM_stage_inst_dmem_n10791) );
NAND2_X1 MEM_stage_inst_dmem_U15179 ( .A1(EX_pipeline_reg_out_17), .A2(MEM_stage_inst_dmem_n17137), .ZN(MEM_stage_inst_dmem_n17112) );
NAND2_X1 MEM_stage_inst_dmem_U15178 ( .A1(MEM_stage_inst_dmem_ram_2540), .A2(MEM_stage_inst_dmem_n17136), .ZN(MEM_stage_inst_dmem_n17113) );
NAND2_X1 MEM_stage_inst_dmem_U15177 ( .A1(MEM_stage_inst_dmem_n17111), .A2(MEM_stage_inst_dmem_n17110), .ZN(MEM_stage_inst_dmem_n10792) );
NAND2_X1 MEM_stage_inst_dmem_U15176 ( .A1(EX_pipeline_reg_out_18), .A2(MEM_stage_inst_dmem_n17137), .ZN(MEM_stage_inst_dmem_n17110) );
NAND2_X1 MEM_stage_inst_dmem_U15175 ( .A1(MEM_stage_inst_dmem_ram_2541), .A2(MEM_stage_inst_dmem_n17136), .ZN(MEM_stage_inst_dmem_n17111) );
NAND2_X1 MEM_stage_inst_dmem_U15174 ( .A1(MEM_stage_inst_dmem_n17109), .A2(MEM_stage_inst_dmem_n17108), .ZN(MEM_stage_inst_dmem_n10793) );
NAND2_X1 MEM_stage_inst_dmem_U15173 ( .A1(EX_pipeline_reg_out_19), .A2(MEM_stage_inst_dmem_n17137), .ZN(MEM_stage_inst_dmem_n17108) );
NAND2_X1 MEM_stage_inst_dmem_U15172 ( .A1(MEM_stage_inst_dmem_ram_2542), .A2(MEM_stage_inst_dmem_n17136), .ZN(MEM_stage_inst_dmem_n17109) );
NAND2_X1 MEM_stage_inst_dmem_U15171 ( .A1(MEM_stage_inst_dmem_n17107), .A2(MEM_stage_inst_dmem_n17106), .ZN(MEM_stage_inst_dmem_n10794) );
NAND2_X1 MEM_stage_inst_dmem_U15170 ( .A1(EX_pipeline_reg_out_20), .A2(MEM_stage_inst_dmem_n17137), .ZN(MEM_stage_inst_dmem_n17106) );
INV_X1 MEM_stage_inst_dmem_U15169 ( .A(MEM_stage_inst_dmem_n17136), .ZN(MEM_stage_inst_dmem_n17137) );
NAND2_X1 MEM_stage_inst_dmem_U15168 ( .A1(MEM_stage_inst_dmem_ram_2543), .A2(MEM_stage_inst_dmem_n17136), .ZN(MEM_stage_inst_dmem_n17107) );
NAND2_X1 MEM_stage_inst_dmem_U15167 ( .A1(MEM_stage_inst_dmem_n20969), .A2(MEM_stage_inst_dmem_n17582), .ZN(MEM_stage_inst_dmem_n17136) );
NAND2_X1 MEM_stage_inst_dmem_U15166 ( .A1(MEM_stage_inst_dmem_n17105), .A2(MEM_stage_inst_dmem_n17104), .ZN(MEM_stage_inst_dmem_n10795) );
NAND2_X1 MEM_stage_inst_dmem_U15165 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n17103), .ZN(MEM_stage_inst_dmem_n17104) );
NAND2_X1 MEM_stage_inst_dmem_U15164 ( .A1(MEM_stage_inst_dmem_ram_2544), .A2(MEM_stage_inst_dmem_n17102), .ZN(MEM_stage_inst_dmem_n17105) );
NAND2_X1 MEM_stage_inst_dmem_U15163 ( .A1(MEM_stage_inst_dmem_n17101), .A2(MEM_stage_inst_dmem_n17100), .ZN(MEM_stage_inst_dmem_n10796) );
NAND2_X1 MEM_stage_inst_dmem_U15162 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n17103), .ZN(MEM_stage_inst_dmem_n17100) );
NAND2_X1 MEM_stage_inst_dmem_U15161 ( .A1(MEM_stage_inst_dmem_ram_2545), .A2(MEM_stage_inst_dmem_n17102), .ZN(MEM_stage_inst_dmem_n17101) );
NAND2_X1 MEM_stage_inst_dmem_U15160 ( .A1(MEM_stage_inst_dmem_n17099), .A2(MEM_stage_inst_dmem_n17098), .ZN(MEM_stage_inst_dmem_n10797) );
NAND2_X1 MEM_stage_inst_dmem_U15159 ( .A1(MEM_stage_inst_dmem_n18027), .A2(MEM_stage_inst_dmem_n17103), .ZN(MEM_stage_inst_dmem_n17098) );
NAND2_X1 MEM_stage_inst_dmem_U15158 ( .A1(MEM_stage_inst_dmem_ram_2546), .A2(MEM_stage_inst_dmem_n17102), .ZN(MEM_stage_inst_dmem_n17099) );
NAND2_X1 MEM_stage_inst_dmem_U15157 ( .A1(MEM_stage_inst_dmem_n17097), .A2(MEM_stage_inst_dmem_n17096), .ZN(MEM_stage_inst_dmem_n10798) );
NAND2_X1 MEM_stage_inst_dmem_U15156 ( .A1(EX_pipeline_reg_out_8), .A2(MEM_stage_inst_dmem_n17103), .ZN(MEM_stage_inst_dmem_n17096) );
NAND2_X1 MEM_stage_inst_dmem_U15155 ( .A1(MEM_stage_inst_dmem_ram_2547), .A2(MEM_stage_inst_dmem_n17102), .ZN(MEM_stage_inst_dmem_n17097) );
NAND2_X1 MEM_stage_inst_dmem_U15154 ( .A1(MEM_stage_inst_dmem_n17095), .A2(MEM_stage_inst_dmem_n17094), .ZN(MEM_stage_inst_dmem_n10799) );
NAND2_X1 MEM_stage_inst_dmem_U15153 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n17103), .ZN(MEM_stage_inst_dmem_n17094) );
NAND2_X1 MEM_stage_inst_dmem_U15152 ( .A1(MEM_stage_inst_dmem_ram_2548), .A2(MEM_stage_inst_dmem_n17102), .ZN(MEM_stage_inst_dmem_n17095) );
NAND2_X1 MEM_stage_inst_dmem_U15151 ( .A1(MEM_stage_inst_dmem_n17093), .A2(MEM_stage_inst_dmem_n17092), .ZN(MEM_stage_inst_dmem_n10800) );
NAND2_X1 MEM_stage_inst_dmem_U15150 ( .A1(EX_pipeline_reg_out_10), .A2(MEM_stage_inst_dmem_n17103), .ZN(MEM_stage_inst_dmem_n17092) );
NAND2_X1 MEM_stage_inst_dmem_U15149 ( .A1(MEM_stage_inst_dmem_ram_2549), .A2(MEM_stage_inst_dmem_n17102), .ZN(MEM_stage_inst_dmem_n17093) );
NAND2_X1 MEM_stage_inst_dmem_U15148 ( .A1(MEM_stage_inst_dmem_n17091), .A2(MEM_stage_inst_dmem_n17090), .ZN(MEM_stage_inst_dmem_n10801) );
NAND2_X1 MEM_stage_inst_dmem_U15147 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n17103), .ZN(MEM_stage_inst_dmem_n17090) );
NAND2_X1 MEM_stage_inst_dmem_U15146 ( .A1(MEM_stage_inst_dmem_ram_2550), .A2(MEM_stage_inst_dmem_n17102), .ZN(MEM_stage_inst_dmem_n17091) );
NAND2_X1 MEM_stage_inst_dmem_U15145 ( .A1(MEM_stage_inst_dmem_n17089), .A2(MEM_stage_inst_dmem_n17088), .ZN(MEM_stage_inst_dmem_n10802) );
NAND2_X1 MEM_stage_inst_dmem_U15144 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n17103), .ZN(MEM_stage_inst_dmem_n17088) );
NAND2_X1 MEM_stage_inst_dmem_U15143 ( .A1(MEM_stage_inst_dmem_ram_2551), .A2(MEM_stage_inst_dmem_n17102), .ZN(MEM_stage_inst_dmem_n17089) );
NAND2_X1 MEM_stage_inst_dmem_U15142 ( .A1(MEM_stage_inst_dmem_n17087), .A2(MEM_stage_inst_dmem_n17086), .ZN(MEM_stage_inst_dmem_n10803) );
NAND2_X1 MEM_stage_inst_dmem_U15141 ( .A1(MEM_stage_inst_dmem_n18013), .A2(MEM_stage_inst_dmem_n17103), .ZN(MEM_stage_inst_dmem_n17086) );
NAND2_X1 MEM_stage_inst_dmem_U15140 ( .A1(MEM_stage_inst_dmem_ram_2552), .A2(MEM_stage_inst_dmem_n17102), .ZN(MEM_stage_inst_dmem_n17087) );
NAND2_X1 MEM_stage_inst_dmem_U15139 ( .A1(MEM_stage_inst_dmem_n17085), .A2(MEM_stage_inst_dmem_n17084), .ZN(MEM_stage_inst_dmem_n10804) );
NAND2_X1 MEM_stage_inst_dmem_U15138 ( .A1(MEM_stage_inst_dmem_n96), .A2(MEM_stage_inst_dmem_n17103), .ZN(MEM_stage_inst_dmem_n17084) );
NAND2_X1 MEM_stage_inst_dmem_U15137 ( .A1(MEM_stage_inst_dmem_ram_2553), .A2(MEM_stage_inst_dmem_n17102), .ZN(MEM_stage_inst_dmem_n17085) );
NAND2_X1 MEM_stage_inst_dmem_U15136 ( .A1(MEM_stage_inst_dmem_n17083), .A2(MEM_stage_inst_dmem_n17082), .ZN(MEM_stage_inst_dmem_n10805) );
NAND2_X1 MEM_stage_inst_dmem_U15135 ( .A1(MEM_stage_inst_dmem_n18007), .A2(MEM_stage_inst_dmem_n17103), .ZN(MEM_stage_inst_dmem_n17082) );
NAND2_X1 MEM_stage_inst_dmem_U15134 ( .A1(MEM_stage_inst_dmem_ram_2554), .A2(MEM_stage_inst_dmem_n17102), .ZN(MEM_stage_inst_dmem_n17083) );
NAND2_X1 MEM_stage_inst_dmem_U15133 ( .A1(MEM_stage_inst_dmem_n17081), .A2(MEM_stage_inst_dmem_n17080), .ZN(MEM_stage_inst_dmem_n10806) );
NAND2_X1 MEM_stage_inst_dmem_U15132 ( .A1(MEM_stage_inst_dmem_n18004), .A2(MEM_stage_inst_dmem_n17103), .ZN(MEM_stage_inst_dmem_n17080) );
NAND2_X1 MEM_stage_inst_dmem_U15131 ( .A1(MEM_stage_inst_dmem_ram_2555), .A2(MEM_stage_inst_dmem_n17102), .ZN(MEM_stage_inst_dmem_n17081) );
NAND2_X1 MEM_stage_inst_dmem_U15130 ( .A1(MEM_stage_inst_dmem_n17079), .A2(MEM_stage_inst_dmem_n17078), .ZN(MEM_stage_inst_dmem_n10807) );
NAND2_X1 MEM_stage_inst_dmem_U15129 ( .A1(MEM_stage_inst_dmem_n18001), .A2(MEM_stage_inst_dmem_n17103), .ZN(MEM_stage_inst_dmem_n17078) );
NAND2_X1 MEM_stage_inst_dmem_U15128 ( .A1(MEM_stage_inst_dmem_ram_2556), .A2(MEM_stage_inst_dmem_n17102), .ZN(MEM_stage_inst_dmem_n17079) );
NAND2_X1 MEM_stage_inst_dmem_U15127 ( .A1(MEM_stage_inst_dmem_n17077), .A2(MEM_stage_inst_dmem_n17076), .ZN(MEM_stage_inst_dmem_n10808) );
NAND2_X1 MEM_stage_inst_dmem_U15126 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n17103), .ZN(MEM_stage_inst_dmem_n17076) );
NAND2_X1 MEM_stage_inst_dmem_U15125 ( .A1(MEM_stage_inst_dmem_ram_2557), .A2(MEM_stage_inst_dmem_n17102), .ZN(MEM_stage_inst_dmem_n17077) );
NAND2_X1 MEM_stage_inst_dmem_U15124 ( .A1(MEM_stage_inst_dmem_n17075), .A2(MEM_stage_inst_dmem_n17074), .ZN(MEM_stage_inst_dmem_n10809) );
NAND2_X1 MEM_stage_inst_dmem_U15123 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n17103), .ZN(MEM_stage_inst_dmem_n17074) );
NAND2_X1 MEM_stage_inst_dmem_U15122 ( .A1(MEM_stage_inst_dmem_ram_2558), .A2(MEM_stage_inst_dmem_n17102), .ZN(MEM_stage_inst_dmem_n17075) );
NAND2_X1 MEM_stage_inst_dmem_U15121 ( .A1(MEM_stage_inst_dmem_n17073), .A2(MEM_stage_inst_dmem_n17072), .ZN(MEM_stage_inst_dmem_n10810) );
NAND2_X1 MEM_stage_inst_dmem_U15120 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n17103), .ZN(MEM_stage_inst_dmem_n17072) );
NAND2_X1 MEM_stage_inst_dmem_U15119 ( .A1(MEM_stage_inst_dmem_ram_2559), .A2(MEM_stage_inst_dmem_n17102), .ZN(MEM_stage_inst_dmem_n17073) );
NAND2_X1 MEM_stage_inst_dmem_U15118 ( .A1(MEM_stage_inst_dmem_n20934), .A2(MEM_stage_inst_dmem_n17582), .ZN(MEM_stage_inst_dmem_n17102) );
NOR2_X2 MEM_stage_inst_dmem_U15117 ( .A1(MEM_stage_inst_dmem_n17619), .A2(MEM_stage_inst_dmem_n20369), .ZN(MEM_stage_inst_dmem_n17582) );
NAND2_X1 MEM_stage_inst_dmem_U15116 ( .A1(EX_pipeline_reg_out_26), .A2(MEM_stage_inst_dmem_n17618), .ZN(MEM_stage_inst_dmem_n20369) );
NOR2_X1 MEM_stage_inst_dmem_U15115 ( .A1(EX_pipeline_reg_out_29), .A2(n3522), .ZN(MEM_stage_inst_dmem_n17618) );
NAND2_X1 MEM_stage_inst_dmem_U15114 ( .A1(MEM_stage_inst_dmem_n17071), .A2(MEM_stage_inst_dmem_n17070), .ZN(MEM_stage_inst_dmem_n10811) );
NAND2_X1 MEM_stage_inst_dmem_U15113 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n17069), .ZN(MEM_stage_inst_dmem_n17070) );
NAND2_X1 MEM_stage_inst_dmem_U15112 ( .A1(MEM_stage_inst_dmem_ram_1536), .A2(MEM_stage_inst_dmem_n17068), .ZN(MEM_stage_inst_dmem_n17071) );
NAND2_X1 MEM_stage_inst_dmem_U15111 ( .A1(MEM_stage_inst_dmem_n17067), .A2(MEM_stage_inst_dmem_n17066), .ZN(MEM_stage_inst_dmem_n10812) );
NAND2_X1 MEM_stage_inst_dmem_U15110 ( .A1(MEM_stage_inst_dmem_n109), .A2(MEM_stage_inst_dmem_n17069), .ZN(MEM_stage_inst_dmem_n17066) );
NAND2_X1 MEM_stage_inst_dmem_U15109 ( .A1(MEM_stage_inst_dmem_ram_1537), .A2(MEM_stage_inst_dmem_n17068), .ZN(MEM_stage_inst_dmem_n17067) );
NAND2_X1 MEM_stage_inst_dmem_U15108 ( .A1(MEM_stage_inst_dmem_n17065), .A2(MEM_stage_inst_dmem_n17064), .ZN(MEM_stage_inst_dmem_n10813) );
NAND2_X1 MEM_stage_inst_dmem_U15107 ( .A1(MEM_stage_inst_dmem_n18027), .A2(MEM_stage_inst_dmem_n17069), .ZN(MEM_stage_inst_dmem_n17064) );
NAND2_X1 MEM_stage_inst_dmem_U15106 ( .A1(MEM_stage_inst_dmem_ram_1538), .A2(MEM_stage_inst_dmem_n17068), .ZN(MEM_stage_inst_dmem_n17065) );
NAND2_X1 MEM_stage_inst_dmem_U15105 ( .A1(MEM_stage_inst_dmem_n17063), .A2(MEM_stage_inst_dmem_n17062), .ZN(MEM_stage_inst_dmem_n10814) );
NAND2_X1 MEM_stage_inst_dmem_U15104 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n17069), .ZN(MEM_stage_inst_dmem_n17062) );
NAND2_X1 MEM_stage_inst_dmem_U15103 ( .A1(MEM_stage_inst_dmem_ram_1539), .A2(MEM_stage_inst_dmem_n17068), .ZN(MEM_stage_inst_dmem_n17063) );
NAND2_X1 MEM_stage_inst_dmem_U15102 ( .A1(MEM_stage_inst_dmem_n17061), .A2(MEM_stage_inst_dmem_n17060), .ZN(MEM_stage_inst_dmem_n10815) );
NAND2_X1 MEM_stage_inst_dmem_U15101 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n17069), .ZN(MEM_stage_inst_dmem_n17060) );
NAND2_X1 MEM_stage_inst_dmem_U15100 ( .A1(MEM_stage_inst_dmem_ram_1540), .A2(MEM_stage_inst_dmem_n17068), .ZN(MEM_stage_inst_dmem_n17061) );
NAND2_X1 MEM_stage_inst_dmem_U15099 ( .A1(MEM_stage_inst_dmem_n17059), .A2(MEM_stage_inst_dmem_n17058), .ZN(MEM_stage_inst_dmem_n10816) );
NAND2_X1 MEM_stage_inst_dmem_U15098 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n17069), .ZN(MEM_stage_inst_dmem_n17058) );
NAND2_X1 MEM_stage_inst_dmem_U15097 ( .A1(MEM_stage_inst_dmem_ram_1541), .A2(MEM_stage_inst_dmem_n17068), .ZN(MEM_stage_inst_dmem_n17059) );
NAND2_X1 MEM_stage_inst_dmem_U15096 ( .A1(MEM_stage_inst_dmem_n17057), .A2(MEM_stage_inst_dmem_n17056), .ZN(MEM_stage_inst_dmem_n10817) );
NAND2_X1 MEM_stage_inst_dmem_U15095 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n17069), .ZN(MEM_stage_inst_dmem_n17056) );
NAND2_X1 MEM_stage_inst_dmem_U15094 ( .A1(MEM_stage_inst_dmem_ram_1542), .A2(MEM_stage_inst_dmem_n17068), .ZN(MEM_stage_inst_dmem_n17057) );
NAND2_X1 MEM_stage_inst_dmem_U15093 ( .A1(MEM_stage_inst_dmem_n17055), .A2(MEM_stage_inst_dmem_n17054), .ZN(MEM_stage_inst_dmem_n10818) );
NAND2_X1 MEM_stage_inst_dmem_U15092 ( .A1(MEM_stage_inst_dmem_n16777), .A2(MEM_stage_inst_dmem_n17069), .ZN(MEM_stage_inst_dmem_n17054) );
NAND2_X1 MEM_stage_inst_dmem_U15091 ( .A1(MEM_stage_inst_dmem_ram_1543), .A2(MEM_stage_inst_dmem_n17068), .ZN(MEM_stage_inst_dmem_n17055) );
NAND2_X1 MEM_stage_inst_dmem_U15090 ( .A1(MEM_stage_inst_dmem_n17053), .A2(MEM_stage_inst_dmem_n17052), .ZN(MEM_stage_inst_dmem_n10819) );
NAND2_X1 MEM_stage_inst_dmem_U15089 ( .A1(MEM_stage_inst_dmem_n18013), .A2(MEM_stage_inst_dmem_n17069), .ZN(MEM_stage_inst_dmem_n17052) );
NAND2_X1 MEM_stage_inst_dmem_U15088 ( .A1(MEM_stage_inst_dmem_ram_1544), .A2(MEM_stage_inst_dmem_n17068), .ZN(MEM_stage_inst_dmem_n17053) );
NAND2_X1 MEM_stage_inst_dmem_U15087 ( .A1(MEM_stage_inst_dmem_n17051), .A2(MEM_stage_inst_dmem_n17050), .ZN(MEM_stage_inst_dmem_n10820) );
NAND2_X1 MEM_stage_inst_dmem_U15086 ( .A1(MEM_stage_inst_dmem_n96), .A2(MEM_stage_inst_dmem_n17069), .ZN(MEM_stage_inst_dmem_n17050) );
NAND2_X1 MEM_stage_inst_dmem_U15085 ( .A1(MEM_stage_inst_dmem_ram_1545), .A2(MEM_stage_inst_dmem_n17068), .ZN(MEM_stage_inst_dmem_n17051) );
NAND2_X1 MEM_stage_inst_dmem_U15084 ( .A1(MEM_stage_inst_dmem_n17049), .A2(MEM_stage_inst_dmem_n17048), .ZN(MEM_stage_inst_dmem_n10821) );
NAND2_X1 MEM_stage_inst_dmem_U15083 ( .A1(MEM_stage_inst_dmem_n18007), .A2(MEM_stage_inst_dmem_n17069), .ZN(MEM_stage_inst_dmem_n17048) );
NAND2_X1 MEM_stage_inst_dmem_U15082 ( .A1(MEM_stage_inst_dmem_ram_1546), .A2(MEM_stage_inst_dmem_n17068), .ZN(MEM_stage_inst_dmem_n17049) );
NAND2_X1 MEM_stage_inst_dmem_U15081 ( .A1(MEM_stage_inst_dmem_n17047), .A2(MEM_stage_inst_dmem_n17046), .ZN(MEM_stage_inst_dmem_n10822) );
NAND2_X1 MEM_stage_inst_dmem_U15080 ( .A1(MEM_stage_inst_dmem_n18004), .A2(MEM_stage_inst_dmem_n17069), .ZN(MEM_stage_inst_dmem_n17046) );
NAND2_X1 MEM_stage_inst_dmem_U15079 ( .A1(MEM_stage_inst_dmem_ram_1547), .A2(MEM_stage_inst_dmem_n17068), .ZN(MEM_stage_inst_dmem_n17047) );
NAND2_X1 MEM_stage_inst_dmem_U15078 ( .A1(MEM_stage_inst_dmem_n17045), .A2(MEM_stage_inst_dmem_n17044), .ZN(MEM_stage_inst_dmem_n10823) );
NAND2_X1 MEM_stage_inst_dmem_U15077 ( .A1(MEM_stage_inst_dmem_n18001), .A2(MEM_stage_inst_dmem_n17069), .ZN(MEM_stage_inst_dmem_n17044) );
NAND2_X1 MEM_stage_inst_dmem_U15076 ( .A1(MEM_stage_inst_dmem_ram_1548), .A2(MEM_stage_inst_dmem_n17068), .ZN(MEM_stage_inst_dmem_n17045) );
NAND2_X1 MEM_stage_inst_dmem_U15075 ( .A1(MEM_stage_inst_dmem_n17043), .A2(MEM_stage_inst_dmem_n17042), .ZN(MEM_stage_inst_dmem_n10824) );
NAND2_X1 MEM_stage_inst_dmem_U15074 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n17069), .ZN(MEM_stage_inst_dmem_n17042) );
NAND2_X1 MEM_stage_inst_dmem_U15073 ( .A1(MEM_stage_inst_dmem_ram_1549), .A2(MEM_stage_inst_dmem_n17068), .ZN(MEM_stage_inst_dmem_n17043) );
NAND2_X1 MEM_stage_inst_dmem_U15072 ( .A1(MEM_stage_inst_dmem_n17041), .A2(MEM_stage_inst_dmem_n17040), .ZN(MEM_stage_inst_dmem_n10825) );
NAND2_X1 MEM_stage_inst_dmem_U15071 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n17069), .ZN(MEM_stage_inst_dmem_n17040) );
NAND2_X1 MEM_stage_inst_dmem_U15070 ( .A1(MEM_stage_inst_dmem_ram_1550), .A2(MEM_stage_inst_dmem_n17068), .ZN(MEM_stage_inst_dmem_n17041) );
NAND2_X1 MEM_stage_inst_dmem_U15069 ( .A1(MEM_stage_inst_dmem_n17039), .A2(MEM_stage_inst_dmem_n17038), .ZN(MEM_stage_inst_dmem_n10826) );
NAND2_X1 MEM_stage_inst_dmem_U15068 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n17069), .ZN(MEM_stage_inst_dmem_n17038) );
INV_X1 MEM_stage_inst_dmem_U15067 ( .A(MEM_stage_inst_dmem_n17068), .ZN(MEM_stage_inst_dmem_n17069) );
NAND2_X1 MEM_stage_inst_dmem_U15066 ( .A1(MEM_stage_inst_dmem_ram_1551), .A2(MEM_stage_inst_dmem_n17068), .ZN(MEM_stage_inst_dmem_n17039) );
NAND2_X1 MEM_stage_inst_dmem_U15065 ( .A1(MEM_stage_inst_dmem_n21465), .A2(MEM_stage_inst_dmem_n17037), .ZN(MEM_stage_inst_dmem_n17068) );
NAND2_X1 MEM_stage_inst_dmem_U15064 ( .A1(MEM_stage_inst_dmem_n17036), .A2(MEM_stage_inst_dmem_n17035), .ZN(MEM_stage_inst_dmem_n10827) );
NAND2_X1 MEM_stage_inst_dmem_U15063 ( .A1(EX_pipeline_reg_out_5), .A2(MEM_stage_inst_dmem_n17034), .ZN(MEM_stage_inst_dmem_n17035) );
NAND2_X1 MEM_stage_inst_dmem_U15062 ( .A1(MEM_stage_inst_dmem_ram_1552), .A2(MEM_stage_inst_dmem_n17033), .ZN(MEM_stage_inst_dmem_n17036) );
NAND2_X1 MEM_stage_inst_dmem_U15061 ( .A1(MEM_stage_inst_dmem_n17032), .A2(MEM_stage_inst_dmem_n17031), .ZN(MEM_stage_inst_dmem_n10828) );
NAND2_X1 MEM_stage_inst_dmem_U15060 ( .A1(EX_pipeline_reg_out_6), .A2(MEM_stage_inst_dmem_n17034), .ZN(MEM_stage_inst_dmem_n17031) );
NAND2_X1 MEM_stage_inst_dmem_U15059 ( .A1(MEM_stage_inst_dmem_ram_1553), .A2(MEM_stage_inst_dmem_n17033), .ZN(MEM_stage_inst_dmem_n17032) );
NAND2_X1 MEM_stage_inst_dmem_U15058 ( .A1(MEM_stage_inst_dmem_n17030), .A2(MEM_stage_inst_dmem_n17029), .ZN(MEM_stage_inst_dmem_n10829) );
NAND2_X1 MEM_stage_inst_dmem_U15057 ( .A1(EX_pipeline_reg_out_7), .A2(MEM_stage_inst_dmem_n17034), .ZN(MEM_stage_inst_dmem_n17029) );
NAND2_X1 MEM_stage_inst_dmem_U15056 ( .A1(MEM_stage_inst_dmem_ram_1554), .A2(MEM_stage_inst_dmem_n17033), .ZN(MEM_stage_inst_dmem_n17030) );
NAND2_X1 MEM_stage_inst_dmem_U15055 ( .A1(MEM_stage_inst_dmem_n17028), .A2(MEM_stage_inst_dmem_n17027), .ZN(MEM_stage_inst_dmem_n10830) );
NAND2_X1 MEM_stage_inst_dmem_U15054 ( .A1(EX_pipeline_reg_out_8), .A2(MEM_stage_inst_dmem_n17034), .ZN(MEM_stage_inst_dmem_n17027) );
NAND2_X1 MEM_stage_inst_dmem_U15053 ( .A1(MEM_stage_inst_dmem_ram_1555), .A2(MEM_stage_inst_dmem_n17033), .ZN(MEM_stage_inst_dmem_n17028) );
NAND2_X1 MEM_stage_inst_dmem_U15052 ( .A1(MEM_stage_inst_dmem_n17026), .A2(MEM_stage_inst_dmem_n17025), .ZN(MEM_stage_inst_dmem_n10831) );
NAND2_X1 MEM_stage_inst_dmem_U15051 ( .A1(EX_pipeline_reg_out_9), .A2(MEM_stage_inst_dmem_n17034), .ZN(MEM_stage_inst_dmem_n17025) );
NAND2_X1 MEM_stage_inst_dmem_U15050 ( .A1(MEM_stage_inst_dmem_ram_1556), .A2(MEM_stage_inst_dmem_n17033), .ZN(MEM_stage_inst_dmem_n17026) );
NAND2_X1 MEM_stage_inst_dmem_U15049 ( .A1(MEM_stage_inst_dmem_n17024), .A2(MEM_stage_inst_dmem_n17023), .ZN(MEM_stage_inst_dmem_n10832) );
NAND2_X1 MEM_stage_inst_dmem_U15048 ( .A1(EX_pipeline_reg_out_10), .A2(MEM_stage_inst_dmem_n17034), .ZN(MEM_stage_inst_dmem_n17023) );
NAND2_X1 MEM_stage_inst_dmem_U15047 ( .A1(MEM_stage_inst_dmem_ram_1557), .A2(MEM_stage_inst_dmem_n17033), .ZN(MEM_stage_inst_dmem_n17024) );
NAND2_X1 MEM_stage_inst_dmem_U15046 ( .A1(MEM_stage_inst_dmem_n17022), .A2(MEM_stage_inst_dmem_n17021), .ZN(MEM_stage_inst_dmem_n10833) );
NAND2_X1 MEM_stage_inst_dmem_U15045 ( .A1(EX_pipeline_reg_out_11), .A2(MEM_stage_inst_dmem_n17034), .ZN(MEM_stage_inst_dmem_n17021) );
NAND2_X1 MEM_stage_inst_dmem_U15044 ( .A1(MEM_stage_inst_dmem_ram_1558), .A2(MEM_stage_inst_dmem_n17033), .ZN(MEM_stage_inst_dmem_n17022) );
NAND2_X1 MEM_stage_inst_dmem_U15043 ( .A1(MEM_stage_inst_dmem_n17020), .A2(MEM_stage_inst_dmem_n17019), .ZN(MEM_stage_inst_dmem_n10834) );
NAND2_X1 MEM_stage_inst_dmem_U15042 ( .A1(EX_pipeline_reg_out_12), .A2(MEM_stage_inst_dmem_n17034), .ZN(MEM_stage_inst_dmem_n17019) );
NAND2_X1 MEM_stage_inst_dmem_U15041 ( .A1(MEM_stage_inst_dmem_ram_1559), .A2(MEM_stage_inst_dmem_n17033), .ZN(MEM_stage_inst_dmem_n17020) );
NAND2_X1 MEM_stage_inst_dmem_U15040 ( .A1(MEM_stage_inst_dmem_n17018), .A2(MEM_stage_inst_dmem_n17017), .ZN(MEM_stage_inst_dmem_n10835) );
NAND2_X1 MEM_stage_inst_dmem_U15039 ( .A1(EX_pipeline_reg_out_13), .A2(MEM_stage_inst_dmem_n17034), .ZN(MEM_stage_inst_dmem_n17017) );
NAND2_X1 MEM_stage_inst_dmem_U15038 ( .A1(MEM_stage_inst_dmem_ram_1560), .A2(MEM_stage_inst_dmem_n17033), .ZN(MEM_stage_inst_dmem_n17018) );
NAND2_X1 MEM_stage_inst_dmem_U15037 ( .A1(MEM_stage_inst_dmem_n17016), .A2(MEM_stage_inst_dmem_n17015), .ZN(MEM_stage_inst_dmem_n10836) );
NAND2_X1 MEM_stage_inst_dmem_U15036 ( .A1(EX_pipeline_reg_out_14), .A2(MEM_stage_inst_dmem_n17034), .ZN(MEM_stage_inst_dmem_n17015) );
NAND2_X1 MEM_stage_inst_dmem_U15035 ( .A1(MEM_stage_inst_dmem_ram_1561), .A2(MEM_stage_inst_dmem_n17033), .ZN(MEM_stage_inst_dmem_n17016) );
NAND2_X1 MEM_stage_inst_dmem_U15034 ( .A1(MEM_stage_inst_dmem_n17014), .A2(MEM_stage_inst_dmem_n17013), .ZN(MEM_stage_inst_dmem_n10837) );
NAND2_X1 MEM_stage_inst_dmem_U15033 ( .A1(EX_pipeline_reg_out_15), .A2(MEM_stage_inst_dmem_n17034), .ZN(MEM_stage_inst_dmem_n17013) );
NAND2_X1 MEM_stage_inst_dmem_U15032 ( .A1(MEM_stage_inst_dmem_ram_1562), .A2(MEM_stage_inst_dmem_n17033), .ZN(MEM_stage_inst_dmem_n17014) );
NAND2_X1 MEM_stage_inst_dmem_U15031 ( .A1(MEM_stage_inst_dmem_n17012), .A2(MEM_stage_inst_dmem_n17011), .ZN(MEM_stage_inst_dmem_n10838) );
NAND2_X1 MEM_stage_inst_dmem_U15030 ( .A1(EX_pipeline_reg_out_16), .A2(MEM_stage_inst_dmem_n17034), .ZN(MEM_stage_inst_dmem_n17011) );
NAND2_X1 MEM_stage_inst_dmem_U15029 ( .A1(MEM_stage_inst_dmem_ram_1563), .A2(MEM_stage_inst_dmem_n17033), .ZN(MEM_stage_inst_dmem_n17012) );
NAND2_X1 MEM_stage_inst_dmem_U15028 ( .A1(MEM_stage_inst_dmem_n17010), .A2(MEM_stage_inst_dmem_n17009), .ZN(MEM_stage_inst_dmem_n10839) );
NAND2_X1 MEM_stage_inst_dmem_U15027 ( .A1(EX_pipeline_reg_out_17), .A2(MEM_stage_inst_dmem_n17034), .ZN(MEM_stage_inst_dmem_n17009) );
NAND2_X1 MEM_stage_inst_dmem_U15026 ( .A1(MEM_stage_inst_dmem_ram_1564), .A2(MEM_stage_inst_dmem_n17033), .ZN(MEM_stage_inst_dmem_n17010) );
NAND2_X1 MEM_stage_inst_dmem_U15025 ( .A1(MEM_stage_inst_dmem_n17008), .A2(MEM_stage_inst_dmem_n17007), .ZN(MEM_stage_inst_dmem_n10840) );
NAND2_X1 MEM_stage_inst_dmem_U15024 ( .A1(EX_pipeline_reg_out_18), .A2(MEM_stage_inst_dmem_n17034), .ZN(MEM_stage_inst_dmem_n17007) );
NAND2_X1 MEM_stage_inst_dmem_U15023 ( .A1(MEM_stage_inst_dmem_ram_1565), .A2(MEM_stage_inst_dmem_n17033), .ZN(MEM_stage_inst_dmem_n17008) );
NAND2_X1 MEM_stage_inst_dmem_U15022 ( .A1(MEM_stage_inst_dmem_n17006), .A2(MEM_stage_inst_dmem_n17005), .ZN(MEM_stage_inst_dmem_n10841) );
NAND2_X1 MEM_stage_inst_dmem_U15021 ( .A1(EX_pipeline_reg_out_19), .A2(MEM_stage_inst_dmem_n17034), .ZN(MEM_stage_inst_dmem_n17005) );
NAND2_X1 MEM_stage_inst_dmem_U15020 ( .A1(MEM_stage_inst_dmem_ram_1566), .A2(MEM_stage_inst_dmem_n17033), .ZN(MEM_stage_inst_dmem_n17006) );
NAND2_X1 MEM_stage_inst_dmem_U15019 ( .A1(MEM_stage_inst_dmem_n17004), .A2(MEM_stage_inst_dmem_n17003), .ZN(MEM_stage_inst_dmem_n10842) );
NAND2_X1 MEM_stage_inst_dmem_U15018 ( .A1(EX_pipeline_reg_out_20), .A2(MEM_stage_inst_dmem_n17034), .ZN(MEM_stage_inst_dmem_n17003) );
INV_X1 MEM_stage_inst_dmem_U15017 ( .A(MEM_stage_inst_dmem_n17033), .ZN(MEM_stage_inst_dmem_n17034) );
NAND2_X1 MEM_stage_inst_dmem_U15016 ( .A1(MEM_stage_inst_dmem_ram_1567), .A2(MEM_stage_inst_dmem_n17033), .ZN(MEM_stage_inst_dmem_n17004) );
NAND2_X1 MEM_stage_inst_dmem_U15015 ( .A1(MEM_stage_inst_dmem_n21429), .A2(MEM_stage_inst_dmem_n17037), .ZN(MEM_stage_inst_dmem_n17033) );
NAND2_X1 MEM_stage_inst_dmem_U15014 ( .A1(MEM_stage_inst_dmem_n17002), .A2(MEM_stage_inst_dmem_n17001), .ZN(MEM_stage_inst_dmem_n10843) );
NAND2_X1 MEM_stage_inst_dmem_U15013 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n17000), .ZN(MEM_stage_inst_dmem_n17001) );
NAND2_X1 MEM_stage_inst_dmem_U15012 ( .A1(MEM_stage_inst_dmem_ram_1568), .A2(MEM_stage_inst_dmem_n16999), .ZN(MEM_stage_inst_dmem_n17002) );
NAND2_X1 MEM_stage_inst_dmem_U15011 ( .A1(MEM_stage_inst_dmem_n16998), .A2(MEM_stage_inst_dmem_n16997), .ZN(MEM_stage_inst_dmem_n10844) );
NAND2_X1 MEM_stage_inst_dmem_U15010 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n17000), .ZN(MEM_stage_inst_dmem_n16997) );
NAND2_X1 MEM_stage_inst_dmem_U15009 ( .A1(MEM_stage_inst_dmem_ram_1569), .A2(MEM_stage_inst_dmem_n16999), .ZN(MEM_stage_inst_dmem_n16998) );
NAND2_X1 MEM_stage_inst_dmem_U15008 ( .A1(MEM_stage_inst_dmem_n16996), .A2(MEM_stage_inst_dmem_n16995), .ZN(MEM_stage_inst_dmem_n10845) );
NAND2_X1 MEM_stage_inst_dmem_U15007 ( .A1(MEM_stage_inst_dmem_n18027), .A2(MEM_stage_inst_dmem_n17000), .ZN(MEM_stage_inst_dmem_n16995) );
NAND2_X1 MEM_stage_inst_dmem_U15006 ( .A1(MEM_stage_inst_dmem_ram_1570), .A2(MEM_stage_inst_dmem_n16999), .ZN(MEM_stage_inst_dmem_n16996) );
NAND2_X1 MEM_stage_inst_dmem_U15005 ( .A1(MEM_stage_inst_dmem_n16994), .A2(MEM_stage_inst_dmem_n16993), .ZN(MEM_stage_inst_dmem_n10846) );
NAND2_X1 MEM_stage_inst_dmem_U15004 ( .A1(MEM_stage_inst_dmem_n13064), .A2(MEM_stage_inst_dmem_n17000), .ZN(MEM_stage_inst_dmem_n16993) );
NAND2_X1 MEM_stage_inst_dmem_U15003 ( .A1(MEM_stage_inst_dmem_ram_1571), .A2(MEM_stage_inst_dmem_n16999), .ZN(MEM_stage_inst_dmem_n16994) );
NAND2_X1 MEM_stage_inst_dmem_U15002 ( .A1(MEM_stage_inst_dmem_n16992), .A2(MEM_stage_inst_dmem_n16991), .ZN(MEM_stage_inst_dmem_n10847) );
NAND2_X1 MEM_stage_inst_dmem_U15001 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n17000), .ZN(MEM_stage_inst_dmem_n16991) );
NAND2_X1 MEM_stage_inst_dmem_U15000 ( .A1(MEM_stage_inst_dmem_ram_1572), .A2(MEM_stage_inst_dmem_n16999), .ZN(MEM_stage_inst_dmem_n16992) );
NAND2_X1 MEM_stage_inst_dmem_U14999 ( .A1(MEM_stage_inst_dmem_n16990), .A2(MEM_stage_inst_dmem_n16989), .ZN(MEM_stage_inst_dmem_n10848) );
NAND2_X1 MEM_stage_inst_dmem_U14998 ( .A1(MEM_stage_inst_dmem_n13059), .A2(MEM_stage_inst_dmem_n17000), .ZN(MEM_stage_inst_dmem_n16989) );
NAND2_X1 MEM_stage_inst_dmem_U14997 ( .A1(MEM_stage_inst_dmem_ram_1573), .A2(MEM_stage_inst_dmem_n16999), .ZN(MEM_stage_inst_dmem_n16990) );
NAND2_X1 MEM_stage_inst_dmem_U14996 ( .A1(MEM_stage_inst_dmem_n16988), .A2(MEM_stage_inst_dmem_n16987), .ZN(MEM_stage_inst_dmem_n10849) );
NAND2_X1 MEM_stage_inst_dmem_U14995 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n17000), .ZN(MEM_stage_inst_dmem_n16987) );
NAND2_X1 MEM_stage_inst_dmem_U14994 ( .A1(MEM_stage_inst_dmem_ram_1574), .A2(MEM_stage_inst_dmem_n16999), .ZN(MEM_stage_inst_dmem_n16988) );
NAND2_X1 MEM_stage_inst_dmem_U14993 ( .A1(MEM_stage_inst_dmem_n16986), .A2(MEM_stage_inst_dmem_n16985), .ZN(MEM_stage_inst_dmem_n10850) );
NAND2_X1 MEM_stage_inst_dmem_U14992 ( .A1(MEM_stage_inst_dmem_n16361), .A2(MEM_stage_inst_dmem_n17000), .ZN(MEM_stage_inst_dmem_n16985) );
NAND2_X1 MEM_stage_inst_dmem_U14991 ( .A1(MEM_stage_inst_dmem_ram_1575), .A2(MEM_stage_inst_dmem_n16999), .ZN(MEM_stage_inst_dmem_n16986) );
NAND2_X1 MEM_stage_inst_dmem_U14990 ( .A1(MEM_stage_inst_dmem_n16984), .A2(MEM_stage_inst_dmem_n16983), .ZN(MEM_stage_inst_dmem_n10851) );
NAND2_X1 MEM_stage_inst_dmem_U14989 ( .A1(MEM_stage_inst_dmem_n18013), .A2(MEM_stage_inst_dmem_n17000), .ZN(MEM_stage_inst_dmem_n16983) );
NAND2_X1 MEM_stage_inst_dmem_U14988 ( .A1(MEM_stage_inst_dmem_ram_1576), .A2(MEM_stage_inst_dmem_n16999), .ZN(MEM_stage_inst_dmem_n16984) );
NAND2_X1 MEM_stage_inst_dmem_U14987 ( .A1(MEM_stage_inst_dmem_n16982), .A2(MEM_stage_inst_dmem_n16981), .ZN(MEM_stage_inst_dmem_n10852) );
NAND2_X1 MEM_stage_inst_dmem_U14986 ( .A1(MEM_stage_inst_dmem_n96), .A2(MEM_stage_inst_dmem_n17000), .ZN(MEM_stage_inst_dmem_n16981) );
NAND2_X1 MEM_stage_inst_dmem_U14985 ( .A1(MEM_stage_inst_dmem_ram_1577), .A2(MEM_stage_inst_dmem_n16999), .ZN(MEM_stage_inst_dmem_n16982) );
NAND2_X1 MEM_stage_inst_dmem_U14984 ( .A1(MEM_stage_inst_dmem_n16980), .A2(MEM_stage_inst_dmem_n16979), .ZN(MEM_stage_inst_dmem_n10853) );
NAND2_X1 MEM_stage_inst_dmem_U14983 ( .A1(MEM_stage_inst_dmem_n18007), .A2(MEM_stage_inst_dmem_n17000), .ZN(MEM_stage_inst_dmem_n16979) );
NAND2_X1 MEM_stage_inst_dmem_U14982 ( .A1(MEM_stage_inst_dmem_ram_1578), .A2(MEM_stage_inst_dmem_n16999), .ZN(MEM_stage_inst_dmem_n16980) );
NAND2_X1 MEM_stage_inst_dmem_U14981 ( .A1(MEM_stage_inst_dmem_n16978), .A2(MEM_stage_inst_dmem_n16977), .ZN(MEM_stage_inst_dmem_n10854) );
NAND2_X1 MEM_stage_inst_dmem_U14980 ( .A1(MEM_stage_inst_dmem_n18004), .A2(MEM_stage_inst_dmem_n17000), .ZN(MEM_stage_inst_dmem_n16977) );
NAND2_X1 MEM_stage_inst_dmem_U14979 ( .A1(MEM_stage_inst_dmem_ram_1579), .A2(MEM_stage_inst_dmem_n16999), .ZN(MEM_stage_inst_dmem_n16978) );
NAND2_X1 MEM_stage_inst_dmem_U14978 ( .A1(MEM_stage_inst_dmem_n16976), .A2(MEM_stage_inst_dmem_n16975), .ZN(MEM_stage_inst_dmem_n10855) );
NAND2_X1 MEM_stage_inst_dmem_U14977 ( .A1(MEM_stage_inst_dmem_n18001), .A2(MEM_stage_inst_dmem_n17000), .ZN(MEM_stage_inst_dmem_n16975) );
NAND2_X1 MEM_stage_inst_dmem_U14976 ( .A1(MEM_stage_inst_dmem_ram_1580), .A2(MEM_stage_inst_dmem_n16999), .ZN(MEM_stage_inst_dmem_n16976) );
NAND2_X1 MEM_stage_inst_dmem_U14975 ( .A1(MEM_stage_inst_dmem_n16974), .A2(MEM_stage_inst_dmem_n16973), .ZN(MEM_stage_inst_dmem_n10856) );
NAND2_X1 MEM_stage_inst_dmem_U14974 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n17000), .ZN(MEM_stage_inst_dmem_n16973) );
NAND2_X1 MEM_stage_inst_dmem_U14973 ( .A1(MEM_stage_inst_dmem_ram_1581), .A2(MEM_stage_inst_dmem_n16999), .ZN(MEM_stage_inst_dmem_n16974) );
NAND2_X1 MEM_stage_inst_dmem_U14972 ( .A1(MEM_stage_inst_dmem_n16972), .A2(MEM_stage_inst_dmem_n16971), .ZN(MEM_stage_inst_dmem_n10857) );
NAND2_X1 MEM_stage_inst_dmem_U14971 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n17000), .ZN(MEM_stage_inst_dmem_n16971) );
NAND2_X1 MEM_stage_inst_dmem_U14970 ( .A1(MEM_stage_inst_dmem_ram_1582), .A2(MEM_stage_inst_dmem_n16999), .ZN(MEM_stage_inst_dmem_n16972) );
NAND2_X1 MEM_stage_inst_dmem_U14969 ( .A1(MEM_stage_inst_dmem_n16970), .A2(MEM_stage_inst_dmem_n16969), .ZN(MEM_stage_inst_dmem_n10858) );
NAND2_X1 MEM_stage_inst_dmem_U14968 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n17000), .ZN(MEM_stage_inst_dmem_n16969) );
INV_X1 MEM_stage_inst_dmem_U14967 ( .A(MEM_stage_inst_dmem_n16999), .ZN(MEM_stage_inst_dmem_n17000) );
NAND2_X1 MEM_stage_inst_dmem_U14966 ( .A1(MEM_stage_inst_dmem_ram_1583), .A2(MEM_stage_inst_dmem_n16999), .ZN(MEM_stage_inst_dmem_n16970) );
NAND2_X1 MEM_stage_inst_dmem_U14965 ( .A1(MEM_stage_inst_dmem_n21394), .A2(MEM_stage_inst_dmem_n17037), .ZN(MEM_stage_inst_dmem_n16999) );
NAND2_X1 MEM_stage_inst_dmem_U14964 ( .A1(MEM_stage_inst_dmem_n16968), .A2(MEM_stage_inst_dmem_n16967), .ZN(MEM_stage_inst_dmem_n10859) );
NAND2_X1 MEM_stage_inst_dmem_U14963 ( .A1(EX_pipeline_reg_out_5), .A2(MEM_stage_inst_dmem_n16966), .ZN(MEM_stage_inst_dmem_n16967) );
NAND2_X1 MEM_stage_inst_dmem_U14962 ( .A1(MEM_stage_inst_dmem_ram_1584), .A2(MEM_stage_inst_dmem_n16965), .ZN(MEM_stage_inst_dmem_n16968) );
NAND2_X1 MEM_stage_inst_dmem_U14961 ( .A1(MEM_stage_inst_dmem_n16964), .A2(MEM_stage_inst_dmem_n16963), .ZN(MEM_stage_inst_dmem_n10860) );
NAND2_X1 MEM_stage_inst_dmem_U14960 ( .A1(EX_pipeline_reg_out_6), .A2(MEM_stage_inst_dmem_n16966), .ZN(MEM_stage_inst_dmem_n16963) );
NAND2_X1 MEM_stage_inst_dmem_U14959 ( .A1(MEM_stage_inst_dmem_ram_1585), .A2(MEM_stage_inst_dmem_n16965), .ZN(MEM_stage_inst_dmem_n16964) );
NAND2_X1 MEM_stage_inst_dmem_U14958 ( .A1(MEM_stage_inst_dmem_n16962), .A2(MEM_stage_inst_dmem_n16961), .ZN(MEM_stage_inst_dmem_n10861) );
NAND2_X1 MEM_stage_inst_dmem_U14957 ( .A1(EX_pipeline_reg_out_7), .A2(MEM_stage_inst_dmem_n16966), .ZN(MEM_stage_inst_dmem_n16961) );
NAND2_X1 MEM_stage_inst_dmem_U14956 ( .A1(MEM_stage_inst_dmem_ram_1586), .A2(MEM_stage_inst_dmem_n16965), .ZN(MEM_stage_inst_dmem_n16962) );
NAND2_X1 MEM_stage_inst_dmem_U14955 ( .A1(MEM_stage_inst_dmem_n16960), .A2(MEM_stage_inst_dmem_n16959), .ZN(MEM_stage_inst_dmem_n10862) );
NAND2_X1 MEM_stage_inst_dmem_U14954 ( .A1(EX_pipeline_reg_out_8), .A2(MEM_stage_inst_dmem_n16966), .ZN(MEM_stage_inst_dmem_n16959) );
NAND2_X1 MEM_stage_inst_dmem_U14953 ( .A1(MEM_stage_inst_dmem_ram_1587), .A2(MEM_stage_inst_dmem_n16965), .ZN(MEM_stage_inst_dmem_n16960) );
NAND2_X1 MEM_stage_inst_dmem_U14952 ( .A1(MEM_stage_inst_dmem_n16958), .A2(MEM_stage_inst_dmem_n16957), .ZN(MEM_stage_inst_dmem_n10863) );
NAND2_X1 MEM_stage_inst_dmem_U14951 ( .A1(EX_pipeline_reg_out_9), .A2(MEM_stage_inst_dmem_n16966), .ZN(MEM_stage_inst_dmem_n16957) );
NAND2_X1 MEM_stage_inst_dmem_U14950 ( .A1(MEM_stage_inst_dmem_ram_1588), .A2(MEM_stage_inst_dmem_n16965), .ZN(MEM_stage_inst_dmem_n16958) );
NAND2_X1 MEM_stage_inst_dmem_U14949 ( .A1(MEM_stage_inst_dmem_n16956), .A2(MEM_stage_inst_dmem_n16955), .ZN(MEM_stage_inst_dmem_n10864) );
NAND2_X1 MEM_stage_inst_dmem_U14948 ( .A1(EX_pipeline_reg_out_10), .A2(MEM_stage_inst_dmem_n16966), .ZN(MEM_stage_inst_dmem_n16955) );
NAND2_X1 MEM_stage_inst_dmem_U14947 ( .A1(MEM_stage_inst_dmem_ram_1589), .A2(MEM_stage_inst_dmem_n16965), .ZN(MEM_stage_inst_dmem_n16956) );
NAND2_X1 MEM_stage_inst_dmem_U14946 ( .A1(MEM_stage_inst_dmem_n16954), .A2(MEM_stage_inst_dmem_n16953), .ZN(MEM_stage_inst_dmem_n10865) );
NAND2_X1 MEM_stage_inst_dmem_U14945 ( .A1(EX_pipeline_reg_out_11), .A2(MEM_stage_inst_dmem_n16966), .ZN(MEM_stage_inst_dmem_n16953) );
NAND2_X1 MEM_stage_inst_dmem_U14944 ( .A1(MEM_stage_inst_dmem_ram_1590), .A2(MEM_stage_inst_dmem_n16965), .ZN(MEM_stage_inst_dmem_n16954) );
NAND2_X1 MEM_stage_inst_dmem_U14943 ( .A1(MEM_stage_inst_dmem_n16952), .A2(MEM_stage_inst_dmem_n16951), .ZN(MEM_stage_inst_dmem_n10866) );
NAND2_X1 MEM_stage_inst_dmem_U14942 ( .A1(EX_pipeline_reg_out_12), .A2(MEM_stage_inst_dmem_n16966), .ZN(MEM_stage_inst_dmem_n16951) );
NAND2_X1 MEM_stage_inst_dmem_U14941 ( .A1(MEM_stage_inst_dmem_ram_1591), .A2(MEM_stage_inst_dmem_n16965), .ZN(MEM_stage_inst_dmem_n16952) );
NAND2_X1 MEM_stage_inst_dmem_U14940 ( .A1(MEM_stage_inst_dmem_n16950), .A2(MEM_stage_inst_dmem_n16949), .ZN(MEM_stage_inst_dmem_n10867) );
NAND2_X1 MEM_stage_inst_dmem_U14939 ( .A1(EX_pipeline_reg_out_13), .A2(MEM_stage_inst_dmem_n16966), .ZN(MEM_stage_inst_dmem_n16949) );
NAND2_X1 MEM_stage_inst_dmem_U14938 ( .A1(MEM_stage_inst_dmem_ram_1592), .A2(MEM_stage_inst_dmem_n16965), .ZN(MEM_stage_inst_dmem_n16950) );
NAND2_X1 MEM_stage_inst_dmem_U14937 ( .A1(MEM_stage_inst_dmem_n16948), .A2(MEM_stage_inst_dmem_n16947), .ZN(MEM_stage_inst_dmem_n10868) );
NAND2_X1 MEM_stage_inst_dmem_U14936 ( .A1(EX_pipeline_reg_out_14), .A2(MEM_stage_inst_dmem_n16966), .ZN(MEM_stage_inst_dmem_n16947) );
NAND2_X1 MEM_stage_inst_dmem_U14935 ( .A1(MEM_stage_inst_dmem_ram_1593), .A2(MEM_stage_inst_dmem_n16965), .ZN(MEM_stage_inst_dmem_n16948) );
NAND2_X1 MEM_stage_inst_dmem_U14934 ( .A1(MEM_stage_inst_dmem_n16946), .A2(MEM_stage_inst_dmem_n16945), .ZN(MEM_stage_inst_dmem_n10869) );
NAND2_X1 MEM_stage_inst_dmem_U14933 ( .A1(EX_pipeline_reg_out_15), .A2(MEM_stage_inst_dmem_n16966), .ZN(MEM_stage_inst_dmem_n16945) );
NAND2_X1 MEM_stage_inst_dmem_U14932 ( .A1(MEM_stage_inst_dmem_ram_1594), .A2(MEM_stage_inst_dmem_n16965), .ZN(MEM_stage_inst_dmem_n16946) );
NAND2_X1 MEM_stage_inst_dmem_U14931 ( .A1(MEM_stage_inst_dmem_n16944), .A2(MEM_stage_inst_dmem_n16943), .ZN(MEM_stage_inst_dmem_n10870) );
NAND2_X1 MEM_stage_inst_dmem_U14930 ( .A1(EX_pipeline_reg_out_16), .A2(MEM_stage_inst_dmem_n16966), .ZN(MEM_stage_inst_dmem_n16943) );
NAND2_X1 MEM_stage_inst_dmem_U14929 ( .A1(MEM_stage_inst_dmem_ram_1595), .A2(MEM_stage_inst_dmem_n16965), .ZN(MEM_stage_inst_dmem_n16944) );
NAND2_X1 MEM_stage_inst_dmem_U14928 ( .A1(MEM_stage_inst_dmem_n16942), .A2(MEM_stage_inst_dmem_n16941), .ZN(MEM_stage_inst_dmem_n10871) );
NAND2_X1 MEM_stage_inst_dmem_U14927 ( .A1(EX_pipeline_reg_out_17), .A2(MEM_stage_inst_dmem_n16966), .ZN(MEM_stage_inst_dmem_n16941) );
NAND2_X1 MEM_stage_inst_dmem_U14926 ( .A1(MEM_stage_inst_dmem_ram_1596), .A2(MEM_stage_inst_dmem_n16965), .ZN(MEM_stage_inst_dmem_n16942) );
NAND2_X1 MEM_stage_inst_dmem_U14925 ( .A1(MEM_stage_inst_dmem_n16940), .A2(MEM_stage_inst_dmem_n16939), .ZN(MEM_stage_inst_dmem_n10872) );
NAND2_X1 MEM_stage_inst_dmem_U14924 ( .A1(EX_pipeline_reg_out_18), .A2(MEM_stage_inst_dmem_n16966), .ZN(MEM_stage_inst_dmem_n16939) );
NAND2_X1 MEM_stage_inst_dmem_U14923 ( .A1(MEM_stage_inst_dmem_ram_1597), .A2(MEM_stage_inst_dmem_n16965), .ZN(MEM_stage_inst_dmem_n16940) );
NAND2_X1 MEM_stage_inst_dmem_U14922 ( .A1(MEM_stage_inst_dmem_n16938), .A2(MEM_stage_inst_dmem_n16937), .ZN(MEM_stage_inst_dmem_n10873) );
NAND2_X1 MEM_stage_inst_dmem_U14921 ( .A1(EX_pipeline_reg_out_19), .A2(MEM_stage_inst_dmem_n16966), .ZN(MEM_stage_inst_dmem_n16937) );
NAND2_X1 MEM_stage_inst_dmem_U14920 ( .A1(MEM_stage_inst_dmem_ram_1598), .A2(MEM_stage_inst_dmem_n16965), .ZN(MEM_stage_inst_dmem_n16938) );
NAND2_X1 MEM_stage_inst_dmem_U14919 ( .A1(MEM_stage_inst_dmem_n16936), .A2(MEM_stage_inst_dmem_n16935), .ZN(MEM_stage_inst_dmem_n10874) );
NAND2_X1 MEM_stage_inst_dmem_U14918 ( .A1(EX_pipeline_reg_out_20), .A2(MEM_stage_inst_dmem_n16966), .ZN(MEM_stage_inst_dmem_n16935) );
INV_X1 MEM_stage_inst_dmem_U14917 ( .A(MEM_stage_inst_dmem_n16965), .ZN(MEM_stage_inst_dmem_n16966) );
NAND2_X1 MEM_stage_inst_dmem_U14916 ( .A1(MEM_stage_inst_dmem_ram_1599), .A2(MEM_stage_inst_dmem_n16965), .ZN(MEM_stage_inst_dmem_n16936) );
NAND2_X1 MEM_stage_inst_dmem_U14915 ( .A1(MEM_stage_inst_dmem_n21359), .A2(MEM_stage_inst_dmem_n17037), .ZN(MEM_stage_inst_dmem_n16965) );
NAND2_X1 MEM_stage_inst_dmem_U14914 ( .A1(MEM_stage_inst_dmem_n16934), .A2(MEM_stage_inst_dmem_n16933), .ZN(MEM_stage_inst_dmem_n10875) );
NAND2_X1 MEM_stage_inst_dmem_U14913 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n16932), .ZN(MEM_stage_inst_dmem_n16933) );
NAND2_X1 MEM_stage_inst_dmem_U14912 ( .A1(MEM_stage_inst_dmem_ram_1600), .A2(MEM_stage_inst_dmem_n16931), .ZN(MEM_stage_inst_dmem_n16934) );
NAND2_X1 MEM_stage_inst_dmem_U14911 ( .A1(MEM_stage_inst_dmem_n16930), .A2(MEM_stage_inst_dmem_n16929), .ZN(MEM_stage_inst_dmem_n10876) );
NAND2_X1 MEM_stage_inst_dmem_U14910 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n16932), .ZN(MEM_stage_inst_dmem_n16929) );
NAND2_X1 MEM_stage_inst_dmem_U14909 ( .A1(MEM_stage_inst_dmem_ram_1601), .A2(MEM_stage_inst_dmem_n16931), .ZN(MEM_stage_inst_dmem_n16930) );
NAND2_X1 MEM_stage_inst_dmem_U14908 ( .A1(MEM_stage_inst_dmem_n16928), .A2(MEM_stage_inst_dmem_n16927), .ZN(MEM_stage_inst_dmem_n10877) );
NAND2_X1 MEM_stage_inst_dmem_U14907 ( .A1(MEM_stage_inst_dmem_n18027), .A2(MEM_stage_inst_dmem_n16932), .ZN(MEM_stage_inst_dmem_n16927) );
NAND2_X1 MEM_stage_inst_dmem_U14906 ( .A1(MEM_stage_inst_dmem_ram_1602), .A2(MEM_stage_inst_dmem_n16931), .ZN(MEM_stage_inst_dmem_n16928) );
NAND2_X1 MEM_stage_inst_dmem_U14905 ( .A1(MEM_stage_inst_dmem_n16926), .A2(MEM_stage_inst_dmem_n16925), .ZN(MEM_stage_inst_dmem_n10878) );
NAND2_X1 MEM_stage_inst_dmem_U14904 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n16932), .ZN(MEM_stage_inst_dmem_n16925) );
NAND2_X1 MEM_stage_inst_dmem_U14903 ( .A1(MEM_stage_inst_dmem_ram_1603), .A2(MEM_stage_inst_dmem_n16931), .ZN(MEM_stage_inst_dmem_n16926) );
NAND2_X1 MEM_stage_inst_dmem_U14902 ( .A1(MEM_stage_inst_dmem_n16924), .A2(MEM_stage_inst_dmem_n16923), .ZN(MEM_stage_inst_dmem_n10879) );
NAND2_X1 MEM_stage_inst_dmem_U14901 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n16932), .ZN(MEM_stage_inst_dmem_n16923) );
NAND2_X1 MEM_stage_inst_dmem_U14900 ( .A1(MEM_stage_inst_dmem_ram_1604), .A2(MEM_stage_inst_dmem_n16931), .ZN(MEM_stage_inst_dmem_n16924) );
NAND2_X1 MEM_stage_inst_dmem_U14899 ( .A1(MEM_stage_inst_dmem_n16922), .A2(MEM_stage_inst_dmem_n16921), .ZN(MEM_stage_inst_dmem_n10880) );
NAND2_X1 MEM_stage_inst_dmem_U14898 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n16932), .ZN(MEM_stage_inst_dmem_n16921) );
NAND2_X1 MEM_stage_inst_dmem_U14897 ( .A1(MEM_stage_inst_dmem_ram_1605), .A2(MEM_stage_inst_dmem_n16931), .ZN(MEM_stage_inst_dmem_n16922) );
NAND2_X1 MEM_stage_inst_dmem_U14896 ( .A1(MEM_stage_inst_dmem_n16920), .A2(MEM_stage_inst_dmem_n16919), .ZN(MEM_stage_inst_dmem_n10881) );
NAND2_X1 MEM_stage_inst_dmem_U14895 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n16932), .ZN(MEM_stage_inst_dmem_n16919) );
NAND2_X1 MEM_stage_inst_dmem_U14894 ( .A1(MEM_stage_inst_dmem_ram_1606), .A2(MEM_stage_inst_dmem_n16931), .ZN(MEM_stage_inst_dmem_n16920) );
NAND2_X1 MEM_stage_inst_dmem_U14893 ( .A1(MEM_stage_inst_dmem_n16918), .A2(MEM_stage_inst_dmem_n16917), .ZN(MEM_stage_inst_dmem_n10882) );
NAND2_X1 MEM_stage_inst_dmem_U14892 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n16932), .ZN(MEM_stage_inst_dmem_n16917) );
NAND2_X1 MEM_stage_inst_dmem_U14891 ( .A1(MEM_stage_inst_dmem_ram_1607), .A2(MEM_stage_inst_dmem_n16931), .ZN(MEM_stage_inst_dmem_n16918) );
NAND2_X1 MEM_stage_inst_dmem_U14890 ( .A1(MEM_stage_inst_dmem_n16916), .A2(MEM_stage_inst_dmem_n16915), .ZN(MEM_stage_inst_dmem_n10883) );
NAND2_X1 MEM_stage_inst_dmem_U14889 ( .A1(MEM_stage_inst_dmem_n18013), .A2(MEM_stage_inst_dmem_n16932), .ZN(MEM_stage_inst_dmem_n16915) );
NAND2_X1 MEM_stage_inst_dmem_U14888 ( .A1(MEM_stage_inst_dmem_ram_1608), .A2(MEM_stage_inst_dmem_n16931), .ZN(MEM_stage_inst_dmem_n16916) );
NAND2_X1 MEM_stage_inst_dmem_U14887 ( .A1(MEM_stage_inst_dmem_n16914), .A2(MEM_stage_inst_dmem_n16913), .ZN(MEM_stage_inst_dmem_n10884) );
NAND2_X1 MEM_stage_inst_dmem_U14886 ( .A1(MEM_stage_inst_dmem_n96), .A2(MEM_stage_inst_dmem_n16932), .ZN(MEM_stage_inst_dmem_n16913) );
NAND2_X1 MEM_stage_inst_dmem_U14885 ( .A1(MEM_stage_inst_dmem_ram_1609), .A2(MEM_stage_inst_dmem_n16931), .ZN(MEM_stage_inst_dmem_n16914) );
NAND2_X1 MEM_stage_inst_dmem_U14884 ( .A1(MEM_stage_inst_dmem_n16912), .A2(MEM_stage_inst_dmem_n16911), .ZN(MEM_stage_inst_dmem_n10885) );
NAND2_X1 MEM_stage_inst_dmem_U14883 ( .A1(MEM_stage_inst_dmem_n18007), .A2(MEM_stage_inst_dmem_n16932), .ZN(MEM_stage_inst_dmem_n16911) );
NAND2_X1 MEM_stage_inst_dmem_U14882 ( .A1(MEM_stage_inst_dmem_ram_1610), .A2(MEM_stage_inst_dmem_n16931), .ZN(MEM_stage_inst_dmem_n16912) );
NAND2_X1 MEM_stage_inst_dmem_U14881 ( .A1(MEM_stage_inst_dmem_n16910), .A2(MEM_stage_inst_dmem_n16909), .ZN(MEM_stage_inst_dmem_n10886) );
NAND2_X1 MEM_stage_inst_dmem_U14880 ( .A1(MEM_stage_inst_dmem_n18004), .A2(MEM_stage_inst_dmem_n16932), .ZN(MEM_stage_inst_dmem_n16909) );
NAND2_X1 MEM_stage_inst_dmem_U14879 ( .A1(MEM_stage_inst_dmem_ram_1611), .A2(MEM_stage_inst_dmem_n16931), .ZN(MEM_stage_inst_dmem_n16910) );
NAND2_X1 MEM_stage_inst_dmem_U14878 ( .A1(MEM_stage_inst_dmem_n16908), .A2(MEM_stage_inst_dmem_n16907), .ZN(MEM_stage_inst_dmem_n10887) );
NAND2_X1 MEM_stage_inst_dmem_U14877 ( .A1(MEM_stage_inst_dmem_n18001), .A2(MEM_stage_inst_dmem_n16932), .ZN(MEM_stage_inst_dmem_n16907) );
NAND2_X1 MEM_stage_inst_dmem_U14876 ( .A1(MEM_stage_inst_dmem_ram_1612), .A2(MEM_stage_inst_dmem_n16931), .ZN(MEM_stage_inst_dmem_n16908) );
NAND2_X1 MEM_stage_inst_dmem_U14875 ( .A1(MEM_stage_inst_dmem_n16906), .A2(MEM_stage_inst_dmem_n16905), .ZN(MEM_stage_inst_dmem_n10888) );
NAND2_X1 MEM_stage_inst_dmem_U14874 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n16932), .ZN(MEM_stage_inst_dmem_n16905) );
NAND2_X1 MEM_stage_inst_dmem_U14873 ( .A1(MEM_stage_inst_dmem_ram_1613), .A2(MEM_stage_inst_dmem_n16931), .ZN(MEM_stage_inst_dmem_n16906) );
NAND2_X1 MEM_stage_inst_dmem_U14872 ( .A1(MEM_stage_inst_dmem_n16904), .A2(MEM_stage_inst_dmem_n16903), .ZN(MEM_stage_inst_dmem_n10889) );
NAND2_X1 MEM_stage_inst_dmem_U14871 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n16932), .ZN(MEM_stage_inst_dmem_n16903) );
NAND2_X1 MEM_stage_inst_dmem_U14870 ( .A1(MEM_stage_inst_dmem_ram_1614), .A2(MEM_stage_inst_dmem_n16931), .ZN(MEM_stage_inst_dmem_n16904) );
NAND2_X1 MEM_stage_inst_dmem_U14869 ( .A1(MEM_stage_inst_dmem_n16902), .A2(MEM_stage_inst_dmem_n16901), .ZN(MEM_stage_inst_dmem_n10890) );
NAND2_X1 MEM_stage_inst_dmem_U14868 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n16932), .ZN(MEM_stage_inst_dmem_n16901) );
INV_X1 MEM_stage_inst_dmem_U14867 ( .A(MEM_stage_inst_dmem_n16931), .ZN(MEM_stage_inst_dmem_n16932) );
NAND2_X1 MEM_stage_inst_dmem_U14866 ( .A1(MEM_stage_inst_dmem_ram_1615), .A2(MEM_stage_inst_dmem_n16931), .ZN(MEM_stage_inst_dmem_n16902) );
NAND2_X1 MEM_stage_inst_dmem_U14865 ( .A1(MEM_stage_inst_dmem_n21319), .A2(MEM_stage_inst_dmem_n17037), .ZN(MEM_stage_inst_dmem_n16931) );
NAND2_X1 MEM_stage_inst_dmem_U14864 ( .A1(MEM_stage_inst_dmem_n16900), .A2(MEM_stage_inst_dmem_n16899), .ZN(MEM_stage_inst_dmem_n10891) );
NAND2_X1 MEM_stage_inst_dmem_U14863 ( .A1(EX_pipeline_reg_out_5), .A2(MEM_stage_inst_dmem_n16898), .ZN(MEM_stage_inst_dmem_n16899) );
NAND2_X1 MEM_stage_inst_dmem_U14862 ( .A1(MEM_stage_inst_dmem_ram_1616), .A2(MEM_stage_inst_dmem_n16897), .ZN(MEM_stage_inst_dmem_n16900) );
NAND2_X1 MEM_stage_inst_dmem_U14861 ( .A1(MEM_stage_inst_dmem_n16896), .A2(MEM_stage_inst_dmem_n16895), .ZN(MEM_stage_inst_dmem_n10892) );
NAND2_X1 MEM_stage_inst_dmem_U14860 ( .A1(EX_pipeline_reg_out_6), .A2(MEM_stage_inst_dmem_n16898), .ZN(MEM_stage_inst_dmem_n16895) );
NAND2_X1 MEM_stage_inst_dmem_U14859 ( .A1(MEM_stage_inst_dmem_ram_1617), .A2(MEM_stage_inst_dmem_n16897), .ZN(MEM_stage_inst_dmem_n16896) );
NAND2_X1 MEM_stage_inst_dmem_U14858 ( .A1(MEM_stage_inst_dmem_n16894), .A2(MEM_stage_inst_dmem_n16893), .ZN(MEM_stage_inst_dmem_n10893) );
NAND2_X1 MEM_stage_inst_dmem_U14857 ( .A1(EX_pipeline_reg_out_7), .A2(MEM_stage_inst_dmem_n16898), .ZN(MEM_stage_inst_dmem_n16893) );
NAND2_X1 MEM_stage_inst_dmem_U14856 ( .A1(MEM_stage_inst_dmem_ram_1618), .A2(MEM_stage_inst_dmem_n16897), .ZN(MEM_stage_inst_dmem_n16894) );
NAND2_X1 MEM_stage_inst_dmem_U14855 ( .A1(MEM_stage_inst_dmem_n16892), .A2(MEM_stage_inst_dmem_n16891), .ZN(MEM_stage_inst_dmem_n10894) );
NAND2_X1 MEM_stage_inst_dmem_U14854 ( .A1(EX_pipeline_reg_out_8), .A2(MEM_stage_inst_dmem_n16898), .ZN(MEM_stage_inst_dmem_n16891) );
NAND2_X1 MEM_stage_inst_dmem_U14853 ( .A1(MEM_stage_inst_dmem_ram_1619), .A2(MEM_stage_inst_dmem_n16897), .ZN(MEM_stage_inst_dmem_n16892) );
NAND2_X1 MEM_stage_inst_dmem_U14852 ( .A1(MEM_stage_inst_dmem_n16890), .A2(MEM_stage_inst_dmem_n16889), .ZN(MEM_stage_inst_dmem_n10895) );
NAND2_X1 MEM_stage_inst_dmem_U14851 ( .A1(EX_pipeline_reg_out_9), .A2(MEM_stage_inst_dmem_n16898), .ZN(MEM_stage_inst_dmem_n16889) );
NAND2_X1 MEM_stage_inst_dmem_U14850 ( .A1(MEM_stage_inst_dmem_ram_1620), .A2(MEM_stage_inst_dmem_n16897), .ZN(MEM_stage_inst_dmem_n16890) );
NAND2_X1 MEM_stage_inst_dmem_U14849 ( .A1(MEM_stage_inst_dmem_n16888), .A2(MEM_stage_inst_dmem_n16887), .ZN(MEM_stage_inst_dmem_n10896) );
NAND2_X1 MEM_stage_inst_dmem_U14848 ( .A1(EX_pipeline_reg_out_10), .A2(MEM_stage_inst_dmem_n16898), .ZN(MEM_stage_inst_dmem_n16887) );
NAND2_X1 MEM_stage_inst_dmem_U14847 ( .A1(MEM_stage_inst_dmem_ram_1621), .A2(MEM_stage_inst_dmem_n16897), .ZN(MEM_stage_inst_dmem_n16888) );
NAND2_X1 MEM_stage_inst_dmem_U14846 ( .A1(MEM_stage_inst_dmem_n16886), .A2(MEM_stage_inst_dmem_n16885), .ZN(MEM_stage_inst_dmem_n10897) );
NAND2_X1 MEM_stage_inst_dmem_U14845 ( .A1(EX_pipeline_reg_out_11), .A2(MEM_stage_inst_dmem_n16898), .ZN(MEM_stage_inst_dmem_n16885) );
NAND2_X1 MEM_stage_inst_dmem_U14844 ( .A1(MEM_stage_inst_dmem_ram_1622), .A2(MEM_stage_inst_dmem_n16897), .ZN(MEM_stage_inst_dmem_n16886) );
NAND2_X1 MEM_stage_inst_dmem_U14843 ( .A1(MEM_stage_inst_dmem_n16884), .A2(MEM_stage_inst_dmem_n16883), .ZN(MEM_stage_inst_dmem_n10898) );
NAND2_X1 MEM_stage_inst_dmem_U14842 ( .A1(EX_pipeline_reg_out_12), .A2(MEM_stage_inst_dmem_n16898), .ZN(MEM_stage_inst_dmem_n16883) );
NAND2_X1 MEM_stage_inst_dmem_U14841 ( .A1(MEM_stage_inst_dmem_ram_1623), .A2(MEM_stage_inst_dmem_n16897), .ZN(MEM_stage_inst_dmem_n16884) );
NAND2_X1 MEM_stage_inst_dmem_U14840 ( .A1(MEM_stage_inst_dmem_n16882), .A2(MEM_stage_inst_dmem_n16881), .ZN(MEM_stage_inst_dmem_n10899) );
NAND2_X1 MEM_stage_inst_dmem_U14839 ( .A1(EX_pipeline_reg_out_13), .A2(MEM_stage_inst_dmem_n16898), .ZN(MEM_stage_inst_dmem_n16881) );
NAND2_X1 MEM_stage_inst_dmem_U14838 ( .A1(MEM_stage_inst_dmem_ram_1624), .A2(MEM_stage_inst_dmem_n16897), .ZN(MEM_stage_inst_dmem_n16882) );
NAND2_X1 MEM_stage_inst_dmem_U14837 ( .A1(MEM_stage_inst_dmem_n16880), .A2(MEM_stage_inst_dmem_n16879), .ZN(MEM_stage_inst_dmem_n10900) );
NAND2_X1 MEM_stage_inst_dmem_U14836 ( .A1(EX_pipeline_reg_out_14), .A2(MEM_stage_inst_dmem_n16898), .ZN(MEM_stage_inst_dmem_n16879) );
NAND2_X1 MEM_stage_inst_dmem_U14835 ( .A1(MEM_stage_inst_dmem_ram_1625), .A2(MEM_stage_inst_dmem_n16897), .ZN(MEM_stage_inst_dmem_n16880) );
NAND2_X1 MEM_stage_inst_dmem_U14834 ( .A1(MEM_stage_inst_dmem_n16878), .A2(MEM_stage_inst_dmem_n16877), .ZN(MEM_stage_inst_dmem_n10901) );
NAND2_X1 MEM_stage_inst_dmem_U14833 ( .A1(EX_pipeline_reg_out_15), .A2(MEM_stage_inst_dmem_n16898), .ZN(MEM_stage_inst_dmem_n16877) );
NAND2_X1 MEM_stage_inst_dmem_U14832 ( .A1(MEM_stage_inst_dmem_ram_1626), .A2(MEM_stage_inst_dmem_n16897), .ZN(MEM_stage_inst_dmem_n16878) );
NAND2_X1 MEM_stage_inst_dmem_U14831 ( .A1(MEM_stage_inst_dmem_n16876), .A2(MEM_stage_inst_dmem_n16875), .ZN(MEM_stage_inst_dmem_n10902) );
NAND2_X1 MEM_stage_inst_dmem_U14830 ( .A1(EX_pipeline_reg_out_16), .A2(MEM_stage_inst_dmem_n16898), .ZN(MEM_stage_inst_dmem_n16875) );
NAND2_X1 MEM_stage_inst_dmem_U14829 ( .A1(MEM_stage_inst_dmem_ram_1627), .A2(MEM_stage_inst_dmem_n16897), .ZN(MEM_stage_inst_dmem_n16876) );
NAND2_X1 MEM_stage_inst_dmem_U14828 ( .A1(MEM_stage_inst_dmem_n16874), .A2(MEM_stage_inst_dmem_n16873), .ZN(MEM_stage_inst_dmem_n10903) );
NAND2_X1 MEM_stage_inst_dmem_U14827 ( .A1(EX_pipeline_reg_out_17), .A2(MEM_stage_inst_dmem_n16898), .ZN(MEM_stage_inst_dmem_n16873) );
NAND2_X1 MEM_stage_inst_dmem_U14826 ( .A1(MEM_stage_inst_dmem_ram_1628), .A2(MEM_stage_inst_dmem_n16897), .ZN(MEM_stage_inst_dmem_n16874) );
NAND2_X1 MEM_stage_inst_dmem_U14825 ( .A1(MEM_stage_inst_dmem_n16872), .A2(MEM_stage_inst_dmem_n16871), .ZN(MEM_stage_inst_dmem_n10904) );
NAND2_X1 MEM_stage_inst_dmem_U14824 ( .A1(EX_pipeline_reg_out_18), .A2(MEM_stage_inst_dmem_n16898), .ZN(MEM_stage_inst_dmem_n16871) );
NAND2_X1 MEM_stage_inst_dmem_U14823 ( .A1(MEM_stage_inst_dmem_ram_1629), .A2(MEM_stage_inst_dmem_n16897), .ZN(MEM_stage_inst_dmem_n16872) );
NAND2_X1 MEM_stage_inst_dmem_U14822 ( .A1(MEM_stage_inst_dmem_n16870), .A2(MEM_stage_inst_dmem_n16869), .ZN(MEM_stage_inst_dmem_n10905) );
NAND2_X1 MEM_stage_inst_dmem_U14821 ( .A1(EX_pipeline_reg_out_19), .A2(MEM_stage_inst_dmem_n16898), .ZN(MEM_stage_inst_dmem_n16869) );
NAND2_X1 MEM_stage_inst_dmem_U14820 ( .A1(MEM_stage_inst_dmem_ram_1630), .A2(MEM_stage_inst_dmem_n16897), .ZN(MEM_stage_inst_dmem_n16870) );
NAND2_X1 MEM_stage_inst_dmem_U14819 ( .A1(MEM_stage_inst_dmem_n16868), .A2(MEM_stage_inst_dmem_n16867), .ZN(MEM_stage_inst_dmem_n10906) );
NAND2_X1 MEM_stage_inst_dmem_U14818 ( .A1(EX_pipeline_reg_out_20), .A2(MEM_stage_inst_dmem_n16898), .ZN(MEM_stage_inst_dmem_n16867) );
INV_X1 MEM_stage_inst_dmem_U14817 ( .A(MEM_stage_inst_dmem_n16897), .ZN(MEM_stage_inst_dmem_n16898) );
NAND2_X1 MEM_stage_inst_dmem_U14816 ( .A1(MEM_stage_inst_dmem_ram_1631), .A2(MEM_stage_inst_dmem_n16897), .ZN(MEM_stage_inst_dmem_n16868) );
NAND2_X1 MEM_stage_inst_dmem_U14815 ( .A1(MEM_stage_inst_dmem_n21284), .A2(MEM_stage_inst_dmem_n17037), .ZN(MEM_stage_inst_dmem_n16897) );
NAND2_X1 MEM_stage_inst_dmem_U14814 ( .A1(MEM_stage_inst_dmem_n16866), .A2(MEM_stage_inst_dmem_n16865), .ZN(MEM_stage_inst_dmem_n10907) );
NAND2_X1 MEM_stage_inst_dmem_U14813 ( .A1(EX_pipeline_reg_out_5), .A2(MEM_stage_inst_dmem_n16864), .ZN(MEM_stage_inst_dmem_n16865) );
NAND2_X1 MEM_stage_inst_dmem_U14812 ( .A1(MEM_stage_inst_dmem_ram_1632), .A2(MEM_stage_inst_dmem_n16863), .ZN(MEM_stage_inst_dmem_n16866) );
NAND2_X1 MEM_stage_inst_dmem_U14811 ( .A1(MEM_stage_inst_dmem_n16862), .A2(MEM_stage_inst_dmem_n16861), .ZN(MEM_stage_inst_dmem_n10908) );
NAND2_X1 MEM_stage_inst_dmem_U14810 ( .A1(EX_pipeline_reg_out_6), .A2(MEM_stage_inst_dmem_n16864), .ZN(MEM_stage_inst_dmem_n16861) );
NAND2_X1 MEM_stage_inst_dmem_U14809 ( .A1(MEM_stage_inst_dmem_ram_1633), .A2(MEM_stage_inst_dmem_n16863), .ZN(MEM_stage_inst_dmem_n16862) );
NAND2_X1 MEM_stage_inst_dmem_U14808 ( .A1(MEM_stage_inst_dmem_n16860), .A2(MEM_stage_inst_dmem_n16859), .ZN(MEM_stage_inst_dmem_n10909) );
NAND2_X1 MEM_stage_inst_dmem_U14807 ( .A1(EX_pipeline_reg_out_7), .A2(MEM_stage_inst_dmem_n16864), .ZN(MEM_stage_inst_dmem_n16859) );
NAND2_X1 MEM_stage_inst_dmem_U14806 ( .A1(MEM_stage_inst_dmem_ram_1634), .A2(MEM_stage_inst_dmem_n16863), .ZN(MEM_stage_inst_dmem_n16860) );
NAND2_X1 MEM_stage_inst_dmem_U14805 ( .A1(MEM_stage_inst_dmem_n16858), .A2(MEM_stage_inst_dmem_n16857), .ZN(MEM_stage_inst_dmem_n10910) );
NAND2_X1 MEM_stage_inst_dmem_U14804 ( .A1(EX_pipeline_reg_out_8), .A2(MEM_stage_inst_dmem_n16864), .ZN(MEM_stage_inst_dmem_n16857) );
NAND2_X1 MEM_stage_inst_dmem_U14803 ( .A1(MEM_stage_inst_dmem_ram_1635), .A2(MEM_stage_inst_dmem_n16863), .ZN(MEM_stage_inst_dmem_n16858) );
NAND2_X1 MEM_stage_inst_dmem_U14802 ( .A1(MEM_stage_inst_dmem_n16856), .A2(MEM_stage_inst_dmem_n16855), .ZN(MEM_stage_inst_dmem_n10911) );
NAND2_X1 MEM_stage_inst_dmem_U14801 ( .A1(EX_pipeline_reg_out_9), .A2(MEM_stage_inst_dmem_n16864), .ZN(MEM_stage_inst_dmem_n16855) );
NAND2_X1 MEM_stage_inst_dmem_U14800 ( .A1(MEM_stage_inst_dmem_ram_1636), .A2(MEM_stage_inst_dmem_n16863), .ZN(MEM_stage_inst_dmem_n16856) );
NAND2_X1 MEM_stage_inst_dmem_U14799 ( .A1(MEM_stage_inst_dmem_n16854), .A2(MEM_stage_inst_dmem_n16853), .ZN(MEM_stage_inst_dmem_n10912) );
NAND2_X1 MEM_stage_inst_dmem_U14798 ( .A1(EX_pipeline_reg_out_10), .A2(MEM_stage_inst_dmem_n16864), .ZN(MEM_stage_inst_dmem_n16853) );
NAND2_X1 MEM_stage_inst_dmem_U14797 ( .A1(MEM_stage_inst_dmem_ram_1637), .A2(MEM_stage_inst_dmem_n16863), .ZN(MEM_stage_inst_dmem_n16854) );
NAND2_X1 MEM_stage_inst_dmem_U14796 ( .A1(MEM_stage_inst_dmem_n16852), .A2(MEM_stage_inst_dmem_n16851), .ZN(MEM_stage_inst_dmem_n10913) );
NAND2_X1 MEM_stage_inst_dmem_U14795 ( .A1(EX_pipeline_reg_out_11), .A2(MEM_stage_inst_dmem_n16864), .ZN(MEM_stage_inst_dmem_n16851) );
NAND2_X1 MEM_stage_inst_dmem_U14794 ( .A1(MEM_stage_inst_dmem_ram_1638), .A2(MEM_stage_inst_dmem_n16863), .ZN(MEM_stage_inst_dmem_n16852) );
NAND2_X1 MEM_stage_inst_dmem_U14793 ( .A1(MEM_stage_inst_dmem_n16850), .A2(MEM_stage_inst_dmem_n16849), .ZN(MEM_stage_inst_dmem_n10914) );
NAND2_X1 MEM_stage_inst_dmem_U14792 ( .A1(EX_pipeline_reg_out_12), .A2(MEM_stage_inst_dmem_n16864), .ZN(MEM_stage_inst_dmem_n16849) );
NAND2_X1 MEM_stage_inst_dmem_U14791 ( .A1(MEM_stage_inst_dmem_ram_1639), .A2(MEM_stage_inst_dmem_n16863), .ZN(MEM_stage_inst_dmem_n16850) );
NAND2_X1 MEM_stage_inst_dmem_U14790 ( .A1(MEM_stage_inst_dmem_n16848), .A2(MEM_stage_inst_dmem_n16847), .ZN(MEM_stage_inst_dmem_n10915) );
NAND2_X1 MEM_stage_inst_dmem_U14789 ( .A1(EX_pipeline_reg_out_13), .A2(MEM_stage_inst_dmem_n16864), .ZN(MEM_stage_inst_dmem_n16847) );
NAND2_X1 MEM_stage_inst_dmem_U14788 ( .A1(MEM_stage_inst_dmem_ram_1640), .A2(MEM_stage_inst_dmem_n16863), .ZN(MEM_stage_inst_dmem_n16848) );
NAND2_X1 MEM_stage_inst_dmem_U14787 ( .A1(MEM_stage_inst_dmem_n16846), .A2(MEM_stage_inst_dmem_n16845), .ZN(MEM_stage_inst_dmem_n10916) );
NAND2_X1 MEM_stage_inst_dmem_U14786 ( .A1(EX_pipeline_reg_out_14), .A2(MEM_stage_inst_dmem_n16864), .ZN(MEM_stage_inst_dmem_n16845) );
NAND2_X1 MEM_stage_inst_dmem_U14785 ( .A1(MEM_stage_inst_dmem_ram_1641), .A2(MEM_stage_inst_dmem_n16863), .ZN(MEM_stage_inst_dmem_n16846) );
NAND2_X1 MEM_stage_inst_dmem_U14784 ( .A1(MEM_stage_inst_dmem_n16844), .A2(MEM_stage_inst_dmem_n16843), .ZN(MEM_stage_inst_dmem_n10917) );
NAND2_X1 MEM_stage_inst_dmem_U14783 ( .A1(EX_pipeline_reg_out_15), .A2(MEM_stage_inst_dmem_n16864), .ZN(MEM_stage_inst_dmem_n16843) );
NAND2_X1 MEM_stage_inst_dmem_U14782 ( .A1(MEM_stage_inst_dmem_ram_1642), .A2(MEM_stage_inst_dmem_n16863), .ZN(MEM_stage_inst_dmem_n16844) );
NAND2_X1 MEM_stage_inst_dmem_U14781 ( .A1(MEM_stage_inst_dmem_n16842), .A2(MEM_stage_inst_dmem_n16841), .ZN(MEM_stage_inst_dmem_n10918) );
NAND2_X1 MEM_stage_inst_dmem_U14780 ( .A1(EX_pipeline_reg_out_16), .A2(MEM_stage_inst_dmem_n16864), .ZN(MEM_stage_inst_dmem_n16841) );
NAND2_X1 MEM_stage_inst_dmem_U14779 ( .A1(MEM_stage_inst_dmem_ram_1643), .A2(MEM_stage_inst_dmem_n16863), .ZN(MEM_stage_inst_dmem_n16842) );
NAND2_X1 MEM_stage_inst_dmem_U14778 ( .A1(MEM_stage_inst_dmem_n16840), .A2(MEM_stage_inst_dmem_n16839), .ZN(MEM_stage_inst_dmem_n10919) );
NAND2_X1 MEM_stage_inst_dmem_U14777 ( .A1(EX_pipeline_reg_out_17), .A2(MEM_stage_inst_dmem_n16864), .ZN(MEM_stage_inst_dmem_n16839) );
NAND2_X1 MEM_stage_inst_dmem_U14776 ( .A1(MEM_stage_inst_dmem_ram_1644), .A2(MEM_stage_inst_dmem_n16863), .ZN(MEM_stage_inst_dmem_n16840) );
NAND2_X1 MEM_stage_inst_dmem_U14775 ( .A1(MEM_stage_inst_dmem_n16838), .A2(MEM_stage_inst_dmem_n16837), .ZN(MEM_stage_inst_dmem_n10920) );
NAND2_X1 MEM_stage_inst_dmem_U14774 ( .A1(EX_pipeline_reg_out_18), .A2(MEM_stage_inst_dmem_n16864), .ZN(MEM_stage_inst_dmem_n16837) );
NAND2_X1 MEM_stage_inst_dmem_U14773 ( .A1(MEM_stage_inst_dmem_ram_1645), .A2(MEM_stage_inst_dmem_n16863), .ZN(MEM_stage_inst_dmem_n16838) );
NAND2_X1 MEM_stage_inst_dmem_U14772 ( .A1(MEM_stage_inst_dmem_n16836), .A2(MEM_stage_inst_dmem_n16835), .ZN(MEM_stage_inst_dmem_n10921) );
NAND2_X1 MEM_stage_inst_dmem_U14771 ( .A1(EX_pipeline_reg_out_19), .A2(MEM_stage_inst_dmem_n16864), .ZN(MEM_stage_inst_dmem_n16835) );
NAND2_X1 MEM_stage_inst_dmem_U14770 ( .A1(MEM_stage_inst_dmem_ram_1646), .A2(MEM_stage_inst_dmem_n16863), .ZN(MEM_stage_inst_dmem_n16836) );
NAND2_X1 MEM_stage_inst_dmem_U14769 ( .A1(MEM_stage_inst_dmem_n16834), .A2(MEM_stage_inst_dmem_n16833), .ZN(MEM_stage_inst_dmem_n10922) );
NAND2_X1 MEM_stage_inst_dmem_U14768 ( .A1(EX_pipeline_reg_out_20), .A2(MEM_stage_inst_dmem_n16864), .ZN(MEM_stage_inst_dmem_n16833) );
NAND2_X1 MEM_stage_inst_dmem_U14767 ( .A1(MEM_stage_inst_dmem_ram_1647), .A2(MEM_stage_inst_dmem_n16863), .ZN(MEM_stage_inst_dmem_n16834) );
NAND2_X1 MEM_stage_inst_dmem_U14766 ( .A1(MEM_stage_inst_dmem_n21249), .A2(MEM_stage_inst_dmem_n17037), .ZN(MEM_stage_inst_dmem_n16863) );
NAND2_X1 MEM_stage_inst_dmem_U14765 ( .A1(MEM_stage_inst_dmem_n16832), .A2(MEM_stage_inst_dmem_n16831), .ZN(MEM_stage_inst_dmem_n10923) );
NAND2_X1 MEM_stage_inst_dmem_U14764 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n16830), .ZN(MEM_stage_inst_dmem_n16831) );
NAND2_X1 MEM_stage_inst_dmem_U14763 ( .A1(MEM_stage_inst_dmem_ram_1648), .A2(MEM_stage_inst_dmem_n16829), .ZN(MEM_stage_inst_dmem_n16832) );
NAND2_X1 MEM_stage_inst_dmem_U14762 ( .A1(MEM_stage_inst_dmem_n16828), .A2(MEM_stage_inst_dmem_n16827), .ZN(MEM_stage_inst_dmem_n10924) );
NAND2_X1 MEM_stage_inst_dmem_U14761 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n16830), .ZN(MEM_stage_inst_dmem_n16827) );
NAND2_X1 MEM_stage_inst_dmem_U14760 ( .A1(MEM_stage_inst_dmem_ram_1649), .A2(MEM_stage_inst_dmem_n16829), .ZN(MEM_stage_inst_dmem_n16828) );
NAND2_X1 MEM_stage_inst_dmem_U14759 ( .A1(MEM_stage_inst_dmem_n16826), .A2(MEM_stage_inst_dmem_n16825), .ZN(MEM_stage_inst_dmem_n10925) );
NAND2_X1 MEM_stage_inst_dmem_U14758 ( .A1(MEM_stage_inst_dmem_n18027), .A2(MEM_stage_inst_dmem_n16830), .ZN(MEM_stage_inst_dmem_n16825) );
BUF_X1 MEM_stage_inst_dmem_U14757 ( .A(EX_pipeline_reg_out_7), .Z(MEM_stage_inst_dmem_n18027) );
NAND2_X1 MEM_stage_inst_dmem_U14756 ( .A1(MEM_stage_inst_dmem_ram_1650), .A2(MEM_stage_inst_dmem_n16829), .ZN(MEM_stage_inst_dmem_n16826) );
NAND2_X1 MEM_stage_inst_dmem_U14755 ( .A1(MEM_stage_inst_dmem_n16824), .A2(MEM_stage_inst_dmem_n16823), .ZN(MEM_stage_inst_dmem_n10926) );
NAND2_X1 MEM_stage_inst_dmem_U14754 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n16830), .ZN(MEM_stage_inst_dmem_n16823) );
NAND2_X1 MEM_stage_inst_dmem_U14753 ( .A1(MEM_stage_inst_dmem_ram_1651), .A2(MEM_stage_inst_dmem_n16829), .ZN(MEM_stage_inst_dmem_n16824) );
NAND2_X1 MEM_stage_inst_dmem_U14752 ( .A1(MEM_stage_inst_dmem_n16822), .A2(MEM_stage_inst_dmem_n16821), .ZN(MEM_stage_inst_dmem_n10927) );
NAND2_X1 MEM_stage_inst_dmem_U14751 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n16830), .ZN(MEM_stage_inst_dmem_n16821) );
NAND2_X1 MEM_stage_inst_dmem_U14750 ( .A1(MEM_stage_inst_dmem_ram_1652), .A2(MEM_stage_inst_dmem_n16829), .ZN(MEM_stage_inst_dmem_n16822) );
NAND2_X1 MEM_stage_inst_dmem_U14749 ( .A1(MEM_stage_inst_dmem_n16820), .A2(MEM_stage_inst_dmem_n16819), .ZN(MEM_stage_inst_dmem_n10928) );
NAND2_X1 MEM_stage_inst_dmem_U14748 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n16830), .ZN(MEM_stage_inst_dmem_n16819) );
NAND2_X1 MEM_stage_inst_dmem_U14747 ( .A1(MEM_stage_inst_dmem_ram_1653), .A2(MEM_stage_inst_dmem_n16829), .ZN(MEM_stage_inst_dmem_n16820) );
NAND2_X1 MEM_stage_inst_dmem_U14746 ( .A1(MEM_stage_inst_dmem_n16818), .A2(MEM_stage_inst_dmem_n16817), .ZN(MEM_stage_inst_dmem_n10929) );
NAND2_X1 MEM_stage_inst_dmem_U14745 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n16830), .ZN(MEM_stage_inst_dmem_n16817) );
NAND2_X1 MEM_stage_inst_dmem_U14744 ( .A1(MEM_stage_inst_dmem_ram_1654), .A2(MEM_stage_inst_dmem_n16829), .ZN(MEM_stage_inst_dmem_n16818) );
NAND2_X1 MEM_stage_inst_dmem_U14743 ( .A1(MEM_stage_inst_dmem_n16816), .A2(MEM_stage_inst_dmem_n16815), .ZN(MEM_stage_inst_dmem_n10930) );
NAND2_X1 MEM_stage_inst_dmem_U14742 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n16830), .ZN(MEM_stage_inst_dmem_n16815) );
NAND2_X1 MEM_stage_inst_dmem_U14741 ( .A1(MEM_stage_inst_dmem_ram_1655), .A2(MEM_stage_inst_dmem_n16829), .ZN(MEM_stage_inst_dmem_n16816) );
NAND2_X1 MEM_stage_inst_dmem_U14740 ( .A1(MEM_stage_inst_dmem_n16814), .A2(MEM_stage_inst_dmem_n16813), .ZN(MEM_stage_inst_dmem_n10931) );
NAND2_X1 MEM_stage_inst_dmem_U14739 ( .A1(MEM_stage_inst_dmem_n18013), .A2(MEM_stage_inst_dmem_n16830), .ZN(MEM_stage_inst_dmem_n16813) );
BUF_X1 MEM_stage_inst_dmem_U14738 ( .A(EX_pipeline_reg_out_13), .Z(MEM_stage_inst_dmem_n18013) );
NAND2_X1 MEM_stage_inst_dmem_U14737 ( .A1(MEM_stage_inst_dmem_ram_1656), .A2(MEM_stage_inst_dmem_n16829), .ZN(MEM_stage_inst_dmem_n16814) );
NAND2_X1 MEM_stage_inst_dmem_U14736 ( .A1(MEM_stage_inst_dmem_n16812), .A2(MEM_stage_inst_dmem_n16811), .ZN(MEM_stage_inst_dmem_n10932) );
NAND2_X1 MEM_stage_inst_dmem_U14735 ( .A1(EX_pipeline_reg_out_14), .A2(MEM_stage_inst_dmem_n16830), .ZN(MEM_stage_inst_dmem_n16811) );
NAND2_X1 MEM_stage_inst_dmem_U14733 ( .A1(MEM_stage_inst_dmem_ram_1657), .A2(MEM_stage_inst_dmem_n16829), .ZN(MEM_stage_inst_dmem_n16812) );
NAND2_X1 MEM_stage_inst_dmem_U14732 ( .A1(MEM_stage_inst_dmem_n16810), .A2(MEM_stage_inst_dmem_n16809), .ZN(MEM_stage_inst_dmem_n10933) );
NAND2_X1 MEM_stage_inst_dmem_U14731 ( .A1(MEM_stage_inst_dmem_n18007), .A2(MEM_stage_inst_dmem_n16830), .ZN(MEM_stage_inst_dmem_n16809) );
BUF_X1 MEM_stage_inst_dmem_U14730 ( .A(EX_pipeline_reg_out_15), .Z(MEM_stage_inst_dmem_n18007) );
NAND2_X1 MEM_stage_inst_dmem_U14729 ( .A1(MEM_stage_inst_dmem_ram_1658), .A2(MEM_stage_inst_dmem_n16829), .ZN(MEM_stage_inst_dmem_n16810) );
NAND2_X1 MEM_stage_inst_dmem_U14728 ( .A1(MEM_stage_inst_dmem_n16808), .A2(MEM_stage_inst_dmem_n16807), .ZN(MEM_stage_inst_dmem_n10934) );
NAND2_X1 MEM_stage_inst_dmem_U14727 ( .A1(MEM_stage_inst_dmem_n18004), .A2(MEM_stage_inst_dmem_n16830), .ZN(MEM_stage_inst_dmem_n16807) );
BUF_X1 MEM_stage_inst_dmem_U14726 ( .A(EX_pipeline_reg_out_16), .Z(MEM_stage_inst_dmem_n18004) );
NAND2_X1 MEM_stage_inst_dmem_U14725 ( .A1(MEM_stage_inst_dmem_ram_1659), .A2(MEM_stage_inst_dmem_n16829), .ZN(MEM_stage_inst_dmem_n16808) );
NAND2_X1 MEM_stage_inst_dmem_U14724 ( .A1(MEM_stage_inst_dmem_n16806), .A2(MEM_stage_inst_dmem_n16805), .ZN(MEM_stage_inst_dmem_n10935) );
NAND2_X1 MEM_stage_inst_dmem_U14723 ( .A1(MEM_stage_inst_dmem_n18001), .A2(MEM_stage_inst_dmem_n16830), .ZN(MEM_stage_inst_dmem_n16805) );
BUF_X1 MEM_stage_inst_dmem_U14722 ( .A(EX_pipeline_reg_out_17), .Z(MEM_stage_inst_dmem_n18001) );
NAND2_X1 MEM_stage_inst_dmem_U14721 ( .A1(MEM_stage_inst_dmem_ram_1660), .A2(MEM_stage_inst_dmem_n16829), .ZN(MEM_stage_inst_dmem_n16806) );
NAND2_X1 MEM_stage_inst_dmem_U14720 ( .A1(MEM_stage_inst_dmem_n16804), .A2(MEM_stage_inst_dmem_n16803), .ZN(MEM_stage_inst_dmem_n10936) );
NAND2_X1 MEM_stage_inst_dmem_U14719 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n16830), .ZN(MEM_stage_inst_dmem_n16803) );
NAND2_X1 MEM_stage_inst_dmem_U14718 ( .A1(MEM_stage_inst_dmem_ram_1661), .A2(MEM_stage_inst_dmem_n16829), .ZN(MEM_stage_inst_dmem_n16804) );
NAND2_X1 MEM_stage_inst_dmem_U14717 ( .A1(MEM_stage_inst_dmem_n16802), .A2(MEM_stage_inst_dmem_n16801), .ZN(MEM_stage_inst_dmem_n10937) );
NAND2_X1 MEM_stage_inst_dmem_U14716 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n16830), .ZN(MEM_stage_inst_dmem_n16801) );
NAND2_X1 MEM_stage_inst_dmem_U14715 ( .A1(MEM_stage_inst_dmem_ram_1662), .A2(MEM_stage_inst_dmem_n16829), .ZN(MEM_stage_inst_dmem_n16802) );
NAND2_X1 MEM_stage_inst_dmem_U14714 ( .A1(MEM_stage_inst_dmem_n16800), .A2(MEM_stage_inst_dmem_n16799), .ZN(MEM_stage_inst_dmem_n10938) );
NAND2_X1 MEM_stage_inst_dmem_U14713 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n16830), .ZN(MEM_stage_inst_dmem_n16799) );
NAND2_X1 MEM_stage_inst_dmem_U14712 ( .A1(MEM_stage_inst_dmem_ram_1663), .A2(MEM_stage_inst_dmem_n16829), .ZN(MEM_stage_inst_dmem_n16800) );
NAND2_X1 MEM_stage_inst_dmem_U14711 ( .A1(MEM_stage_inst_dmem_n21214), .A2(MEM_stage_inst_dmem_n17037), .ZN(MEM_stage_inst_dmem_n16829) );
NAND2_X1 MEM_stage_inst_dmem_U14710 ( .A1(MEM_stage_inst_dmem_n16798), .A2(MEM_stage_inst_dmem_n16797), .ZN(MEM_stage_inst_dmem_n10939) );
NAND2_X1 MEM_stage_inst_dmem_U14709 ( .A1(MEM_stage_inst_dmem_n19275), .A2(MEM_stage_inst_dmem_n16796), .ZN(MEM_stage_inst_dmem_n16797) );
NAND2_X1 MEM_stage_inst_dmem_U14708 ( .A1(MEM_stage_inst_dmem_ram_1664), .A2(MEM_stage_inst_dmem_n16795), .ZN(MEM_stage_inst_dmem_n16798) );
NAND2_X1 MEM_stage_inst_dmem_U14707 ( .A1(MEM_stage_inst_dmem_n16794), .A2(MEM_stage_inst_dmem_n16793), .ZN(MEM_stage_inst_dmem_n10940) );
NAND2_X1 MEM_stage_inst_dmem_U14706 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n16796), .ZN(MEM_stage_inst_dmem_n16793) );
NAND2_X1 MEM_stage_inst_dmem_U14705 ( .A1(MEM_stage_inst_dmem_ram_1665), .A2(MEM_stage_inst_dmem_n16795), .ZN(MEM_stage_inst_dmem_n16794) );
NAND2_X1 MEM_stage_inst_dmem_U14704 ( .A1(MEM_stage_inst_dmem_n16791), .A2(MEM_stage_inst_dmem_n16790), .ZN(MEM_stage_inst_dmem_n10941) );
NAND2_X1 MEM_stage_inst_dmem_U14703 ( .A1(MEM_stage_inst_dmem_n16789), .A2(MEM_stage_inst_dmem_n16796), .ZN(MEM_stage_inst_dmem_n16790) );
NAND2_X1 MEM_stage_inst_dmem_U14702 ( .A1(MEM_stage_inst_dmem_ram_1666), .A2(MEM_stage_inst_dmem_n16795), .ZN(MEM_stage_inst_dmem_n16791) );
NAND2_X1 MEM_stage_inst_dmem_U14701 ( .A1(MEM_stage_inst_dmem_n16788), .A2(MEM_stage_inst_dmem_n16787), .ZN(MEM_stage_inst_dmem_n10942) );
NAND2_X1 MEM_stage_inst_dmem_U14700 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n16796), .ZN(MEM_stage_inst_dmem_n16787) );
NAND2_X1 MEM_stage_inst_dmem_U14699 ( .A1(MEM_stage_inst_dmem_ram_1667), .A2(MEM_stage_inst_dmem_n16795), .ZN(MEM_stage_inst_dmem_n16788) );
NAND2_X1 MEM_stage_inst_dmem_U14698 ( .A1(MEM_stage_inst_dmem_n16786), .A2(MEM_stage_inst_dmem_n16785), .ZN(MEM_stage_inst_dmem_n10943) );
NAND2_X1 MEM_stage_inst_dmem_U14697 ( .A1(MEM_stage_inst_dmem_n16784), .A2(MEM_stage_inst_dmem_n16796), .ZN(MEM_stage_inst_dmem_n16785) );
NAND2_X1 MEM_stage_inst_dmem_U14696 ( .A1(MEM_stage_inst_dmem_ram_1668), .A2(MEM_stage_inst_dmem_n16795), .ZN(MEM_stage_inst_dmem_n16786) );
NAND2_X1 MEM_stage_inst_dmem_U14695 ( .A1(MEM_stage_inst_dmem_n16783), .A2(MEM_stage_inst_dmem_n16782), .ZN(MEM_stage_inst_dmem_n10944) );
NAND2_X1 MEM_stage_inst_dmem_U14694 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n16796), .ZN(MEM_stage_inst_dmem_n16782) );
NAND2_X1 MEM_stage_inst_dmem_U14693 ( .A1(MEM_stage_inst_dmem_ram_1669), .A2(MEM_stage_inst_dmem_n16795), .ZN(MEM_stage_inst_dmem_n16783) );
NAND2_X1 MEM_stage_inst_dmem_U14692 ( .A1(MEM_stage_inst_dmem_n16781), .A2(MEM_stage_inst_dmem_n16780), .ZN(MEM_stage_inst_dmem_n10945) );
NAND2_X1 MEM_stage_inst_dmem_U14691 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n16796), .ZN(MEM_stage_inst_dmem_n16780) );
NAND2_X1 MEM_stage_inst_dmem_U14690 ( .A1(MEM_stage_inst_dmem_ram_1670), .A2(MEM_stage_inst_dmem_n16795), .ZN(MEM_stage_inst_dmem_n16781) );
NAND2_X1 MEM_stage_inst_dmem_U14689 ( .A1(MEM_stage_inst_dmem_n16779), .A2(MEM_stage_inst_dmem_n16778), .ZN(MEM_stage_inst_dmem_n10946) );
NAND2_X1 MEM_stage_inst_dmem_U14688 ( .A1(MEM_stage_inst_dmem_n16777), .A2(MEM_stage_inst_dmem_n16796), .ZN(MEM_stage_inst_dmem_n16778) );
NAND2_X1 MEM_stage_inst_dmem_U14687 ( .A1(MEM_stage_inst_dmem_ram_1671), .A2(MEM_stage_inst_dmem_n16795), .ZN(MEM_stage_inst_dmem_n16779) );
NAND2_X1 MEM_stage_inst_dmem_U14686 ( .A1(MEM_stage_inst_dmem_n16776), .A2(MEM_stage_inst_dmem_n16775), .ZN(MEM_stage_inst_dmem_n10947) );
NAND2_X1 MEM_stage_inst_dmem_U14685 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n16796), .ZN(MEM_stage_inst_dmem_n16775) );
NAND2_X1 MEM_stage_inst_dmem_U14684 ( .A1(MEM_stage_inst_dmem_ram_1672), .A2(MEM_stage_inst_dmem_n16795), .ZN(MEM_stage_inst_dmem_n16776) );
NAND2_X1 MEM_stage_inst_dmem_U14683 ( .A1(MEM_stage_inst_dmem_n16774), .A2(MEM_stage_inst_dmem_n16773), .ZN(MEM_stage_inst_dmem_n10948) );
NAND2_X1 MEM_stage_inst_dmem_U14682 ( .A1(MEM_stage_inst_dmem_n16772), .A2(MEM_stage_inst_dmem_n16796), .ZN(MEM_stage_inst_dmem_n16773) );
NAND2_X1 MEM_stage_inst_dmem_U14681 ( .A1(MEM_stage_inst_dmem_ram_1673), .A2(MEM_stage_inst_dmem_n16795), .ZN(MEM_stage_inst_dmem_n16774) );
NAND2_X1 MEM_stage_inst_dmem_U14680 ( .A1(MEM_stage_inst_dmem_n16771), .A2(MEM_stage_inst_dmem_n16770), .ZN(MEM_stage_inst_dmem_n10949) );
NAND2_X1 MEM_stage_inst_dmem_U14679 ( .A1(MEM_stage_inst_dmem_n16769), .A2(MEM_stage_inst_dmem_n16796), .ZN(MEM_stage_inst_dmem_n16770) );
NAND2_X1 MEM_stage_inst_dmem_U14678 ( .A1(MEM_stage_inst_dmem_ram_1674), .A2(MEM_stage_inst_dmem_n16795), .ZN(MEM_stage_inst_dmem_n16771) );
NAND2_X1 MEM_stage_inst_dmem_U14677 ( .A1(MEM_stage_inst_dmem_n16768), .A2(MEM_stage_inst_dmem_n16767), .ZN(MEM_stage_inst_dmem_n10950) );
NAND2_X1 MEM_stage_inst_dmem_U14676 ( .A1(MEM_stage_inst_dmem_n14705), .A2(MEM_stage_inst_dmem_n16796), .ZN(MEM_stage_inst_dmem_n16767) );
NAND2_X1 MEM_stage_inst_dmem_U14675 ( .A1(MEM_stage_inst_dmem_ram_1675), .A2(MEM_stage_inst_dmem_n16795), .ZN(MEM_stage_inst_dmem_n16768) );
NAND2_X1 MEM_stage_inst_dmem_U14674 ( .A1(MEM_stage_inst_dmem_n16766), .A2(MEM_stage_inst_dmem_n16765), .ZN(MEM_stage_inst_dmem_n10951) );
NAND2_X1 MEM_stage_inst_dmem_U14673 ( .A1(MEM_stage_inst_dmem_n14702), .A2(MEM_stage_inst_dmem_n16796), .ZN(MEM_stage_inst_dmem_n16765) );
NAND2_X1 MEM_stage_inst_dmem_U14672 ( .A1(MEM_stage_inst_dmem_ram_1676), .A2(MEM_stage_inst_dmem_n16795), .ZN(MEM_stage_inst_dmem_n16766) );
NAND2_X1 MEM_stage_inst_dmem_U14671 ( .A1(MEM_stage_inst_dmem_n16764), .A2(MEM_stage_inst_dmem_n16763), .ZN(MEM_stage_inst_dmem_n10952) );
NAND2_X1 MEM_stage_inst_dmem_U14670 ( .A1(MEM_stage_inst_dmem_n19242), .A2(MEM_stage_inst_dmem_n16796), .ZN(MEM_stage_inst_dmem_n16763) );
NAND2_X1 MEM_stage_inst_dmem_U14669 ( .A1(MEM_stage_inst_dmem_ram_1677), .A2(MEM_stage_inst_dmem_n16795), .ZN(MEM_stage_inst_dmem_n16764) );
NAND2_X1 MEM_stage_inst_dmem_U14668 ( .A1(MEM_stage_inst_dmem_n16762), .A2(MEM_stage_inst_dmem_n16761), .ZN(MEM_stage_inst_dmem_n10953) );
NAND2_X1 MEM_stage_inst_dmem_U14667 ( .A1(MEM_stage_inst_dmem_n115), .A2(MEM_stage_inst_dmem_n16796), .ZN(MEM_stage_inst_dmem_n16761) );
NAND2_X1 MEM_stage_inst_dmem_U14666 ( .A1(MEM_stage_inst_dmem_ram_1678), .A2(MEM_stage_inst_dmem_n16795), .ZN(MEM_stage_inst_dmem_n16762) );
NAND2_X1 MEM_stage_inst_dmem_U14665 ( .A1(MEM_stage_inst_dmem_n16760), .A2(MEM_stage_inst_dmem_n16759), .ZN(MEM_stage_inst_dmem_n10954) );
NAND2_X1 MEM_stage_inst_dmem_U14664 ( .A1(MEM_stage_inst_dmem_n16758), .A2(MEM_stage_inst_dmem_n16796), .ZN(MEM_stage_inst_dmem_n16759) );
INV_X1 MEM_stage_inst_dmem_U14663 ( .A(MEM_stage_inst_dmem_n16795), .ZN(MEM_stage_inst_dmem_n16796) );
NAND2_X1 MEM_stage_inst_dmem_U14662 ( .A1(MEM_stage_inst_dmem_ram_1679), .A2(MEM_stage_inst_dmem_n16795), .ZN(MEM_stage_inst_dmem_n16760) );
NAND2_X1 MEM_stage_inst_dmem_U14661 ( .A1(MEM_stage_inst_dmem_n21179), .A2(MEM_stage_inst_dmem_n17037), .ZN(MEM_stage_inst_dmem_n16795) );
NAND2_X1 MEM_stage_inst_dmem_U14660 ( .A1(MEM_stage_inst_dmem_n16757), .A2(MEM_stage_inst_dmem_n16756), .ZN(MEM_stage_inst_dmem_n10955) );
NAND2_X1 MEM_stage_inst_dmem_U14659 ( .A1(MEM_stage_inst_dmem_n20551), .A2(MEM_stage_inst_dmem_n16755), .ZN(MEM_stage_inst_dmem_n16756) );
NAND2_X1 MEM_stage_inst_dmem_U14658 ( .A1(MEM_stage_inst_dmem_ram_1680), .A2(MEM_stage_inst_dmem_n16754), .ZN(MEM_stage_inst_dmem_n16757) );
NAND2_X1 MEM_stage_inst_dmem_U14657 ( .A1(MEM_stage_inst_dmem_n16753), .A2(MEM_stage_inst_dmem_n16752), .ZN(MEM_stage_inst_dmem_n10956) );
NAND2_X1 MEM_stage_inst_dmem_U14656 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n16755), .ZN(MEM_stage_inst_dmem_n16752) );
NAND2_X1 MEM_stage_inst_dmem_U14655 ( .A1(MEM_stage_inst_dmem_ram_1681), .A2(MEM_stage_inst_dmem_n16754), .ZN(MEM_stage_inst_dmem_n16753) );
NAND2_X1 MEM_stage_inst_dmem_U14654 ( .A1(MEM_stage_inst_dmem_n16751), .A2(MEM_stage_inst_dmem_n16750), .ZN(MEM_stage_inst_dmem_n10957) );
NAND2_X1 MEM_stage_inst_dmem_U14653 ( .A1(MEM_stage_inst_dmem_n16789), .A2(MEM_stage_inst_dmem_n16755), .ZN(MEM_stage_inst_dmem_n16750) );
NAND2_X1 MEM_stage_inst_dmem_U14652 ( .A1(MEM_stage_inst_dmem_ram_1682), .A2(MEM_stage_inst_dmem_n16754), .ZN(MEM_stage_inst_dmem_n16751) );
NAND2_X1 MEM_stage_inst_dmem_U14651 ( .A1(MEM_stage_inst_dmem_n16749), .A2(MEM_stage_inst_dmem_n16748), .ZN(MEM_stage_inst_dmem_n10958) );
NAND2_X1 MEM_stage_inst_dmem_U14650 ( .A1(MEM_stage_inst_dmem_n13064), .A2(MEM_stage_inst_dmem_n16755), .ZN(MEM_stage_inst_dmem_n16748) );
NAND2_X1 MEM_stage_inst_dmem_U14649 ( .A1(MEM_stage_inst_dmem_ram_1683), .A2(MEM_stage_inst_dmem_n16754), .ZN(MEM_stage_inst_dmem_n16749) );
NAND2_X1 MEM_stage_inst_dmem_U14648 ( .A1(MEM_stage_inst_dmem_n16747), .A2(MEM_stage_inst_dmem_n16746), .ZN(MEM_stage_inst_dmem_n10959) );
NAND2_X1 MEM_stage_inst_dmem_U14647 ( .A1(MEM_stage_inst_dmem_n16784), .A2(MEM_stage_inst_dmem_n16755), .ZN(MEM_stage_inst_dmem_n16746) );
NAND2_X1 MEM_stage_inst_dmem_U14646 ( .A1(MEM_stage_inst_dmem_ram_1684), .A2(MEM_stage_inst_dmem_n16754), .ZN(MEM_stage_inst_dmem_n16747) );
NAND2_X1 MEM_stage_inst_dmem_U14645 ( .A1(MEM_stage_inst_dmem_n16745), .A2(MEM_stage_inst_dmem_n16744), .ZN(MEM_stage_inst_dmem_n10960) );
NAND2_X1 MEM_stage_inst_dmem_U14644 ( .A1(MEM_stage_inst_dmem_n13059), .A2(MEM_stage_inst_dmem_n16755), .ZN(MEM_stage_inst_dmem_n16744) );
NAND2_X1 MEM_stage_inst_dmem_U14643 ( .A1(MEM_stage_inst_dmem_ram_1685), .A2(MEM_stage_inst_dmem_n16754), .ZN(MEM_stage_inst_dmem_n16745) );
NAND2_X1 MEM_stage_inst_dmem_U14642 ( .A1(MEM_stage_inst_dmem_n16743), .A2(MEM_stage_inst_dmem_n16742), .ZN(MEM_stage_inst_dmem_n10961) );
NAND2_X1 MEM_stage_inst_dmem_U14641 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n16755), .ZN(MEM_stage_inst_dmem_n16742) );
NAND2_X1 MEM_stage_inst_dmem_U14640 ( .A1(MEM_stage_inst_dmem_ram_1686), .A2(MEM_stage_inst_dmem_n16754), .ZN(MEM_stage_inst_dmem_n16743) );
NAND2_X1 MEM_stage_inst_dmem_U14639 ( .A1(MEM_stage_inst_dmem_n16741), .A2(MEM_stage_inst_dmem_n16740), .ZN(MEM_stage_inst_dmem_n10962) );
NAND2_X1 MEM_stage_inst_dmem_U14638 ( .A1(MEM_stage_inst_dmem_n16777), .A2(MEM_stage_inst_dmem_n16755), .ZN(MEM_stage_inst_dmem_n16740) );
NAND2_X1 MEM_stage_inst_dmem_U14637 ( .A1(MEM_stage_inst_dmem_ram_1687), .A2(MEM_stage_inst_dmem_n16754), .ZN(MEM_stage_inst_dmem_n16741) );
NAND2_X1 MEM_stage_inst_dmem_U14636 ( .A1(MEM_stage_inst_dmem_n16739), .A2(MEM_stage_inst_dmem_n16738), .ZN(MEM_stage_inst_dmem_n10963) );
NAND2_X1 MEM_stage_inst_dmem_U14635 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n16755), .ZN(MEM_stage_inst_dmem_n16738) );
NAND2_X1 MEM_stage_inst_dmem_U14634 ( .A1(MEM_stage_inst_dmem_ram_1688), .A2(MEM_stage_inst_dmem_n16754), .ZN(MEM_stage_inst_dmem_n16739) );
NAND2_X1 MEM_stage_inst_dmem_U14633 ( .A1(MEM_stage_inst_dmem_n16737), .A2(MEM_stage_inst_dmem_n16736), .ZN(MEM_stage_inst_dmem_n10964) );
NAND2_X1 MEM_stage_inst_dmem_U14632 ( .A1(MEM_stage_inst_dmem_n16772), .A2(MEM_stage_inst_dmem_n16755), .ZN(MEM_stage_inst_dmem_n16736) );
NAND2_X1 MEM_stage_inst_dmem_U14631 ( .A1(MEM_stage_inst_dmem_ram_1689), .A2(MEM_stage_inst_dmem_n16754), .ZN(MEM_stage_inst_dmem_n16737) );
NAND2_X1 MEM_stage_inst_dmem_U14630 ( .A1(MEM_stage_inst_dmem_n16735), .A2(MEM_stage_inst_dmem_n16734), .ZN(MEM_stage_inst_dmem_n10965) );
NAND2_X1 MEM_stage_inst_dmem_U14629 ( .A1(MEM_stage_inst_dmem_n16769), .A2(MEM_stage_inst_dmem_n16755), .ZN(MEM_stage_inst_dmem_n16734) );
NAND2_X1 MEM_stage_inst_dmem_U14628 ( .A1(MEM_stage_inst_dmem_ram_1690), .A2(MEM_stage_inst_dmem_n16754), .ZN(MEM_stage_inst_dmem_n16735) );
NAND2_X1 MEM_stage_inst_dmem_U14627 ( .A1(MEM_stage_inst_dmem_n16733), .A2(MEM_stage_inst_dmem_n16732), .ZN(MEM_stage_inst_dmem_n10966) );
NAND2_X1 MEM_stage_inst_dmem_U14626 ( .A1(MEM_stage_inst_dmem_n20518), .A2(MEM_stage_inst_dmem_n16755), .ZN(MEM_stage_inst_dmem_n16732) );
NAND2_X1 MEM_stage_inst_dmem_U14625 ( .A1(MEM_stage_inst_dmem_ram_1691), .A2(MEM_stage_inst_dmem_n16754), .ZN(MEM_stage_inst_dmem_n16733) );
NAND2_X1 MEM_stage_inst_dmem_U14624 ( .A1(MEM_stage_inst_dmem_n16731), .A2(MEM_stage_inst_dmem_n16730), .ZN(MEM_stage_inst_dmem_n10967) );
NAND2_X1 MEM_stage_inst_dmem_U14623 ( .A1(MEM_stage_inst_dmem_n20515), .A2(MEM_stage_inst_dmem_n16755), .ZN(MEM_stage_inst_dmem_n16730) );
NAND2_X1 MEM_stage_inst_dmem_U14622 ( .A1(MEM_stage_inst_dmem_ram_1692), .A2(MEM_stage_inst_dmem_n16754), .ZN(MEM_stage_inst_dmem_n16731) );
NAND2_X1 MEM_stage_inst_dmem_U14621 ( .A1(MEM_stage_inst_dmem_n16729), .A2(MEM_stage_inst_dmem_n16728), .ZN(MEM_stage_inst_dmem_n10968) );
NAND2_X1 MEM_stage_inst_dmem_U14620 ( .A1(MEM_stage_inst_dmem_n20512), .A2(MEM_stage_inst_dmem_n16755), .ZN(MEM_stage_inst_dmem_n16728) );
NAND2_X1 MEM_stage_inst_dmem_U14619 ( .A1(MEM_stage_inst_dmem_ram_1693), .A2(MEM_stage_inst_dmem_n16754), .ZN(MEM_stage_inst_dmem_n16729) );
NAND2_X1 MEM_stage_inst_dmem_U14618 ( .A1(MEM_stage_inst_dmem_n16727), .A2(MEM_stage_inst_dmem_n16726), .ZN(MEM_stage_inst_dmem_n10969) );
NAND2_X1 MEM_stage_inst_dmem_U14617 ( .A1(MEM_stage_inst_dmem_n20509), .A2(MEM_stage_inst_dmem_n16755), .ZN(MEM_stage_inst_dmem_n16726) );
NAND2_X1 MEM_stage_inst_dmem_U14616 ( .A1(MEM_stage_inst_dmem_ram_1694), .A2(MEM_stage_inst_dmem_n16754), .ZN(MEM_stage_inst_dmem_n16727) );
NAND2_X1 MEM_stage_inst_dmem_U14615 ( .A1(MEM_stage_inst_dmem_n16725), .A2(MEM_stage_inst_dmem_n16724), .ZN(MEM_stage_inst_dmem_n10970) );
NAND2_X1 MEM_stage_inst_dmem_U14614 ( .A1(MEM_stage_inst_dmem_n16758), .A2(MEM_stage_inst_dmem_n16755), .ZN(MEM_stage_inst_dmem_n16724) );
INV_X1 MEM_stage_inst_dmem_U14613 ( .A(MEM_stage_inst_dmem_n16754), .ZN(MEM_stage_inst_dmem_n16755) );
NAND2_X1 MEM_stage_inst_dmem_U14612 ( .A1(MEM_stage_inst_dmem_ram_1695), .A2(MEM_stage_inst_dmem_n16754), .ZN(MEM_stage_inst_dmem_n16725) );
NAND2_X1 MEM_stage_inst_dmem_U14611 ( .A1(MEM_stage_inst_dmem_n21144), .A2(MEM_stage_inst_dmem_n17037), .ZN(MEM_stage_inst_dmem_n16754) );
NAND2_X1 MEM_stage_inst_dmem_U14610 ( .A1(MEM_stage_inst_dmem_n16723), .A2(MEM_stage_inst_dmem_n16722), .ZN(MEM_stage_inst_dmem_n10971) );
NAND2_X1 MEM_stage_inst_dmem_U14609 ( .A1(EX_pipeline_reg_out_5), .A2(MEM_stage_inst_dmem_n16721), .ZN(MEM_stage_inst_dmem_n16722) );
NAND2_X1 MEM_stage_inst_dmem_U14608 ( .A1(MEM_stage_inst_dmem_ram_1696), .A2(MEM_stage_inst_dmem_n16720), .ZN(MEM_stage_inst_dmem_n16723) );
NAND2_X1 MEM_stage_inst_dmem_U14607 ( .A1(MEM_stage_inst_dmem_n16719), .A2(MEM_stage_inst_dmem_n16718), .ZN(MEM_stage_inst_dmem_n10972) );
NAND2_X1 MEM_stage_inst_dmem_U14606 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n16721), .ZN(MEM_stage_inst_dmem_n16718) );
NAND2_X1 MEM_stage_inst_dmem_U14605 ( .A1(MEM_stage_inst_dmem_ram_1697), .A2(MEM_stage_inst_dmem_n16720), .ZN(MEM_stage_inst_dmem_n16719) );
NAND2_X1 MEM_stage_inst_dmem_U14604 ( .A1(MEM_stage_inst_dmem_n16717), .A2(MEM_stage_inst_dmem_n16716), .ZN(MEM_stage_inst_dmem_n10973) );
NAND2_X1 MEM_stage_inst_dmem_U14603 ( .A1(MEM_stage_inst_dmem_n16789), .A2(MEM_stage_inst_dmem_n16721), .ZN(MEM_stage_inst_dmem_n16716) );
NAND2_X1 MEM_stage_inst_dmem_U14602 ( .A1(MEM_stage_inst_dmem_ram_1698), .A2(MEM_stage_inst_dmem_n16720), .ZN(MEM_stage_inst_dmem_n16717) );
NAND2_X1 MEM_stage_inst_dmem_U14601 ( .A1(MEM_stage_inst_dmem_n16715), .A2(MEM_stage_inst_dmem_n16714), .ZN(MEM_stage_inst_dmem_n10974) );
NAND2_X1 MEM_stage_inst_dmem_U14600 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n16721), .ZN(MEM_stage_inst_dmem_n16714) );
NAND2_X1 MEM_stage_inst_dmem_U14599 ( .A1(MEM_stage_inst_dmem_ram_1699), .A2(MEM_stage_inst_dmem_n16720), .ZN(MEM_stage_inst_dmem_n16715) );
NAND2_X1 MEM_stage_inst_dmem_U14598 ( .A1(MEM_stage_inst_dmem_n16713), .A2(MEM_stage_inst_dmem_n16712), .ZN(MEM_stage_inst_dmem_n10975) );
NAND2_X1 MEM_stage_inst_dmem_U14597 ( .A1(MEM_stage_inst_dmem_n16784), .A2(MEM_stage_inst_dmem_n16721), .ZN(MEM_stage_inst_dmem_n16712) );
NAND2_X1 MEM_stage_inst_dmem_U14596 ( .A1(MEM_stage_inst_dmem_ram_1700), .A2(MEM_stage_inst_dmem_n16720), .ZN(MEM_stage_inst_dmem_n16713) );
NAND2_X1 MEM_stage_inst_dmem_U14595 ( .A1(MEM_stage_inst_dmem_n16711), .A2(MEM_stage_inst_dmem_n16710), .ZN(MEM_stage_inst_dmem_n10976) );
NAND2_X1 MEM_stage_inst_dmem_U14594 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n16721), .ZN(MEM_stage_inst_dmem_n16710) );
NAND2_X1 MEM_stage_inst_dmem_U14593 ( .A1(MEM_stage_inst_dmem_ram_1701), .A2(MEM_stage_inst_dmem_n16720), .ZN(MEM_stage_inst_dmem_n16711) );
NAND2_X1 MEM_stage_inst_dmem_U14592 ( .A1(MEM_stage_inst_dmem_n16709), .A2(MEM_stage_inst_dmem_n16708), .ZN(MEM_stage_inst_dmem_n10977) );
NAND2_X1 MEM_stage_inst_dmem_U14591 ( .A1(MEM_stage_inst_dmem_n13056), .A2(MEM_stage_inst_dmem_n16721), .ZN(MEM_stage_inst_dmem_n16708) );
NAND2_X1 MEM_stage_inst_dmem_U14590 ( .A1(MEM_stage_inst_dmem_ram_1702), .A2(MEM_stage_inst_dmem_n16720), .ZN(MEM_stage_inst_dmem_n16709) );
NAND2_X1 MEM_stage_inst_dmem_U14589 ( .A1(MEM_stage_inst_dmem_n16707), .A2(MEM_stage_inst_dmem_n16706), .ZN(MEM_stage_inst_dmem_n10978) );
NAND2_X1 MEM_stage_inst_dmem_U14588 ( .A1(MEM_stage_inst_dmem_n16777), .A2(MEM_stage_inst_dmem_n16721), .ZN(MEM_stage_inst_dmem_n16706) );
NAND2_X1 MEM_stage_inst_dmem_U14587 ( .A1(MEM_stage_inst_dmem_ram_1703), .A2(MEM_stage_inst_dmem_n16720), .ZN(MEM_stage_inst_dmem_n16707) );
NAND2_X1 MEM_stage_inst_dmem_U14586 ( .A1(MEM_stage_inst_dmem_n16705), .A2(MEM_stage_inst_dmem_n16704), .ZN(MEM_stage_inst_dmem_n10979) );
NAND2_X1 MEM_stage_inst_dmem_U14585 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n16721), .ZN(MEM_stage_inst_dmem_n16704) );
NAND2_X1 MEM_stage_inst_dmem_U14584 ( .A1(MEM_stage_inst_dmem_ram_1704), .A2(MEM_stage_inst_dmem_n16720), .ZN(MEM_stage_inst_dmem_n16705) );
NAND2_X1 MEM_stage_inst_dmem_U14583 ( .A1(MEM_stage_inst_dmem_n16703), .A2(MEM_stage_inst_dmem_n16702), .ZN(MEM_stage_inst_dmem_n10980) );
NAND2_X1 MEM_stage_inst_dmem_U14582 ( .A1(MEM_stage_inst_dmem_n16772), .A2(MEM_stage_inst_dmem_n16721), .ZN(MEM_stage_inst_dmem_n16702) );
NAND2_X1 MEM_stage_inst_dmem_U14581 ( .A1(MEM_stage_inst_dmem_ram_1705), .A2(MEM_stage_inst_dmem_n16720), .ZN(MEM_stage_inst_dmem_n16703) );
NAND2_X1 MEM_stage_inst_dmem_U14580 ( .A1(MEM_stage_inst_dmem_n16701), .A2(MEM_stage_inst_dmem_n16700), .ZN(MEM_stage_inst_dmem_n10981) );
NAND2_X1 MEM_stage_inst_dmem_U14579 ( .A1(MEM_stage_inst_dmem_n16769), .A2(MEM_stage_inst_dmem_n16721), .ZN(MEM_stage_inst_dmem_n16700) );
NAND2_X1 MEM_stage_inst_dmem_U14578 ( .A1(MEM_stage_inst_dmem_ram_1706), .A2(MEM_stage_inst_dmem_n16720), .ZN(MEM_stage_inst_dmem_n16701) );
NAND2_X1 MEM_stage_inst_dmem_U14577 ( .A1(MEM_stage_inst_dmem_n16699), .A2(MEM_stage_inst_dmem_n16698), .ZN(MEM_stage_inst_dmem_n10982) );
NAND2_X1 MEM_stage_inst_dmem_U14576 ( .A1(MEM_stage_inst_dmem_n13044), .A2(MEM_stage_inst_dmem_n16721), .ZN(MEM_stage_inst_dmem_n16698) );
NAND2_X1 MEM_stage_inst_dmem_U14575 ( .A1(MEM_stage_inst_dmem_ram_1707), .A2(MEM_stage_inst_dmem_n16720), .ZN(MEM_stage_inst_dmem_n16699) );
NAND2_X1 MEM_stage_inst_dmem_U14574 ( .A1(MEM_stage_inst_dmem_n16697), .A2(MEM_stage_inst_dmem_n16696), .ZN(MEM_stage_inst_dmem_n10983) );
NAND2_X1 MEM_stage_inst_dmem_U14573 ( .A1(MEM_stage_inst_dmem_n13041), .A2(MEM_stage_inst_dmem_n16721), .ZN(MEM_stage_inst_dmem_n16696) );
NAND2_X1 MEM_stage_inst_dmem_U14572 ( .A1(MEM_stage_inst_dmem_ram_1708), .A2(MEM_stage_inst_dmem_n16720), .ZN(MEM_stage_inst_dmem_n16697) );
NAND2_X1 MEM_stage_inst_dmem_U14571 ( .A1(MEM_stage_inst_dmem_n16695), .A2(MEM_stage_inst_dmem_n16694), .ZN(MEM_stage_inst_dmem_n10984) );
NAND2_X1 MEM_stage_inst_dmem_U14570 ( .A1(EX_pipeline_reg_out_18), .A2(MEM_stage_inst_dmem_n16721), .ZN(MEM_stage_inst_dmem_n16694) );
NAND2_X1 MEM_stage_inst_dmem_U14569 ( .A1(MEM_stage_inst_dmem_ram_1709), .A2(MEM_stage_inst_dmem_n16720), .ZN(MEM_stage_inst_dmem_n16695) );
NAND2_X1 MEM_stage_inst_dmem_U14568 ( .A1(MEM_stage_inst_dmem_n16693), .A2(MEM_stage_inst_dmem_n16692), .ZN(MEM_stage_inst_dmem_n10985) );
NAND2_X1 MEM_stage_inst_dmem_U14567 ( .A1(EX_pipeline_reg_out_19), .A2(MEM_stage_inst_dmem_n16721), .ZN(MEM_stage_inst_dmem_n16692) );
NAND2_X1 MEM_stage_inst_dmem_U14566 ( .A1(MEM_stage_inst_dmem_ram_1710), .A2(MEM_stage_inst_dmem_n16720), .ZN(MEM_stage_inst_dmem_n16693) );
NAND2_X1 MEM_stage_inst_dmem_U14565 ( .A1(MEM_stage_inst_dmem_n16691), .A2(MEM_stage_inst_dmem_n16690), .ZN(MEM_stage_inst_dmem_n10986) );
NAND2_X1 MEM_stage_inst_dmem_U14564 ( .A1(MEM_stage_inst_dmem_n16758), .A2(MEM_stage_inst_dmem_n16721), .ZN(MEM_stage_inst_dmem_n16690) );
INV_X1 MEM_stage_inst_dmem_U14563 ( .A(MEM_stage_inst_dmem_n16720), .ZN(MEM_stage_inst_dmem_n16721) );
NAND2_X1 MEM_stage_inst_dmem_U14562 ( .A1(MEM_stage_inst_dmem_ram_1711), .A2(MEM_stage_inst_dmem_n16720), .ZN(MEM_stage_inst_dmem_n16691) );
NAND2_X1 MEM_stage_inst_dmem_U14561 ( .A1(MEM_stage_inst_dmem_n21109), .A2(MEM_stage_inst_dmem_n17037), .ZN(MEM_stage_inst_dmem_n16720) );
NAND2_X1 MEM_stage_inst_dmem_U14560 ( .A1(MEM_stage_inst_dmem_n16689), .A2(MEM_stage_inst_dmem_n16688), .ZN(MEM_stage_inst_dmem_n10987) );
NAND2_X1 MEM_stage_inst_dmem_U14559 ( .A1(MEM_stage_inst_dmem_n14732), .A2(MEM_stage_inst_dmem_n16687), .ZN(MEM_stage_inst_dmem_n16688) );
NAND2_X1 MEM_stage_inst_dmem_U14558 ( .A1(MEM_stage_inst_dmem_ram_1712), .A2(MEM_stage_inst_dmem_n16686), .ZN(MEM_stage_inst_dmem_n16689) );
NAND2_X1 MEM_stage_inst_dmem_U14557 ( .A1(MEM_stage_inst_dmem_n16685), .A2(MEM_stage_inst_dmem_n16684), .ZN(MEM_stage_inst_dmem_n10988) );
NAND2_X1 MEM_stage_inst_dmem_U14556 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n16687), .ZN(MEM_stage_inst_dmem_n16684) );
NAND2_X1 MEM_stage_inst_dmem_U14555 ( .A1(MEM_stage_inst_dmem_ram_1713), .A2(MEM_stage_inst_dmem_n16686), .ZN(MEM_stage_inst_dmem_n16685) );
NAND2_X1 MEM_stage_inst_dmem_U14554 ( .A1(MEM_stage_inst_dmem_n16683), .A2(MEM_stage_inst_dmem_n16682), .ZN(MEM_stage_inst_dmem_n10989) );
NAND2_X1 MEM_stage_inst_dmem_U14553 ( .A1(MEM_stage_inst_dmem_n16789), .A2(MEM_stage_inst_dmem_n16687), .ZN(MEM_stage_inst_dmem_n16682) );
NAND2_X1 MEM_stage_inst_dmem_U14552 ( .A1(MEM_stage_inst_dmem_ram_1714), .A2(MEM_stage_inst_dmem_n16686), .ZN(MEM_stage_inst_dmem_n16683) );
NAND2_X1 MEM_stage_inst_dmem_U14551 ( .A1(MEM_stage_inst_dmem_n16681), .A2(MEM_stage_inst_dmem_n16680), .ZN(MEM_stage_inst_dmem_n10990) );
NAND2_X1 MEM_stage_inst_dmem_U14550 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n16687), .ZN(MEM_stage_inst_dmem_n16680) );
NAND2_X1 MEM_stage_inst_dmem_U14549 ( .A1(MEM_stage_inst_dmem_ram_1715), .A2(MEM_stage_inst_dmem_n16686), .ZN(MEM_stage_inst_dmem_n16681) );
NAND2_X1 MEM_stage_inst_dmem_U14548 ( .A1(MEM_stage_inst_dmem_n16679), .A2(MEM_stage_inst_dmem_n16678), .ZN(MEM_stage_inst_dmem_n10991) );
NAND2_X1 MEM_stage_inst_dmem_U14547 ( .A1(MEM_stage_inst_dmem_n16784), .A2(MEM_stage_inst_dmem_n16687), .ZN(MEM_stage_inst_dmem_n16678) );
NAND2_X1 MEM_stage_inst_dmem_U14546 ( .A1(MEM_stage_inst_dmem_ram_1716), .A2(MEM_stage_inst_dmem_n16686), .ZN(MEM_stage_inst_dmem_n16679) );
NAND2_X1 MEM_stage_inst_dmem_U14545 ( .A1(MEM_stage_inst_dmem_n16677), .A2(MEM_stage_inst_dmem_n16676), .ZN(MEM_stage_inst_dmem_n10992) );
NAND2_X1 MEM_stage_inst_dmem_U14544 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n16687), .ZN(MEM_stage_inst_dmem_n16676) );
NAND2_X1 MEM_stage_inst_dmem_U14543 ( .A1(MEM_stage_inst_dmem_ram_1717), .A2(MEM_stage_inst_dmem_n16686), .ZN(MEM_stage_inst_dmem_n16677) );
NAND2_X1 MEM_stage_inst_dmem_U14542 ( .A1(MEM_stage_inst_dmem_n16675), .A2(MEM_stage_inst_dmem_n16674), .ZN(MEM_stage_inst_dmem_n10993) );
NAND2_X1 MEM_stage_inst_dmem_U14541 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n16687), .ZN(MEM_stage_inst_dmem_n16674) );
NAND2_X1 MEM_stage_inst_dmem_U14540 ( .A1(MEM_stage_inst_dmem_ram_1718), .A2(MEM_stage_inst_dmem_n16686), .ZN(MEM_stage_inst_dmem_n16675) );
NAND2_X1 MEM_stage_inst_dmem_U14539 ( .A1(MEM_stage_inst_dmem_n16673), .A2(MEM_stage_inst_dmem_n16672), .ZN(MEM_stage_inst_dmem_n10994) );
NAND2_X1 MEM_stage_inst_dmem_U14538 ( .A1(MEM_stage_inst_dmem_n16777), .A2(MEM_stage_inst_dmem_n16687), .ZN(MEM_stage_inst_dmem_n16672) );
NAND2_X1 MEM_stage_inst_dmem_U14537 ( .A1(MEM_stage_inst_dmem_ram_1719), .A2(MEM_stage_inst_dmem_n16686), .ZN(MEM_stage_inst_dmem_n16673) );
NAND2_X1 MEM_stage_inst_dmem_U14536 ( .A1(MEM_stage_inst_dmem_n16671), .A2(MEM_stage_inst_dmem_n16670), .ZN(MEM_stage_inst_dmem_n10995) );
NAND2_X1 MEM_stage_inst_dmem_U14535 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n16687), .ZN(MEM_stage_inst_dmem_n16670) );
NAND2_X1 MEM_stage_inst_dmem_U14534 ( .A1(MEM_stage_inst_dmem_ram_1720), .A2(MEM_stage_inst_dmem_n16686), .ZN(MEM_stage_inst_dmem_n16671) );
NAND2_X1 MEM_stage_inst_dmem_U14533 ( .A1(MEM_stage_inst_dmem_n16669), .A2(MEM_stage_inst_dmem_n16668), .ZN(MEM_stage_inst_dmem_n10996) );
NAND2_X1 MEM_stage_inst_dmem_U14532 ( .A1(MEM_stage_inst_dmem_n16772), .A2(MEM_stage_inst_dmem_n16687), .ZN(MEM_stage_inst_dmem_n16668) );
NAND2_X1 MEM_stage_inst_dmem_U14531 ( .A1(MEM_stage_inst_dmem_ram_1721), .A2(MEM_stage_inst_dmem_n16686), .ZN(MEM_stage_inst_dmem_n16669) );
NAND2_X1 MEM_stage_inst_dmem_U14530 ( .A1(MEM_stage_inst_dmem_n16667), .A2(MEM_stage_inst_dmem_n16666), .ZN(MEM_stage_inst_dmem_n10997) );
NAND2_X1 MEM_stage_inst_dmem_U14529 ( .A1(MEM_stage_inst_dmem_n16769), .A2(MEM_stage_inst_dmem_n16687), .ZN(MEM_stage_inst_dmem_n16666) );
NAND2_X1 MEM_stage_inst_dmem_U14528 ( .A1(MEM_stage_inst_dmem_ram_1722), .A2(MEM_stage_inst_dmem_n16686), .ZN(MEM_stage_inst_dmem_n16667) );
NAND2_X1 MEM_stage_inst_dmem_U14527 ( .A1(MEM_stage_inst_dmem_n16665), .A2(MEM_stage_inst_dmem_n16664), .ZN(MEM_stage_inst_dmem_n10998) );
NAND2_X1 MEM_stage_inst_dmem_U14526 ( .A1(MEM_stage_inst_dmem_n13044), .A2(MEM_stage_inst_dmem_n16687), .ZN(MEM_stage_inst_dmem_n16664) );
NAND2_X1 MEM_stage_inst_dmem_U14525 ( .A1(MEM_stage_inst_dmem_ram_1723), .A2(MEM_stage_inst_dmem_n16686), .ZN(MEM_stage_inst_dmem_n16665) );
NAND2_X1 MEM_stage_inst_dmem_U14524 ( .A1(MEM_stage_inst_dmem_n16663), .A2(MEM_stage_inst_dmem_n16662), .ZN(MEM_stage_inst_dmem_n10999) );
NAND2_X1 MEM_stage_inst_dmem_U14523 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n16687), .ZN(MEM_stage_inst_dmem_n16662) );
NAND2_X1 MEM_stage_inst_dmem_U14522 ( .A1(MEM_stage_inst_dmem_ram_1724), .A2(MEM_stage_inst_dmem_n16686), .ZN(MEM_stage_inst_dmem_n16663) );
NAND2_X1 MEM_stage_inst_dmem_U14521 ( .A1(MEM_stage_inst_dmem_n16661), .A2(MEM_stage_inst_dmem_n16660), .ZN(MEM_stage_inst_dmem_n11000) );
NAND2_X1 MEM_stage_inst_dmem_U14520 ( .A1(MEM_stage_inst_dmem_n116), .A2(MEM_stage_inst_dmem_n16687), .ZN(MEM_stage_inst_dmem_n16660) );
NAND2_X1 MEM_stage_inst_dmem_U14519 ( .A1(MEM_stage_inst_dmem_ram_1725), .A2(MEM_stage_inst_dmem_n16686), .ZN(MEM_stage_inst_dmem_n16661) );
NAND2_X1 MEM_stage_inst_dmem_U14518 ( .A1(MEM_stage_inst_dmem_n16659), .A2(MEM_stage_inst_dmem_n16658), .ZN(MEM_stage_inst_dmem_n11001) );
NAND2_X1 MEM_stage_inst_dmem_U14517 ( .A1(MEM_stage_inst_dmem_n14696), .A2(MEM_stage_inst_dmem_n16687), .ZN(MEM_stage_inst_dmem_n16658) );
NAND2_X1 MEM_stage_inst_dmem_U14516 ( .A1(MEM_stage_inst_dmem_ram_1726), .A2(MEM_stage_inst_dmem_n16686), .ZN(MEM_stage_inst_dmem_n16659) );
NAND2_X1 MEM_stage_inst_dmem_U14515 ( .A1(MEM_stage_inst_dmem_n16657), .A2(MEM_stage_inst_dmem_n16656), .ZN(MEM_stage_inst_dmem_n11002) );
NAND2_X1 MEM_stage_inst_dmem_U14514 ( .A1(MEM_stage_inst_dmem_n16758), .A2(MEM_stage_inst_dmem_n16687), .ZN(MEM_stage_inst_dmem_n16656) );
INV_X1 MEM_stage_inst_dmem_U14513 ( .A(MEM_stage_inst_dmem_n16686), .ZN(MEM_stage_inst_dmem_n16687) );
NAND2_X1 MEM_stage_inst_dmem_U14512 ( .A1(MEM_stage_inst_dmem_ram_1727), .A2(MEM_stage_inst_dmem_n16686), .ZN(MEM_stage_inst_dmem_n16657) );
NAND2_X1 MEM_stage_inst_dmem_U14511 ( .A1(MEM_stage_inst_dmem_n21074), .A2(MEM_stage_inst_dmem_n17037), .ZN(MEM_stage_inst_dmem_n16686) );
NAND2_X1 MEM_stage_inst_dmem_U14510 ( .A1(MEM_stage_inst_dmem_n16655), .A2(MEM_stage_inst_dmem_n16654), .ZN(MEM_stage_inst_dmem_n11003) );
NAND2_X1 MEM_stage_inst_dmem_U14509 ( .A1(MEM_stage_inst_dmem_n20551), .A2(MEM_stage_inst_dmem_n16653), .ZN(MEM_stage_inst_dmem_n16654) );
NAND2_X1 MEM_stage_inst_dmem_U14508 ( .A1(MEM_stage_inst_dmem_ram_1728), .A2(MEM_stage_inst_dmem_n16652), .ZN(MEM_stage_inst_dmem_n16655) );
NAND2_X1 MEM_stage_inst_dmem_U14507 ( .A1(MEM_stage_inst_dmem_n16651), .A2(MEM_stage_inst_dmem_n16650), .ZN(MEM_stage_inst_dmem_n11004) );
NAND2_X1 MEM_stage_inst_dmem_U14506 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n16653), .ZN(MEM_stage_inst_dmem_n16650) );
NAND2_X1 MEM_stage_inst_dmem_U14505 ( .A1(MEM_stage_inst_dmem_ram_1729), .A2(MEM_stage_inst_dmem_n16652), .ZN(MEM_stage_inst_dmem_n16651) );
NAND2_X1 MEM_stage_inst_dmem_U14504 ( .A1(MEM_stage_inst_dmem_n16649), .A2(MEM_stage_inst_dmem_n16648), .ZN(MEM_stage_inst_dmem_n11005) );
NAND2_X1 MEM_stage_inst_dmem_U14503 ( .A1(MEM_stage_inst_dmem_n16789), .A2(MEM_stage_inst_dmem_n16653), .ZN(MEM_stage_inst_dmem_n16648) );
NAND2_X1 MEM_stage_inst_dmem_U14502 ( .A1(MEM_stage_inst_dmem_ram_1730), .A2(MEM_stage_inst_dmem_n16652), .ZN(MEM_stage_inst_dmem_n16649) );
NAND2_X1 MEM_stage_inst_dmem_U14501 ( .A1(MEM_stage_inst_dmem_n16647), .A2(MEM_stage_inst_dmem_n16646), .ZN(MEM_stage_inst_dmem_n11006) );
NAND2_X1 MEM_stage_inst_dmem_U14500 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n16653), .ZN(MEM_stage_inst_dmem_n16646) );
NAND2_X1 MEM_stage_inst_dmem_U14499 ( .A1(MEM_stage_inst_dmem_ram_1731), .A2(MEM_stage_inst_dmem_n16652), .ZN(MEM_stage_inst_dmem_n16647) );
NAND2_X1 MEM_stage_inst_dmem_U14498 ( .A1(MEM_stage_inst_dmem_n16645), .A2(MEM_stage_inst_dmem_n16644), .ZN(MEM_stage_inst_dmem_n11007) );
NAND2_X1 MEM_stage_inst_dmem_U14497 ( .A1(MEM_stage_inst_dmem_n16784), .A2(MEM_stage_inst_dmem_n16653), .ZN(MEM_stage_inst_dmem_n16644) );
NAND2_X1 MEM_stage_inst_dmem_U14496 ( .A1(MEM_stage_inst_dmem_ram_1732), .A2(MEM_stage_inst_dmem_n16652), .ZN(MEM_stage_inst_dmem_n16645) );
NAND2_X1 MEM_stage_inst_dmem_U14495 ( .A1(MEM_stage_inst_dmem_n16643), .A2(MEM_stage_inst_dmem_n16642), .ZN(MEM_stage_inst_dmem_n11008) );
NAND2_X1 MEM_stage_inst_dmem_U14494 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n16653), .ZN(MEM_stage_inst_dmem_n16642) );
NAND2_X1 MEM_stage_inst_dmem_U14493 ( .A1(MEM_stage_inst_dmem_ram_1733), .A2(MEM_stage_inst_dmem_n16652), .ZN(MEM_stage_inst_dmem_n16643) );
NAND2_X1 MEM_stage_inst_dmem_U14492 ( .A1(MEM_stage_inst_dmem_n16641), .A2(MEM_stage_inst_dmem_n16640), .ZN(MEM_stage_inst_dmem_n11009) );
NAND2_X1 MEM_stage_inst_dmem_U14491 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n16653), .ZN(MEM_stage_inst_dmem_n16640) );
NAND2_X1 MEM_stage_inst_dmem_U14490 ( .A1(MEM_stage_inst_dmem_ram_1734), .A2(MEM_stage_inst_dmem_n16652), .ZN(MEM_stage_inst_dmem_n16641) );
NAND2_X1 MEM_stage_inst_dmem_U14489 ( .A1(MEM_stage_inst_dmem_n16639), .A2(MEM_stage_inst_dmem_n16638), .ZN(MEM_stage_inst_dmem_n11010) );
NAND2_X1 MEM_stage_inst_dmem_U14488 ( .A1(MEM_stage_inst_dmem_n16777), .A2(MEM_stage_inst_dmem_n16653), .ZN(MEM_stage_inst_dmem_n16638) );
NAND2_X1 MEM_stage_inst_dmem_U14487 ( .A1(MEM_stage_inst_dmem_ram_1735), .A2(MEM_stage_inst_dmem_n16652), .ZN(MEM_stage_inst_dmem_n16639) );
NAND2_X1 MEM_stage_inst_dmem_U14486 ( .A1(MEM_stage_inst_dmem_n16637), .A2(MEM_stage_inst_dmem_n16636), .ZN(MEM_stage_inst_dmem_n11011) );
NAND2_X1 MEM_stage_inst_dmem_U14485 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n16653), .ZN(MEM_stage_inst_dmem_n16636) );
NAND2_X1 MEM_stage_inst_dmem_U14484 ( .A1(MEM_stage_inst_dmem_ram_1736), .A2(MEM_stage_inst_dmem_n16652), .ZN(MEM_stage_inst_dmem_n16637) );
NAND2_X1 MEM_stage_inst_dmem_U14483 ( .A1(MEM_stage_inst_dmem_n16635), .A2(MEM_stage_inst_dmem_n16634), .ZN(MEM_stage_inst_dmem_n11012) );
NAND2_X1 MEM_stage_inst_dmem_U14482 ( .A1(MEM_stage_inst_dmem_n16772), .A2(MEM_stage_inst_dmem_n16653), .ZN(MEM_stage_inst_dmem_n16634) );
NAND2_X1 MEM_stage_inst_dmem_U14481 ( .A1(MEM_stage_inst_dmem_ram_1737), .A2(MEM_stage_inst_dmem_n16652), .ZN(MEM_stage_inst_dmem_n16635) );
NAND2_X1 MEM_stage_inst_dmem_U14480 ( .A1(MEM_stage_inst_dmem_n16633), .A2(MEM_stage_inst_dmem_n16632), .ZN(MEM_stage_inst_dmem_n11013) );
NAND2_X1 MEM_stage_inst_dmem_U14479 ( .A1(MEM_stage_inst_dmem_n16769), .A2(MEM_stage_inst_dmem_n16653), .ZN(MEM_stage_inst_dmem_n16632) );
NAND2_X1 MEM_stage_inst_dmem_U14478 ( .A1(MEM_stage_inst_dmem_ram_1738), .A2(MEM_stage_inst_dmem_n16652), .ZN(MEM_stage_inst_dmem_n16633) );
NAND2_X1 MEM_stage_inst_dmem_U14477 ( .A1(MEM_stage_inst_dmem_n16631), .A2(MEM_stage_inst_dmem_n16630), .ZN(MEM_stage_inst_dmem_n11014) );
NAND2_X1 MEM_stage_inst_dmem_U14476 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n16653), .ZN(MEM_stage_inst_dmem_n16630) );
NAND2_X1 MEM_stage_inst_dmem_U14475 ( .A1(MEM_stage_inst_dmem_ram_1739), .A2(MEM_stage_inst_dmem_n16652), .ZN(MEM_stage_inst_dmem_n16631) );
NAND2_X1 MEM_stage_inst_dmem_U14474 ( .A1(MEM_stage_inst_dmem_n16629), .A2(MEM_stage_inst_dmem_n16628), .ZN(MEM_stage_inst_dmem_n11015) );
NAND2_X1 MEM_stage_inst_dmem_U14473 ( .A1(MEM_stage_inst_dmem_n21474), .A2(MEM_stage_inst_dmem_n16653), .ZN(MEM_stage_inst_dmem_n16628) );
NAND2_X1 MEM_stage_inst_dmem_U14472 ( .A1(MEM_stage_inst_dmem_ram_1740), .A2(MEM_stage_inst_dmem_n16652), .ZN(MEM_stage_inst_dmem_n16629) );
NAND2_X1 MEM_stage_inst_dmem_U14471 ( .A1(MEM_stage_inst_dmem_n16627), .A2(MEM_stage_inst_dmem_n16626), .ZN(MEM_stage_inst_dmem_n11016) );
NAND2_X1 MEM_stage_inst_dmem_U14470 ( .A1(MEM_stage_inst_dmem_n20512), .A2(MEM_stage_inst_dmem_n16653), .ZN(MEM_stage_inst_dmem_n16626) );
NAND2_X1 MEM_stage_inst_dmem_U14469 ( .A1(MEM_stage_inst_dmem_ram_1741), .A2(MEM_stage_inst_dmem_n16652), .ZN(MEM_stage_inst_dmem_n16627) );
NAND2_X1 MEM_stage_inst_dmem_U14468 ( .A1(MEM_stage_inst_dmem_n16625), .A2(MEM_stage_inst_dmem_n16624), .ZN(MEM_stage_inst_dmem_n11017) );
NAND2_X1 MEM_stage_inst_dmem_U14467 ( .A1(MEM_stage_inst_dmem_n20509), .A2(MEM_stage_inst_dmem_n16653), .ZN(MEM_stage_inst_dmem_n16624) );
NAND2_X1 MEM_stage_inst_dmem_U14466 ( .A1(MEM_stage_inst_dmem_ram_1742), .A2(MEM_stage_inst_dmem_n16652), .ZN(MEM_stage_inst_dmem_n16625) );
NAND2_X1 MEM_stage_inst_dmem_U14465 ( .A1(MEM_stage_inst_dmem_n16623), .A2(MEM_stage_inst_dmem_n16622), .ZN(MEM_stage_inst_dmem_n11018) );
NAND2_X1 MEM_stage_inst_dmem_U14464 ( .A1(MEM_stage_inst_dmem_n16758), .A2(MEM_stage_inst_dmem_n16653), .ZN(MEM_stage_inst_dmem_n16622) );
INV_X1 MEM_stage_inst_dmem_U14463 ( .A(MEM_stage_inst_dmem_n16652), .ZN(MEM_stage_inst_dmem_n16653) );
NAND2_X1 MEM_stage_inst_dmem_U14462 ( .A1(MEM_stage_inst_dmem_ram_1743), .A2(MEM_stage_inst_dmem_n16652), .ZN(MEM_stage_inst_dmem_n16623) );
NAND2_X1 MEM_stage_inst_dmem_U14461 ( .A1(MEM_stage_inst_dmem_n21039), .A2(MEM_stage_inst_dmem_n17037), .ZN(MEM_stage_inst_dmem_n16652) );
NAND2_X1 MEM_stage_inst_dmem_U14460 ( .A1(MEM_stage_inst_dmem_n16621), .A2(MEM_stage_inst_dmem_n16620), .ZN(MEM_stage_inst_dmem_n11019) );
NAND2_X1 MEM_stage_inst_dmem_U14459 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n16619), .ZN(MEM_stage_inst_dmem_n16620) );
NAND2_X1 MEM_stage_inst_dmem_U14458 ( .A1(MEM_stage_inst_dmem_ram_1744), .A2(MEM_stage_inst_dmem_n16618), .ZN(MEM_stage_inst_dmem_n16621) );
NAND2_X1 MEM_stage_inst_dmem_U14457 ( .A1(MEM_stage_inst_dmem_n16617), .A2(MEM_stage_inst_dmem_n16616), .ZN(MEM_stage_inst_dmem_n11020) );
NAND2_X1 MEM_stage_inst_dmem_U14456 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n16619), .ZN(MEM_stage_inst_dmem_n16616) );
NAND2_X1 MEM_stage_inst_dmem_U14455 ( .A1(MEM_stage_inst_dmem_ram_1745), .A2(MEM_stage_inst_dmem_n16618), .ZN(MEM_stage_inst_dmem_n16617) );
NAND2_X1 MEM_stage_inst_dmem_U14454 ( .A1(MEM_stage_inst_dmem_n16615), .A2(MEM_stage_inst_dmem_n16614), .ZN(MEM_stage_inst_dmem_n11021) );
NAND2_X1 MEM_stage_inst_dmem_U14453 ( .A1(MEM_stage_inst_dmem_n16789), .A2(MEM_stage_inst_dmem_n16619), .ZN(MEM_stage_inst_dmem_n16614) );
NAND2_X1 MEM_stage_inst_dmem_U14452 ( .A1(MEM_stage_inst_dmem_ram_1746), .A2(MEM_stage_inst_dmem_n16618), .ZN(MEM_stage_inst_dmem_n16615) );
NAND2_X1 MEM_stage_inst_dmem_U14451 ( .A1(MEM_stage_inst_dmem_n16613), .A2(MEM_stage_inst_dmem_n16612), .ZN(MEM_stage_inst_dmem_n11022) );
NAND2_X1 MEM_stage_inst_dmem_U14450 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n16619), .ZN(MEM_stage_inst_dmem_n16612) );
NAND2_X1 MEM_stage_inst_dmem_U14449 ( .A1(MEM_stage_inst_dmem_ram_1747), .A2(MEM_stage_inst_dmem_n16618), .ZN(MEM_stage_inst_dmem_n16613) );
NAND2_X1 MEM_stage_inst_dmem_U14448 ( .A1(MEM_stage_inst_dmem_n16611), .A2(MEM_stage_inst_dmem_n16610), .ZN(MEM_stage_inst_dmem_n11023) );
NAND2_X1 MEM_stage_inst_dmem_U14447 ( .A1(MEM_stage_inst_dmem_n16784), .A2(MEM_stage_inst_dmem_n16619), .ZN(MEM_stage_inst_dmem_n16610) );
NAND2_X1 MEM_stage_inst_dmem_U14446 ( .A1(MEM_stage_inst_dmem_ram_1748), .A2(MEM_stage_inst_dmem_n16618), .ZN(MEM_stage_inst_dmem_n16611) );
NAND2_X1 MEM_stage_inst_dmem_U14445 ( .A1(MEM_stage_inst_dmem_n16609), .A2(MEM_stage_inst_dmem_n16608), .ZN(MEM_stage_inst_dmem_n11024) );
NAND2_X1 MEM_stage_inst_dmem_U14444 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n16619), .ZN(MEM_stage_inst_dmem_n16608) );
NAND2_X1 MEM_stage_inst_dmem_U14443 ( .A1(MEM_stage_inst_dmem_ram_1749), .A2(MEM_stage_inst_dmem_n16618), .ZN(MEM_stage_inst_dmem_n16609) );
NAND2_X1 MEM_stage_inst_dmem_U14442 ( .A1(MEM_stage_inst_dmem_n16607), .A2(MEM_stage_inst_dmem_n16606), .ZN(MEM_stage_inst_dmem_n11025) );
NAND2_X1 MEM_stage_inst_dmem_U14441 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n16619), .ZN(MEM_stage_inst_dmem_n16606) );
NAND2_X1 MEM_stage_inst_dmem_U14440 ( .A1(MEM_stage_inst_dmem_ram_1750), .A2(MEM_stage_inst_dmem_n16618), .ZN(MEM_stage_inst_dmem_n16607) );
NAND2_X1 MEM_stage_inst_dmem_U14439 ( .A1(MEM_stage_inst_dmem_n16605), .A2(MEM_stage_inst_dmem_n16604), .ZN(MEM_stage_inst_dmem_n11026) );
NAND2_X1 MEM_stage_inst_dmem_U14438 ( .A1(MEM_stage_inst_dmem_n16777), .A2(MEM_stage_inst_dmem_n16619), .ZN(MEM_stage_inst_dmem_n16604) );
NAND2_X1 MEM_stage_inst_dmem_U14437 ( .A1(MEM_stage_inst_dmem_ram_1751), .A2(MEM_stage_inst_dmem_n16618), .ZN(MEM_stage_inst_dmem_n16605) );
NAND2_X1 MEM_stage_inst_dmem_U14436 ( .A1(MEM_stage_inst_dmem_n16603), .A2(MEM_stage_inst_dmem_n16602), .ZN(MEM_stage_inst_dmem_n11027) );
NAND2_X1 MEM_stage_inst_dmem_U14435 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n16619), .ZN(MEM_stage_inst_dmem_n16602) );
NAND2_X1 MEM_stage_inst_dmem_U14434 ( .A1(MEM_stage_inst_dmem_ram_1752), .A2(MEM_stage_inst_dmem_n16618), .ZN(MEM_stage_inst_dmem_n16603) );
NAND2_X1 MEM_stage_inst_dmem_U14433 ( .A1(MEM_stage_inst_dmem_n16601), .A2(MEM_stage_inst_dmem_n16600), .ZN(MEM_stage_inst_dmem_n11028) );
NAND2_X1 MEM_stage_inst_dmem_U14432 ( .A1(MEM_stage_inst_dmem_n16772), .A2(MEM_stage_inst_dmem_n16619), .ZN(MEM_stage_inst_dmem_n16600) );
NAND2_X1 MEM_stage_inst_dmem_U14431 ( .A1(MEM_stage_inst_dmem_ram_1753), .A2(MEM_stage_inst_dmem_n16618), .ZN(MEM_stage_inst_dmem_n16601) );
NAND2_X1 MEM_stage_inst_dmem_U14430 ( .A1(MEM_stage_inst_dmem_n16599), .A2(MEM_stage_inst_dmem_n16598), .ZN(MEM_stage_inst_dmem_n11029) );
NAND2_X1 MEM_stage_inst_dmem_U14429 ( .A1(MEM_stage_inst_dmem_n16769), .A2(MEM_stage_inst_dmem_n16619), .ZN(MEM_stage_inst_dmem_n16598) );
NAND2_X1 MEM_stage_inst_dmem_U14428 ( .A1(MEM_stage_inst_dmem_ram_1754), .A2(MEM_stage_inst_dmem_n16618), .ZN(MEM_stage_inst_dmem_n16599) );
NAND2_X1 MEM_stage_inst_dmem_U14427 ( .A1(MEM_stage_inst_dmem_n16597), .A2(MEM_stage_inst_dmem_n16596), .ZN(MEM_stage_inst_dmem_n11030) );
NAND2_X1 MEM_stage_inst_dmem_U14426 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n16619), .ZN(MEM_stage_inst_dmem_n16596) );
NAND2_X1 MEM_stage_inst_dmem_U14425 ( .A1(MEM_stage_inst_dmem_ram_1755), .A2(MEM_stage_inst_dmem_n16618), .ZN(MEM_stage_inst_dmem_n16597) );
NAND2_X1 MEM_stage_inst_dmem_U14424 ( .A1(MEM_stage_inst_dmem_n16595), .A2(MEM_stage_inst_dmem_n16594), .ZN(MEM_stage_inst_dmem_n11031) );
NAND2_X1 MEM_stage_inst_dmem_U14423 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n16619), .ZN(MEM_stage_inst_dmem_n16594) );
NAND2_X1 MEM_stage_inst_dmem_U14422 ( .A1(MEM_stage_inst_dmem_ram_1756), .A2(MEM_stage_inst_dmem_n16618), .ZN(MEM_stage_inst_dmem_n16595) );
NAND2_X1 MEM_stage_inst_dmem_U14421 ( .A1(MEM_stage_inst_dmem_n16593), .A2(MEM_stage_inst_dmem_n16592), .ZN(MEM_stage_inst_dmem_n11032) );
NAND2_X1 MEM_stage_inst_dmem_U14420 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n16619), .ZN(MEM_stage_inst_dmem_n16592) );
NAND2_X1 MEM_stage_inst_dmem_U14419 ( .A1(MEM_stage_inst_dmem_ram_1757), .A2(MEM_stage_inst_dmem_n16618), .ZN(MEM_stage_inst_dmem_n16593) );
NAND2_X1 MEM_stage_inst_dmem_U14418 ( .A1(MEM_stage_inst_dmem_n16591), .A2(MEM_stage_inst_dmem_n16590), .ZN(MEM_stage_inst_dmem_n11033) );
NAND2_X1 MEM_stage_inst_dmem_U14417 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n16619), .ZN(MEM_stage_inst_dmem_n16590) );
NAND2_X1 MEM_stage_inst_dmem_U14416 ( .A1(MEM_stage_inst_dmem_ram_1758), .A2(MEM_stage_inst_dmem_n16618), .ZN(MEM_stage_inst_dmem_n16591) );
NAND2_X1 MEM_stage_inst_dmem_U14415 ( .A1(MEM_stage_inst_dmem_n16589), .A2(MEM_stage_inst_dmem_n16588), .ZN(MEM_stage_inst_dmem_n11034) );
NAND2_X1 MEM_stage_inst_dmem_U14414 ( .A1(MEM_stage_inst_dmem_n16758), .A2(MEM_stage_inst_dmem_n16619), .ZN(MEM_stage_inst_dmem_n16588) );
NAND2_X1 MEM_stage_inst_dmem_U14413 ( .A1(MEM_stage_inst_dmem_ram_1759), .A2(MEM_stage_inst_dmem_n16618), .ZN(MEM_stage_inst_dmem_n16589) );
NAND2_X1 MEM_stage_inst_dmem_U14412 ( .A1(MEM_stage_inst_dmem_n21004), .A2(MEM_stage_inst_dmem_n17037), .ZN(MEM_stage_inst_dmem_n16618) );
NAND2_X1 MEM_stage_inst_dmem_U14411 ( .A1(MEM_stage_inst_dmem_n16587), .A2(MEM_stage_inst_dmem_n16586), .ZN(MEM_stage_inst_dmem_n11035) );
NAND2_X1 MEM_stage_inst_dmem_U14410 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n16585), .ZN(MEM_stage_inst_dmem_n16586) );
NAND2_X1 MEM_stage_inst_dmem_U14409 ( .A1(MEM_stage_inst_dmem_ram_1760), .A2(MEM_stage_inst_dmem_n16584), .ZN(MEM_stage_inst_dmem_n16587) );
NAND2_X1 MEM_stage_inst_dmem_U14408 ( .A1(MEM_stage_inst_dmem_n16583), .A2(MEM_stage_inst_dmem_n16582), .ZN(MEM_stage_inst_dmem_n11036) );
NAND2_X1 MEM_stage_inst_dmem_U14407 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n16585), .ZN(MEM_stage_inst_dmem_n16582) );
NAND2_X1 MEM_stage_inst_dmem_U14406 ( .A1(MEM_stage_inst_dmem_ram_1761), .A2(MEM_stage_inst_dmem_n16584), .ZN(MEM_stage_inst_dmem_n16583) );
NAND2_X1 MEM_stage_inst_dmem_U14405 ( .A1(MEM_stage_inst_dmem_n16581), .A2(MEM_stage_inst_dmem_n16580), .ZN(MEM_stage_inst_dmem_n11037) );
NAND2_X1 MEM_stage_inst_dmem_U14404 ( .A1(MEM_stage_inst_dmem_n16789), .A2(MEM_stage_inst_dmem_n16585), .ZN(MEM_stage_inst_dmem_n16580) );
NAND2_X1 MEM_stage_inst_dmem_U14403 ( .A1(MEM_stage_inst_dmem_ram_1762), .A2(MEM_stage_inst_dmem_n16584), .ZN(MEM_stage_inst_dmem_n16581) );
NAND2_X1 MEM_stage_inst_dmem_U14402 ( .A1(MEM_stage_inst_dmem_n16579), .A2(MEM_stage_inst_dmem_n16578), .ZN(MEM_stage_inst_dmem_n11038) );
NAND2_X1 MEM_stage_inst_dmem_U14401 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n16585), .ZN(MEM_stage_inst_dmem_n16578) );
NAND2_X1 MEM_stage_inst_dmem_U14400 ( .A1(MEM_stage_inst_dmem_ram_1763), .A2(MEM_stage_inst_dmem_n16584), .ZN(MEM_stage_inst_dmem_n16579) );
NAND2_X1 MEM_stage_inst_dmem_U14399 ( .A1(MEM_stage_inst_dmem_n16577), .A2(MEM_stage_inst_dmem_n16576), .ZN(MEM_stage_inst_dmem_n11039) );
NAND2_X1 MEM_stage_inst_dmem_U14398 ( .A1(MEM_stage_inst_dmem_n16784), .A2(MEM_stage_inst_dmem_n16585), .ZN(MEM_stage_inst_dmem_n16576) );
NAND2_X1 MEM_stage_inst_dmem_U14397 ( .A1(MEM_stage_inst_dmem_ram_1764), .A2(MEM_stage_inst_dmem_n16584), .ZN(MEM_stage_inst_dmem_n16577) );
NAND2_X1 MEM_stage_inst_dmem_U14396 ( .A1(MEM_stage_inst_dmem_n16575), .A2(MEM_stage_inst_dmem_n16574), .ZN(MEM_stage_inst_dmem_n11040) );
NAND2_X1 MEM_stage_inst_dmem_U14395 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n16585), .ZN(MEM_stage_inst_dmem_n16574) );
NAND2_X1 MEM_stage_inst_dmem_U14394 ( .A1(MEM_stage_inst_dmem_ram_1765), .A2(MEM_stage_inst_dmem_n16584), .ZN(MEM_stage_inst_dmem_n16575) );
NAND2_X1 MEM_stage_inst_dmem_U14393 ( .A1(MEM_stage_inst_dmem_n16573), .A2(MEM_stage_inst_dmem_n16572), .ZN(MEM_stage_inst_dmem_n11041) );
NAND2_X1 MEM_stage_inst_dmem_U14392 ( .A1(MEM_stage_inst_dmem_n14717), .A2(MEM_stage_inst_dmem_n16585), .ZN(MEM_stage_inst_dmem_n16572) );
NAND2_X1 MEM_stage_inst_dmem_U14391 ( .A1(MEM_stage_inst_dmem_ram_1766), .A2(MEM_stage_inst_dmem_n16584), .ZN(MEM_stage_inst_dmem_n16573) );
NAND2_X1 MEM_stage_inst_dmem_U14390 ( .A1(MEM_stage_inst_dmem_n16571), .A2(MEM_stage_inst_dmem_n16570), .ZN(MEM_stage_inst_dmem_n11042) );
NAND2_X1 MEM_stage_inst_dmem_U14389 ( .A1(MEM_stage_inst_dmem_n16777), .A2(MEM_stage_inst_dmem_n16585), .ZN(MEM_stage_inst_dmem_n16570) );
NAND2_X1 MEM_stage_inst_dmem_U14388 ( .A1(MEM_stage_inst_dmem_ram_1767), .A2(MEM_stage_inst_dmem_n16584), .ZN(MEM_stage_inst_dmem_n16571) );
NAND2_X1 MEM_stage_inst_dmem_U14387 ( .A1(MEM_stage_inst_dmem_n16569), .A2(MEM_stage_inst_dmem_n16568), .ZN(MEM_stage_inst_dmem_n11043) );
NAND2_X1 MEM_stage_inst_dmem_U14386 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n16585), .ZN(MEM_stage_inst_dmem_n16568) );
NAND2_X1 MEM_stage_inst_dmem_U14385 ( .A1(MEM_stage_inst_dmem_ram_1768), .A2(MEM_stage_inst_dmem_n16584), .ZN(MEM_stage_inst_dmem_n16569) );
NAND2_X1 MEM_stage_inst_dmem_U14384 ( .A1(MEM_stage_inst_dmem_n16567), .A2(MEM_stage_inst_dmem_n16566), .ZN(MEM_stage_inst_dmem_n11044) );
NAND2_X1 MEM_stage_inst_dmem_U14383 ( .A1(MEM_stage_inst_dmem_n16772), .A2(MEM_stage_inst_dmem_n16585), .ZN(MEM_stage_inst_dmem_n16566) );
NAND2_X1 MEM_stage_inst_dmem_U14382 ( .A1(MEM_stage_inst_dmem_ram_1769), .A2(MEM_stage_inst_dmem_n16584), .ZN(MEM_stage_inst_dmem_n16567) );
NAND2_X1 MEM_stage_inst_dmem_U14381 ( .A1(MEM_stage_inst_dmem_n16565), .A2(MEM_stage_inst_dmem_n16564), .ZN(MEM_stage_inst_dmem_n11045) );
NAND2_X1 MEM_stage_inst_dmem_U14380 ( .A1(MEM_stage_inst_dmem_n16769), .A2(MEM_stage_inst_dmem_n16585), .ZN(MEM_stage_inst_dmem_n16564) );
NAND2_X1 MEM_stage_inst_dmem_U14379 ( .A1(MEM_stage_inst_dmem_ram_1770), .A2(MEM_stage_inst_dmem_n16584), .ZN(MEM_stage_inst_dmem_n16565) );
NAND2_X1 MEM_stage_inst_dmem_U14378 ( .A1(MEM_stage_inst_dmem_n16563), .A2(MEM_stage_inst_dmem_n16562), .ZN(MEM_stage_inst_dmem_n11046) );
NAND2_X1 MEM_stage_inst_dmem_U14377 ( .A1(MEM_stage_inst_dmem_n20904), .A2(MEM_stage_inst_dmem_n16585), .ZN(MEM_stage_inst_dmem_n16562) );
NAND2_X1 MEM_stage_inst_dmem_U14376 ( .A1(MEM_stage_inst_dmem_ram_1771), .A2(MEM_stage_inst_dmem_n16584), .ZN(MEM_stage_inst_dmem_n16563) );
NAND2_X1 MEM_stage_inst_dmem_U14375 ( .A1(MEM_stage_inst_dmem_n16561), .A2(MEM_stage_inst_dmem_n16560), .ZN(MEM_stage_inst_dmem_n11047) );
NAND2_X1 MEM_stage_inst_dmem_U14374 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n16585), .ZN(MEM_stage_inst_dmem_n16560) );
NAND2_X1 MEM_stage_inst_dmem_U14373 ( .A1(MEM_stage_inst_dmem_ram_1772), .A2(MEM_stage_inst_dmem_n16584), .ZN(MEM_stage_inst_dmem_n16561) );
NAND2_X1 MEM_stage_inst_dmem_U14372 ( .A1(MEM_stage_inst_dmem_n16559), .A2(MEM_stage_inst_dmem_n16558), .ZN(MEM_stage_inst_dmem_n11048) );
NAND2_X1 MEM_stage_inst_dmem_U14371 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n16585), .ZN(MEM_stage_inst_dmem_n16558) );
NAND2_X1 MEM_stage_inst_dmem_U14370 ( .A1(MEM_stage_inst_dmem_ram_1773), .A2(MEM_stage_inst_dmem_n16584), .ZN(MEM_stage_inst_dmem_n16559) );
NAND2_X1 MEM_stage_inst_dmem_U14369 ( .A1(MEM_stage_inst_dmem_n16557), .A2(MEM_stage_inst_dmem_n16556), .ZN(MEM_stage_inst_dmem_n11049) );
NAND2_X1 MEM_stage_inst_dmem_U14368 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n16585), .ZN(MEM_stage_inst_dmem_n16556) );
NAND2_X1 MEM_stage_inst_dmem_U14367 ( .A1(MEM_stage_inst_dmem_ram_1774), .A2(MEM_stage_inst_dmem_n16584), .ZN(MEM_stage_inst_dmem_n16557) );
NAND2_X1 MEM_stage_inst_dmem_U14366 ( .A1(MEM_stage_inst_dmem_n16555), .A2(MEM_stage_inst_dmem_n16554), .ZN(MEM_stage_inst_dmem_n11050) );
NAND2_X1 MEM_stage_inst_dmem_U14365 ( .A1(MEM_stage_inst_dmem_n16758), .A2(MEM_stage_inst_dmem_n16585), .ZN(MEM_stage_inst_dmem_n16554) );
INV_X1 MEM_stage_inst_dmem_U14364 ( .A(MEM_stage_inst_dmem_n16584), .ZN(MEM_stage_inst_dmem_n16585) );
NAND2_X1 MEM_stage_inst_dmem_U14363 ( .A1(MEM_stage_inst_dmem_ram_1775), .A2(MEM_stage_inst_dmem_n16584), .ZN(MEM_stage_inst_dmem_n16555) );
NAND2_X1 MEM_stage_inst_dmem_U14362 ( .A1(MEM_stage_inst_dmem_n20969), .A2(MEM_stage_inst_dmem_n17037), .ZN(MEM_stage_inst_dmem_n16584) );
NAND2_X1 MEM_stage_inst_dmem_U14361 ( .A1(MEM_stage_inst_dmem_n16553), .A2(MEM_stage_inst_dmem_n16552), .ZN(MEM_stage_inst_dmem_n11051) );
NAND2_X1 MEM_stage_inst_dmem_U14360 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n16551), .ZN(MEM_stage_inst_dmem_n16552) );
NAND2_X1 MEM_stage_inst_dmem_U14359 ( .A1(MEM_stage_inst_dmem_ram_1776), .A2(MEM_stage_inst_dmem_n16550), .ZN(MEM_stage_inst_dmem_n16553) );
NAND2_X1 MEM_stage_inst_dmem_U14358 ( .A1(MEM_stage_inst_dmem_n16549), .A2(MEM_stage_inst_dmem_n16548), .ZN(MEM_stage_inst_dmem_n11052) );
NAND2_X1 MEM_stage_inst_dmem_U14357 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n16551), .ZN(MEM_stage_inst_dmem_n16548) );
NAND2_X1 MEM_stage_inst_dmem_U14356 ( .A1(MEM_stage_inst_dmem_ram_1777), .A2(MEM_stage_inst_dmem_n16550), .ZN(MEM_stage_inst_dmem_n16549) );
NAND2_X1 MEM_stage_inst_dmem_U14355 ( .A1(MEM_stage_inst_dmem_n16547), .A2(MEM_stage_inst_dmem_n16546), .ZN(MEM_stage_inst_dmem_n11053) );
NAND2_X1 MEM_stage_inst_dmem_U14354 ( .A1(MEM_stage_inst_dmem_n16789), .A2(MEM_stage_inst_dmem_n16551), .ZN(MEM_stage_inst_dmem_n16546) );
NAND2_X1 MEM_stage_inst_dmem_U14353 ( .A1(MEM_stage_inst_dmem_ram_1778), .A2(MEM_stage_inst_dmem_n16550), .ZN(MEM_stage_inst_dmem_n16547) );
NAND2_X1 MEM_stage_inst_dmem_U14352 ( .A1(MEM_stage_inst_dmem_n16545), .A2(MEM_stage_inst_dmem_n16544), .ZN(MEM_stage_inst_dmem_n11054) );
NAND2_X1 MEM_stage_inst_dmem_U14351 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n16551), .ZN(MEM_stage_inst_dmem_n16544) );
NAND2_X1 MEM_stage_inst_dmem_U14350 ( .A1(MEM_stage_inst_dmem_ram_1779), .A2(MEM_stage_inst_dmem_n16550), .ZN(MEM_stage_inst_dmem_n16545) );
NAND2_X1 MEM_stage_inst_dmem_U14349 ( .A1(MEM_stage_inst_dmem_n16543), .A2(MEM_stage_inst_dmem_n16542), .ZN(MEM_stage_inst_dmem_n11055) );
NAND2_X1 MEM_stage_inst_dmem_U14348 ( .A1(MEM_stage_inst_dmem_n16784), .A2(MEM_stage_inst_dmem_n16551), .ZN(MEM_stage_inst_dmem_n16542) );
NAND2_X1 MEM_stage_inst_dmem_U14347 ( .A1(MEM_stage_inst_dmem_ram_1780), .A2(MEM_stage_inst_dmem_n16550), .ZN(MEM_stage_inst_dmem_n16543) );
NAND2_X1 MEM_stage_inst_dmem_U14346 ( .A1(MEM_stage_inst_dmem_n16541), .A2(MEM_stage_inst_dmem_n16540), .ZN(MEM_stage_inst_dmem_n11056) );
NAND2_X1 MEM_stage_inst_dmem_U14345 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n16551), .ZN(MEM_stage_inst_dmem_n16540) );
NAND2_X1 MEM_stage_inst_dmem_U14344 ( .A1(MEM_stage_inst_dmem_ram_1781), .A2(MEM_stage_inst_dmem_n16550), .ZN(MEM_stage_inst_dmem_n16541) );
NAND2_X1 MEM_stage_inst_dmem_U14343 ( .A1(MEM_stage_inst_dmem_n16539), .A2(MEM_stage_inst_dmem_n16538), .ZN(MEM_stage_inst_dmem_n11057) );
NAND2_X1 MEM_stage_inst_dmem_U14342 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n16551), .ZN(MEM_stage_inst_dmem_n16538) );
NAND2_X1 MEM_stage_inst_dmem_U14341 ( .A1(MEM_stage_inst_dmem_ram_1782), .A2(MEM_stage_inst_dmem_n16550), .ZN(MEM_stage_inst_dmem_n16539) );
NAND2_X1 MEM_stage_inst_dmem_U14340 ( .A1(MEM_stage_inst_dmem_n16537), .A2(MEM_stage_inst_dmem_n16536), .ZN(MEM_stage_inst_dmem_n11058) );
NAND2_X1 MEM_stage_inst_dmem_U14339 ( .A1(MEM_stage_inst_dmem_n16777), .A2(MEM_stage_inst_dmem_n16551), .ZN(MEM_stage_inst_dmem_n16536) );
NAND2_X1 MEM_stage_inst_dmem_U14338 ( .A1(MEM_stage_inst_dmem_ram_1783), .A2(MEM_stage_inst_dmem_n16550), .ZN(MEM_stage_inst_dmem_n16537) );
NAND2_X1 MEM_stage_inst_dmem_U14337 ( .A1(MEM_stage_inst_dmem_n16535), .A2(MEM_stage_inst_dmem_n16534), .ZN(MEM_stage_inst_dmem_n11059) );
NAND2_X1 MEM_stage_inst_dmem_U14336 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n16551), .ZN(MEM_stage_inst_dmem_n16534) );
NAND2_X1 MEM_stage_inst_dmem_U14335 ( .A1(MEM_stage_inst_dmem_ram_1784), .A2(MEM_stage_inst_dmem_n16550), .ZN(MEM_stage_inst_dmem_n16535) );
NAND2_X1 MEM_stage_inst_dmem_U14334 ( .A1(MEM_stage_inst_dmem_n16533), .A2(MEM_stage_inst_dmem_n16532), .ZN(MEM_stage_inst_dmem_n11060) );
NAND2_X1 MEM_stage_inst_dmem_U14333 ( .A1(MEM_stage_inst_dmem_n16772), .A2(MEM_stage_inst_dmem_n16551), .ZN(MEM_stage_inst_dmem_n16532) );
NAND2_X1 MEM_stage_inst_dmem_U14332 ( .A1(MEM_stage_inst_dmem_ram_1785), .A2(MEM_stage_inst_dmem_n16550), .ZN(MEM_stage_inst_dmem_n16533) );
NAND2_X1 MEM_stage_inst_dmem_U14331 ( .A1(MEM_stage_inst_dmem_n16531), .A2(MEM_stage_inst_dmem_n16530), .ZN(MEM_stage_inst_dmem_n11061) );
NAND2_X1 MEM_stage_inst_dmem_U14330 ( .A1(MEM_stage_inst_dmem_n16769), .A2(MEM_stage_inst_dmem_n16551), .ZN(MEM_stage_inst_dmem_n16530) );
NAND2_X1 MEM_stage_inst_dmem_U14329 ( .A1(MEM_stage_inst_dmem_ram_1786), .A2(MEM_stage_inst_dmem_n16550), .ZN(MEM_stage_inst_dmem_n16531) );
NAND2_X1 MEM_stage_inst_dmem_U14328 ( .A1(MEM_stage_inst_dmem_n16529), .A2(MEM_stage_inst_dmem_n16528), .ZN(MEM_stage_inst_dmem_n11062) );
NAND2_X1 MEM_stage_inst_dmem_U14327 ( .A1(MEM_stage_inst_dmem_n18004), .A2(MEM_stage_inst_dmem_n16551), .ZN(MEM_stage_inst_dmem_n16528) );
NAND2_X1 MEM_stage_inst_dmem_U14326 ( .A1(MEM_stage_inst_dmem_ram_1787), .A2(MEM_stage_inst_dmem_n16550), .ZN(MEM_stage_inst_dmem_n16529) );
NAND2_X1 MEM_stage_inst_dmem_U14325 ( .A1(MEM_stage_inst_dmem_n16527), .A2(MEM_stage_inst_dmem_n16526), .ZN(MEM_stage_inst_dmem_n11063) );
NAND2_X1 MEM_stage_inst_dmem_U14324 ( .A1(MEM_stage_inst_dmem_n18001), .A2(MEM_stage_inst_dmem_n16551), .ZN(MEM_stage_inst_dmem_n16526) );
NAND2_X1 MEM_stage_inst_dmem_U14323 ( .A1(MEM_stage_inst_dmem_ram_1788), .A2(MEM_stage_inst_dmem_n16550), .ZN(MEM_stage_inst_dmem_n16527) );
NAND2_X1 MEM_stage_inst_dmem_U14322 ( .A1(MEM_stage_inst_dmem_n16525), .A2(MEM_stage_inst_dmem_n16524), .ZN(MEM_stage_inst_dmem_n11064) );
NAND2_X1 MEM_stage_inst_dmem_U14321 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n16551), .ZN(MEM_stage_inst_dmem_n16524) );
NAND2_X1 MEM_stage_inst_dmem_U14320 ( .A1(MEM_stage_inst_dmem_ram_1789), .A2(MEM_stage_inst_dmem_n16550), .ZN(MEM_stage_inst_dmem_n16525) );
NAND2_X1 MEM_stage_inst_dmem_U14319 ( .A1(MEM_stage_inst_dmem_n16523), .A2(MEM_stage_inst_dmem_n16522), .ZN(MEM_stage_inst_dmem_n11065) );
NAND2_X1 MEM_stage_inst_dmem_U14318 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n16551), .ZN(MEM_stage_inst_dmem_n16522) );
NAND2_X1 MEM_stage_inst_dmem_U14317 ( .A1(MEM_stage_inst_dmem_ram_1790), .A2(MEM_stage_inst_dmem_n16550), .ZN(MEM_stage_inst_dmem_n16523) );
NAND2_X1 MEM_stage_inst_dmem_U14316 ( .A1(MEM_stage_inst_dmem_n16521), .A2(MEM_stage_inst_dmem_n16520), .ZN(MEM_stage_inst_dmem_n11066) );
NAND2_X1 MEM_stage_inst_dmem_U14315 ( .A1(MEM_stage_inst_dmem_n16758), .A2(MEM_stage_inst_dmem_n16551), .ZN(MEM_stage_inst_dmem_n16520) );
INV_X1 MEM_stage_inst_dmem_U14314 ( .A(MEM_stage_inst_dmem_n16550), .ZN(MEM_stage_inst_dmem_n16551) );
NAND2_X1 MEM_stage_inst_dmem_U14313 ( .A1(MEM_stage_inst_dmem_ram_1791), .A2(MEM_stage_inst_dmem_n16550), .ZN(MEM_stage_inst_dmem_n16521) );
NAND2_X1 MEM_stage_inst_dmem_U14312 ( .A1(MEM_stage_inst_dmem_n20934), .A2(MEM_stage_inst_dmem_n17037), .ZN(MEM_stage_inst_dmem_n16550) );
NOR2_X2 MEM_stage_inst_dmem_U14311 ( .A1(MEM_stage_inst_dmem_n16519), .A2(MEM_stage_inst_dmem_n20933), .ZN(MEM_stage_inst_dmem_n17037) );
NAND2_X1 MEM_stage_inst_dmem_U14310 ( .A1(MEM_stage_inst_dmem_n16518), .A2(MEM_stage_inst_dmem_n16517), .ZN(MEM_stage_inst_dmem_n11067) );
NAND2_X1 MEM_stage_inst_dmem_U14309 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n16516), .ZN(MEM_stage_inst_dmem_n16517) );
NAND2_X1 MEM_stage_inst_dmem_U14308 ( .A1(MEM_stage_inst_dmem_ram_1792), .A2(MEM_stage_inst_dmem_n16515), .ZN(MEM_stage_inst_dmem_n16518) );
NAND2_X1 MEM_stage_inst_dmem_U14307 ( .A1(MEM_stage_inst_dmem_n16514), .A2(MEM_stage_inst_dmem_n16513), .ZN(MEM_stage_inst_dmem_n11068) );
NAND2_X1 MEM_stage_inst_dmem_U14306 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n16516), .ZN(MEM_stage_inst_dmem_n16513) );
NAND2_X1 MEM_stage_inst_dmem_U14305 ( .A1(MEM_stage_inst_dmem_ram_1793), .A2(MEM_stage_inst_dmem_n16515), .ZN(MEM_stage_inst_dmem_n16514) );
NAND2_X1 MEM_stage_inst_dmem_U14304 ( .A1(MEM_stage_inst_dmem_n16512), .A2(MEM_stage_inst_dmem_n16511), .ZN(MEM_stage_inst_dmem_n11069) );
NAND2_X1 MEM_stage_inst_dmem_U14303 ( .A1(MEM_stage_inst_dmem_n16789), .A2(MEM_stage_inst_dmem_n16516), .ZN(MEM_stage_inst_dmem_n16511) );
NAND2_X1 MEM_stage_inst_dmem_U14302 ( .A1(MEM_stage_inst_dmem_ram_1794), .A2(MEM_stage_inst_dmem_n16515), .ZN(MEM_stage_inst_dmem_n16512) );
NAND2_X1 MEM_stage_inst_dmem_U14301 ( .A1(MEM_stage_inst_dmem_n16510), .A2(MEM_stage_inst_dmem_n16509), .ZN(MEM_stage_inst_dmem_n11070) );
NAND2_X1 MEM_stage_inst_dmem_U14300 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n16516), .ZN(MEM_stage_inst_dmem_n16509) );
NAND2_X1 MEM_stage_inst_dmem_U14299 ( .A1(MEM_stage_inst_dmem_ram_1795), .A2(MEM_stage_inst_dmem_n16515), .ZN(MEM_stage_inst_dmem_n16510) );
NAND2_X1 MEM_stage_inst_dmem_U14298 ( .A1(MEM_stage_inst_dmem_n16508), .A2(MEM_stage_inst_dmem_n16507), .ZN(MEM_stage_inst_dmem_n11071) );
NAND2_X1 MEM_stage_inst_dmem_U14297 ( .A1(MEM_stage_inst_dmem_n16784), .A2(MEM_stage_inst_dmem_n16516), .ZN(MEM_stage_inst_dmem_n16507) );
NAND2_X1 MEM_stage_inst_dmem_U14296 ( .A1(MEM_stage_inst_dmem_ram_1796), .A2(MEM_stage_inst_dmem_n16515), .ZN(MEM_stage_inst_dmem_n16508) );
NAND2_X1 MEM_stage_inst_dmem_U14295 ( .A1(MEM_stage_inst_dmem_n16506), .A2(MEM_stage_inst_dmem_n16505), .ZN(MEM_stage_inst_dmem_n11072) );
NAND2_X1 MEM_stage_inst_dmem_U14294 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n16516), .ZN(MEM_stage_inst_dmem_n16505) );
NAND2_X1 MEM_stage_inst_dmem_U14293 ( .A1(MEM_stage_inst_dmem_ram_1797), .A2(MEM_stage_inst_dmem_n16515), .ZN(MEM_stage_inst_dmem_n16506) );
NAND2_X1 MEM_stage_inst_dmem_U14292 ( .A1(MEM_stage_inst_dmem_n16504), .A2(MEM_stage_inst_dmem_n16503), .ZN(MEM_stage_inst_dmem_n11073) );
NAND2_X1 MEM_stage_inst_dmem_U14291 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n16516), .ZN(MEM_stage_inst_dmem_n16503) );
NAND2_X1 MEM_stage_inst_dmem_U14290 ( .A1(MEM_stage_inst_dmem_ram_1798), .A2(MEM_stage_inst_dmem_n16515), .ZN(MEM_stage_inst_dmem_n16504) );
NAND2_X1 MEM_stage_inst_dmem_U14289 ( .A1(MEM_stage_inst_dmem_n16502), .A2(MEM_stage_inst_dmem_n16501), .ZN(MEM_stage_inst_dmem_n11074) );
NAND2_X1 MEM_stage_inst_dmem_U14288 ( .A1(MEM_stage_inst_dmem_n16777), .A2(MEM_stage_inst_dmem_n16516), .ZN(MEM_stage_inst_dmem_n16501) );
NAND2_X1 MEM_stage_inst_dmem_U14287 ( .A1(MEM_stage_inst_dmem_ram_1799), .A2(MEM_stage_inst_dmem_n16515), .ZN(MEM_stage_inst_dmem_n16502) );
NAND2_X1 MEM_stage_inst_dmem_U14286 ( .A1(MEM_stage_inst_dmem_n16500), .A2(MEM_stage_inst_dmem_n16499), .ZN(MEM_stage_inst_dmem_n11075) );
NAND2_X1 MEM_stage_inst_dmem_U14285 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n16516), .ZN(MEM_stage_inst_dmem_n16499) );
NAND2_X1 MEM_stage_inst_dmem_U14284 ( .A1(MEM_stage_inst_dmem_ram_1800), .A2(MEM_stage_inst_dmem_n16515), .ZN(MEM_stage_inst_dmem_n16500) );
NAND2_X1 MEM_stage_inst_dmem_U14283 ( .A1(MEM_stage_inst_dmem_n16498), .A2(MEM_stage_inst_dmem_n16497), .ZN(MEM_stage_inst_dmem_n11076) );
NAND2_X1 MEM_stage_inst_dmem_U14282 ( .A1(MEM_stage_inst_dmem_n16772), .A2(MEM_stage_inst_dmem_n16516), .ZN(MEM_stage_inst_dmem_n16497) );
NAND2_X1 MEM_stage_inst_dmem_U14281 ( .A1(MEM_stage_inst_dmem_ram_1801), .A2(MEM_stage_inst_dmem_n16515), .ZN(MEM_stage_inst_dmem_n16498) );
NAND2_X1 MEM_stage_inst_dmem_U14280 ( .A1(MEM_stage_inst_dmem_n16496), .A2(MEM_stage_inst_dmem_n16495), .ZN(MEM_stage_inst_dmem_n11077) );
NAND2_X1 MEM_stage_inst_dmem_U14279 ( .A1(MEM_stage_inst_dmem_n16769), .A2(MEM_stage_inst_dmem_n16516), .ZN(MEM_stage_inst_dmem_n16495) );
NAND2_X1 MEM_stage_inst_dmem_U14278 ( .A1(MEM_stage_inst_dmem_ram_1802), .A2(MEM_stage_inst_dmem_n16515), .ZN(MEM_stage_inst_dmem_n16496) );
NAND2_X1 MEM_stage_inst_dmem_U14277 ( .A1(MEM_stage_inst_dmem_n16494), .A2(MEM_stage_inst_dmem_n16493), .ZN(MEM_stage_inst_dmem_n11078) );
NAND2_X1 MEM_stage_inst_dmem_U14276 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n16516), .ZN(MEM_stage_inst_dmem_n16493) );
NAND2_X1 MEM_stage_inst_dmem_U14275 ( .A1(MEM_stage_inst_dmem_ram_1803), .A2(MEM_stage_inst_dmem_n16515), .ZN(MEM_stage_inst_dmem_n16494) );
NAND2_X1 MEM_stage_inst_dmem_U14274 ( .A1(MEM_stage_inst_dmem_n16492), .A2(MEM_stage_inst_dmem_n16491), .ZN(MEM_stage_inst_dmem_n11079) );
NAND2_X1 MEM_stage_inst_dmem_U14273 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n16516), .ZN(MEM_stage_inst_dmem_n16491) );
NAND2_X1 MEM_stage_inst_dmem_U14272 ( .A1(MEM_stage_inst_dmem_ram_1804), .A2(MEM_stage_inst_dmem_n16515), .ZN(MEM_stage_inst_dmem_n16492) );
NAND2_X1 MEM_stage_inst_dmem_U14271 ( .A1(MEM_stage_inst_dmem_n16490), .A2(MEM_stage_inst_dmem_n16489), .ZN(MEM_stage_inst_dmem_n11080) );
NAND2_X1 MEM_stage_inst_dmem_U14270 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n16516), .ZN(MEM_stage_inst_dmem_n16489) );
NAND2_X1 MEM_stage_inst_dmem_U14269 ( .A1(MEM_stage_inst_dmem_ram_1805), .A2(MEM_stage_inst_dmem_n16515), .ZN(MEM_stage_inst_dmem_n16490) );
NAND2_X1 MEM_stage_inst_dmem_U14268 ( .A1(MEM_stage_inst_dmem_n16488), .A2(MEM_stage_inst_dmem_n16487), .ZN(MEM_stage_inst_dmem_n11081) );
NAND2_X1 MEM_stage_inst_dmem_U14267 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n16516), .ZN(MEM_stage_inst_dmem_n16487) );
NAND2_X1 MEM_stage_inst_dmem_U14266 ( .A1(MEM_stage_inst_dmem_ram_1806), .A2(MEM_stage_inst_dmem_n16515), .ZN(MEM_stage_inst_dmem_n16488) );
NAND2_X1 MEM_stage_inst_dmem_U14265 ( .A1(MEM_stage_inst_dmem_n16486), .A2(MEM_stage_inst_dmem_n16485), .ZN(MEM_stage_inst_dmem_n11082) );
NAND2_X1 MEM_stage_inst_dmem_U14264 ( .A1(MEM_stage_inst_dmem_n16758), .A2(MEM_stage_inst_dmem_n16516), .ZN(MEM_stage_inst_dmem_n16485) );
INV_X1 MEM_stage_inst_dmem_U14263 ( .A(MEM_stage_inst_dmem_n16515), .ZN(MEM_stage_inst_dmem_n16516) );
NAND2_X1 MEM_stage_inst_dmem_U14262 ( .A1(MEM_stage_inst_dmem_ram_1807), .A2(MEM_stage_inst_dmem_n16515), .ZN(MEM_stage_inst_dmem_n16486) );
NAND2_X1 MEM_stage_inst_dmem_U14261 ( .A1(MEM_stage_inst_dmem_n21465), .A2(MEM_stage_inst_dmem_n16484), .ZN(MEM_stage_inst_dmem_n16515) );
NAND2_X1 MEM_stage_inst_dmem_U14260 ( .A1(MEM_stage_inst_dmem_n16483), .A2(MEM_stage_inst_dmem_n16482), .ZN(MEM_stage_inst_dmem_n11083) );
NAND2_X1 MEM_stage_inst_dmem_U14259 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n16481), .ZN(MEM_stage_inst_dmem_n16482) );
NAND2_X1 MEM_stage_inst_dmem_U14258 ( .A1(MEM_stage_inst_dmem_ram_1808), .A2(MEM_stage_inst_dmem_n16480), .ZN(MEM_stage_inst_dmem_n16483) );
NAND2_X1 MEM_stage_inst_dmem_U14257 ( .A1(MEM_stage_inst_dmem_n16479), .A2(MEM_stage_inst_dmem_n16478), .ZN(MEM_stage_inst_dmem_n11084) );
NAND2_X1 MEM_stage_inst_dmem_U14256 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n16481), .ZN(MEM_stage_inst_dmem_n16478) );
NAND2_X1 MEM_stage_inst_dmem_U14255 ( .A1(MEM_stage_inst_dmem_ram_1809), .A2(MEM_stage_inst_dmem_n16480), .ZN(MEM_stage_inst_dmem_n16479) );
NAND2_X1 MEM_stage_inst_dmem_U14254 ( .A1(MEM_stage_inst_dmem_n16477), .A2(MEM_stage_inst_dmem_n16476), .ZN(MEM_stage_inst_dmem_n11085) );
NAND2_X1 MEM_stage_inst_dmem_U14253 ( .A1(MEM_stage_inst_dmem_n16789), .A2(MEM_stage_inst_dmem_n16481), .ZN(MEM_stage_inst_dmem_n16476) );
NAND2_X1 MEM_stage_inst_dmem_U14252 ( .A1(MEM_stage_inst_dmem_ram_1810), .A2(MEM_stage_inst_dmem_n16480), .ZN(MEM_stage_inst_dmem_n16477) );
NAND2_X1 MEM_stage_inst_dmem_U14251 ( .A1(MEM_stage_inst_dmem_n16475), .A2(MEM_stage_inst_dmem_n16474), .ZN(MEM_stage_inst_dmem_n11086) );
NAND2_X1 MEM_stage_inst_dmem_U14250 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n16481), .ZN(MEM_stage_inst_dmem_n16474) );
NAND2_X1 MEM_stage_inst_dmem_U14249 ( .A1(MEM_stage_inst_dmem_ram_1811), .A2(MEM_stage_inst_dmem_n16480), .ZN(MEM_stage_inst_dmem_n16475) );
NAND2_X1 MEM_stage_inst_dmem_U14248 ( .A1(MEM_stage_inst_dmem_n16473), .A2(MEM_stage_inst_dmem_n16472), .ZN(MEM_stage_inst_dmem_n11087) );
NAND2_X1 MEM_stage_inst_dmem_U14247 ( .A1(MEM_stage_inst_dmem_n16784), .A2(MEM_stage_inst_dmem_n16481), .ZN(MEM_stage_inst_dmem_n16472) );
NAND2_X1 MEM_stage_inst_dmem_U14246 ( .A1(MEM_stage_inst_dmem_ram_1812), .A2(MEM_stage_inst_dmem_n16480), .ZN(MEM_stage_inst_dmem_n16473) );
NAND2_X1 MEM_stage_inst_dmem_U14245 ( .A1(MEM_stage_inst_dmem_n16471), .A2(MEM_stage_inst_dmem_n16470), .ZN(MEM_stage_inst_dmem_n11088) );
NAND2_X1 MEM_stage_inst_dmem_U14244 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n16481), .ZN(MEM_stage_inst_dmem_n16470) );
NAND2_X1 MEM_stage_inst_dmem_U14243 ( .A1(MEM_stage_inst_dmem_ram_1813), .A2(MEM_stage_inst_dmem_n16480), .ZN(MEM_stage_inst_dmem_n16471) );
NAND2_X1 MEM_stage_inst_dmem_U14242 ( .A1(MEM_stage_inst_dmem_n16469), .A2(MEM_stage_inst_dmem_n16468), .ZN(MEM_stage_inst_dmem_n11089) );
NAND2_X1 MEM_stage_inst_dmem_U14241 ( .A1(MEM_stage_inst_dmem_n21340), .A2(MEM_stage_inst_dmem_n16481), .ZN(MEM_stage_inst_dmem_n16468) );
NAND2_X1 MEM_stage_inst_dmem_U14240 ( .A1(MEM_stage_inst_dmem_ram_1814), .A2(MEM_stage_inst_dmem_n16480), .ZN(MEM_stage_inst_dmem_n16469) );
NAND2_X1 MEM_stage_inst_dmem_U14239 ( .A1(MEM_stage_inst_dmem_n16467), .A2(MEM_stage_inst_dmem_n16466), .ZN(MEM_stage_inst_dmem_n11090) );
NAND2_X1 MEM_stage_inst_dmem_U14238 ( .A1(MEM_stage_inst_dmem_n16777), .A2(MEM_stage_inst_dmem_n16481), .ZN(MEM_stage_inst_dmem_n16466) );
NAND2_X1 MEM_stage_inst_dmem_U14237 ( .A1(MEM_stage_inst_dmem_ram_1815), .A2(MEM_stage_inst_dmem_n16480), .ZN(MEM_stage_inst_dmem_n16467) );
NAND2_X1 MEM_stage_inst_dmem_U14236 ( .A1(MEM_stage_inst_dmem_n16465), .A2(MEM_stage_inst_dmem_n16464), .ZN(MEM_stage_inst_dmem_n11091) );
NAND2_X1 MEM_stage_inst_dmem_U14235 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n16481), .ZN(MEM_stage_inst_dmem_n16464) );
NAND2_X1 MEM_stage_inst_dmem_U14234 ( .A1(MEM_stage_inst_dmem_ram_1816), .A2(MEM_stage_inst_dmem_n16480), .ZN(MEM_stage_inst_dmem_n16465) );
NAND2_X1 MEM_stage_inst_dmem_U14233 ( .A1(MEM_stage_inst_dmem_n16463), .A2(MEM_stage_inst_dmem_n16462), .ZN(MEM_stage_inst_dmem_n11092) );
NAND2_X1 MEM_stage_inst_dmem_U14232 ( .A1(MEM_stage_inst_dmem_n16772), .A2(MEM_stage_inst_dmem_n16481), .ZN(MEM_stage_inst_dmem_n16462) );
NAND2_X1 MEM_stage_inst_dmem_U14231 ( .A1(MEM_stage_inst_dmem_ram_1817), .A2(MEM_stage_inst_dmem_n16480), .ZN(MEM_stage_inst_dmem_n16463) );
NAND2_X1 MEM_stage_inst_dmem_U14230 ( .A1(MEM_stage_inst_dmem_n16461), .A2(MEM_stage_inst_dmem_n16460), .ZN(MEM_stage_inst_dmem_n11093) );
NAND2_X1 MEM_stage_inst_dmem_U14229 ( .A1(MEM_stage_inst_dmem_n16769), .A2(MEM_stage_inst_dmem_n16481), .ZN(MEM_stage_inst_dmem_n16460) );
NAND2_X1 MEM_stage_inst_dmem_U14228 ( .A1(MEM_stage_inst_dmem_ram_1818), .A2(MEM_stage_inst_dmem_n16480), .ZN(MEM_stage_inst_dmem_n16461) );
NAND2_X1 MEM_stage_inst_dmem_U14227 ( .A1(MEM_stage_inst_dmem_n16459), .A2(MEM_stage_inst_dmem_n16458), .ZN(MEM_stage_inst_dmem_n11094) );
NAND2_X1 MEM_stage_inst_dmem_U14226 ( .A1(MEM_stage_inst_dmem_n18864), .A2(MEM_stage_inst_dmem_n16481), .ZN(MEM_stage_inst_dmem_n16458) );
NAND2_X1 MEM_stage_inst_dmem_U14225 ( .A1(MEM_stage_inst_dmem_ram_1819), .A2(MEM_stage_inst_dmem_n16480), .ZN(MEM_stage_inst_dmem_n16459) );
NAND2_X1 MEM_stage_inst_dmem_U14224 ( .A1(MEM_stage_inst_dmem_n16457), .A2(MEM_stage_inst_dmem_n16456), .ZN(MEM_stage_inst_dmem_n11095) );
NAND2_X1 MEM_stage_inst_dmem_U14223 ( .A1(MEM_stage_inst_dmem_n18861), .A2(MEM_stage_inst_dmem_n16481), .ZN(MEM_stage_inst_dmem_n16456) );
NAND2_X1 MEM_stage_inst_dmem_U14222 ( .A1(MEM_stage_inst_dmem_ram_1820), .A2(MEM_stage_inst_dmem_n16480), .ZN(MEM_stage_inst_dmem_n16457) );
NAND2_X1 MEM_stage_inst_dmem_U14221 ( .A1(MEM_stage_inst_dmem_n16455), .A2(MEM_stage_inst_dmem_n16454), .ZN(MEM_stage_inst_dmem_n11096) );
NAND2_X1 MEM_stage_inst_dmem_U14220 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n16481), .ZN(MEM_stage_inst_dmem_n16454) );
NAND2_X1 MEM_stage_inst_dmem_U14219 ( .A1(MEM_stage_inst_dmem_ram_1821), .A2(MEM_stage_inst_dmem_n16480), .ZN(MEM_stage_inst_dmem_n16455) );
NAND2_X1 MEM_stage_inst_dmem_U14218 ( .A1(MEM_stage_inst_dmem_n16453), .A2(MEM_stage_inst_dmem_n16452), .ZN(MEM_stage_inst_dmem_n11097) );
NAND2_X1 MEM_stage_inst_dmem_U14217 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n16481), .ZN(MEM_stage_inst_dmem_n16452) );
NAND2_X1 MEM_stage_inst_dmem_U14216 ( .A1(MEM_stage_inst_dmem_ram_1822), .A2(MEM_stage_inst_dmem_n16480), .ZN(MEM_stage_inst_dmem_n16453) );
NAND2_X1 MEM_stage_inst_dmem_U14215 ( .A1(MEM_stage_inst_dmem_n16451), .A2(MEM_stage_inst_dmem_n16450), .ZN(MEM_stage_inst_dmem_n11098) );
NAND2_X1 MEM_stage_inst_dmem_U14214 ( .A1(MEM_stage_inst_dmem_n16758), .A2(MEM_stage_inst_dmem_n16481), .ZN(MEM_stage_inst_dmem_n16450) );
INV_X1 MEM_stage_inst_dmem_U14213 ( .A(MEM_stage_inst_dmem_n16480), .ZN(MEM_stage_inst_dmem_n16481) );
NAND2_X1 MEM_stage_inst_dmem_U14212 ( .A1(MEM_stage_inst_dmem_ram_1823), .A2(MEM_stage_inst_dmem_n16480), .ZN(MEM_stage_inst_dmem_n16451) );
NAND2_X1 MEM_stage_inst_dmem_U14211 ( .A1(MEM_stage_inst_dmem_n21429), .A2(MEM_stage_inst_dmem_n16484), .ZN(MEM_stage_inst_dmem_n16480) );
NAND2_X1 MEM_stage_inst_dmem_U14210 ( .A1(MEM_stage_inst_dmem_n16449), .A2(MEM_stage_inst_dmem_n16448), .ZN(MEM_stage_inst_dmem_n11099) );
NAND2_X1 MEM_stage_inst_dmem_U14209 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n16447), .ZN(MEM_stage_inst_dmem_n16448) );
NAND2_X1 MEM_stage_inst_dmem_U14208 ( .A1(MEM_stage_inst_dmem_ram_1824), .A2(MEM_stage_inst_dmem_n16446), .ZN(MEM_stage_inst_dmem_n16449) );
NAND2_X1 MEM_stage_inst_dmem_U14207 ( .A1(MEM_stage_inst_dmem_n16445), .A2(MEM_stage_inst_dmem_n16444), .ZN(MEM_stage_inst_dmem_n11100) );
NAND2_X1 MEM_stage_inst_dmem_U14206 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n16447), .ZN(MEM_stage_inst_dmem_n16444) );
NAND2_X1 MEM_stage_inst_dmem_U14205 ( .A1(MEM_stage_inst_dmem_ram_1825), .A2(MEM_stage_inst_dmem_n16446), .ZN(MEM_stage_inst_dmem_n16445) );
NAND2_X1 MEM_stage_inst_dmem_U14204 ( .A1(MEM_stage_inst_dmem_n16443), .A2(MEM_stage_inst_dmem_n16442), .ZN(MEM_stage_inst_dmem_n11101) );
NAND2_X1 MEM_stage_inst_dmem_U14203 ( .A1(MEM_stage_inst_dmem_n16789), .A2(MEM_stage_inst_dmem_n16447), .ZN(MEM_stage_inst_dmem_n16442) );
NAND2_X1 MEM_stage_inst_dmem_U14202 ( .A1(MEM_stage_inst_dmem_ram_1826), .A2(MEM_stage_inst_dmem_n16446), .ZN(MEM_stage_inst_dmem_n16443) );
NAND2_X1 MEM_stage_inst_dmem_U14201 ( .A1(MEM_stage_inst_dmem_n16441), .A2(MEM_stage_inst_dmem_n16440), .ZN(MEM_stage_inst_dmem_n11102) );
NAND2_X1 MEM_stage_inst_dmem_U14200 ( .A1(EX_pipeline_reg_out_8), .A2(MEM_stage_inst_dmem_n16447), .ZN(MEM_stage_inst_dmem_n16440) );
NAND2_X1 MEM_stage_inst_dmem_U14199 ( .A1(MEM_stage_inst_dmem_ram_1827), .A2(MEM_stage_inst_dmem_n16446), .ZN(MEM_stage_inst_dmem_n16441) );
NAND2_X1 MEM_stage_inst_dmem_U14198 ( .A1(MEM_stage_inst_dmem_n16439), .A2(MEM_stage_inst_dmem_n16438), .ZN(MEM_stage_inst_dmem_n11103) );
NAND2_X1 MEM_stage_inst_dmem_U14197 ( .A1(MEM_stage_inst_dmem_n16784), .A2(MEM_stage_inst_dmem_n16447), .ZN(MEM_stage_inst_dmem_n16438) );
NAND2_X1 MEM_stage_inst_dmem_U14196 ( .A1(MEM_stage_inst_dmem_ram_1828), .A2(MEM_stage_inst_dmem_n16446), .ZN(MEM_stage_inst_dmem_n16439) );
NAND2_X1 MEM_stage_inst_dmem_U14195 ( .A1(MEM_stage_inst_dmem_n16437), .A2(MEM_stage_inst_dmem_n16436), .ZN(MEM_stage_inst_dmem_n11104) );
NAND2_X1 MEM_stage_inst_dmem_U14194 ( .A1(EX_pipeline_reg_out_10), .A2(MEM_stage_inst_dmem_n16447), .ZN(MEM_stage_inst_dmem_n16436) );
NAND2_X1 MEM_stage_inst_dmem_U14193 ( .A1(MEM_stage_inst_dmem_ram_1829), .A2(MEM_stage_inst_dmem_n16446), .ZN(MEM_stage_inst_dmem_n16437) );
NAND2_X1 MEM_stage_inst_dmem_U14192 ( .A1(MEM_stage_inst_dmem_n16435), .A2(MEM_stage_inst_dmem_n16434), .ZN(MEM_stage_inst_dmem_n11105) );
NAND2_X1 MEM_stage_inst_dmem_U14191 ( .A1(EX_pipeline_reg_out_11), .A2(MEM_stage_inst_dmem_n16447), .ZN(MEM_stage_inst_dmem_n16434) );
NAND2_X1 MEM_stage_inst_dmem_U14190 ( .A1(MEM_stage_inst_dmem_ram_1830), .A2(MEM_stage_inst_dmem_n16446), .ZN(MEM_stage_inst_dmem_n16435) );
NAND2_X1 MEM_stage_inst_dmem_U14189 ( .A1(MEM_stage_inst_dmem_n16433), .A2(MEM_stage_inst_dmem_n16432), .ZN(MEM_stage_inst_dmem_n11106) );
NAND2_X1 MEM_stage_inst_dmem_U14188 ( .A1(MEM_stage_inst_dmem_n16777), .A2(MEM_stage_inst_dmem_n16447), .ZN(MEM_stage_inst_dmem_n16432) );
NAND2_X1 MEM_stage_inst_dmem_U14187 ( .A1(MEM_stage_inst_dmem_ram_1831), .A2(MEM_stage_inst_dmem_n16446), .ZN(MEM_stage_inst_dmem_n16433) );
NAND2_X1 MEM_stage_inst_dmem_U14186 ( .A1(MEM_stage_inst_dmem_n16431), .A2(MEM_stage_inst_dmem_n16430), .ZN(MEM_stage_inst_dmem_n11107) );
NAND2_X1 MEM_stage_inst_dmem_U14185 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n16447), .ZN(MEM_stage_inst_dmem_n16430) );
NAND2_X1 MEM_stage_inst_dmem_U14184 ( .A1(MEM_stage_inst_dmem_ram_1832), .A2(MEM_stage_inst_dmem_n16446), .ZN(MEM_stage_inst_dmem_n16431) );
NAND2_X1 MEM_stage_inst_dmem_U14183 ( .A1(MEM_stage_inst_dmem_n16429), .A2(MEM_stage_inst_dmem_n16428), .ZN(MEM_stage_inst_dmem_n11108) );
NAND2_X1 MEM_stage_inst_dmem_U14182 ( .A1(MEM_stage_inst_dmem_n16772), .A2(MEM_stage_inst_dmem_n16447), .ZN(MEM_stage_inst_dmem_n16428) );
NAND2_X1 MEM_stage_inst_dmem_U14181 ( .A1(MEM_stage_inst_dmem_ram_1833), .A2(MEM_stage_inst_dmem_n16446), .ZN(MEM_stage_inst_dmem_n16429) );
NAND2_X1 MEM_stage_inst_dmem_U14180 ( .A1(MEM_stage_inst_dmem_n16427), .A2(MEM_stage_inst_dmem_n16426), .ZN(MEM_stage_inst_dmem_n11109) );
NAND2_X1 MEM_stage_inst_dmem_U14179 ( .A1(MEM_stage_inst_dmem_n16769), .A2(MEM_stage_inst_dmem_n16447), .ZN(MEM_stage_inst_dmem_n16426) );
NAND2_X1 MEM_stage_inst_dmem_U14178 ( .A1(MEM_stage_inst_dmem_ram_1834), .A2(MEM_stage_inst_dmem_n16446), .ZN(MEM_stage_inst_dmem_n16427) );
NAND2_X1 MEM_stage_inst_dmem_U14177 ( .A1(MEM_stage_inst_dmem_n16425), .A2(MEM_stage_inst_dmem_n16424), .ZN(MEM_stage_inst_dmem_n11110) );
NAND2_X1 MEM_stage_inst_dmem_U14176 ( .A1(EX_pipeline_reg_out_16), .A2(MEM_stage_inst_dmem_n16447), .ZN(MEM_stage_inst_dmem_n16424) );
NAND2_X1 MEM_stage_inst_dmem_U14175 ( .A1(MEM_stage_inst_dmem_ram_1835), .A2(MEM_stage_inst_dmem_n16446), .ZN(MEM_stage_inst_dmem_n16425) );
NAND2_X1 MEM_stage_inst_dmem_U14174 ( .A1(MEM_stage_inst_dmem_n16423), .A2(MEM_stage_inst_dmem_n16422), .ZN(MEM_stage_inst_dmem_n11111) );
NAND2_X1 MEM_stage_inst_dmem_U14173 ( .A1(EX_pipeline_reg_out_17), .A2(MEM_stage_inst_dmem_n16447), .ZN(MEM_stage_inst_dmem_n16422) );
NAND2_X1 MEM_stage_inst_dmem_U14172 ( .A1(MEM_stage_inst_dmem_ram_1836), .A2(MEM_stage_inst_dmem_n16446), .ZN(MEM_stage_inst_dmem_n16423) );
NAND2_X1 MEM_stage_inst_dmem_U14171 ( .A1(MEM_stage_inst_dmem_n16421), .A2(MEM_stage_inst_dmem_n16420), .ZN(MEM_stage_inst_dmem_n11112) );
NAND2_X1 MEM_stage_inst_dmem_U14170 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n16447), .ZN(MEM_stage_inst_dmem_n16420) );
NAND2_X1 MEM_stage_inst_dmem_U14169 ( .A1(MEM_stage_inst_dmem_ram_1837), .A2(MEM_stage_inst_dmem_n16446), .ZN(MEM_stage_inst_dmem_n16421) );
NAND2_X1 MEM_stage_inst_dmem_U14168 ( .A1(MEM_stage_inst_dmem_n16419), .A2(MEM_stage_inst_dmem_n16418), .ZN(MEM_stage_inst_dmem_n11113) );
NAND2_X1 MEM_stage_inst_dmem_U14167 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n16447), .ZN(MEM_stage_inst_dmem_n16418) );
NAND2_X1 MEM_stage_inst_dmem_U14166 ( .A1(MEM_stage_inst_dmem_ram_1838), .A2(MEM_stage_inst_dmem_n16446), .ZN(MEM_stage_inst_dmem_n16419) );
NAND2_X1 MEM_stage_inst_dmem_U14165 ( .A1(MEM_stage_inst_dmem_n16417), .A2(MEM_stage_inst_dmem_n16416), .ZN(MEM_stage_inst_dmem_n11114) );
NAND2_X1 MEM_stage_inst_dmem_U14164 ( .A1(MEM_stage_inst_dmem_n16758), .A2(MEM_stage_inst_dmem_n16447), .ZN(MEM_stage_inst_dmem_n16416) );
INV_X1 MEM_stage_inst_dmem_U14163 ( .A(MEM_stage_inst_dmem_n16446), .ZN(MEM_stage_inst_dmem_n16447) );
NAND2_X1 MEM_stage_inst_dmem_U14162 ( .A1(MEM_stage_inst_dmem_ram_1839), .A2(MEM_stage_inst_dmem_n16446), .ZN(MEM_stage_inst_dmem_n16417) );
NAND2_X1 MEM_stage_inst_dmem_U14161 ( .A1(MEM_stage_inst_dmem_n21394), .A2(MEM_stage_inst_dmem_n16484), .ZN(MEM_stage_inst_dmem_n16446) );
NAND2_X1 MEM_stage_inst_dmem_U14160 ( .A1(MEM_stage_inst_dmem_n16415), .A2(MEM_stage_inst_dmem_n16414), .ZN(MEM_stage_inst_dmem_n11115) );
NAND2_X1 MEM_stage_inst_dmem_U14159 ( .A1(MEM_stage_inst_dmem_n15145), .A2(MEM_stage_inst_dmem_n16413), .ZN(MEM_stage_inst_dmem_n16414) );
NAND2_X1 MEM_stage_inst_dmem_U14158 ( .A1(MEM_stage_inst_dmem_ram_1840), .A2(MEM_stage_inst_dmem_n16412), .ZN(MEM_stage_inst_dmem_n16415) );
NAND2_X1 MEM_stage_inst_dmem_U14157 ( .A1(MEM_stage_inst_dmem_n16411), .A2(MEM_stage_inst_dmem_n16410), .ZN(MEM_stage_inst_dmem_n11116) );
NAND2_X1 MEM_stage_inst_dmem_U14156 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n16413), .ZN(MEM_stage_inst_dmem_n16410) );
NAND2_X1 MEM_stage_inst_dmem_U14155 ( .A1(MEM_stage_inst_dmem_ram_1841), .A2(MEM_stage_inst_dmem_n16412), .ZN(MEM_stage_inst_dmem_n16411) );
NAND2_X1 MEM_stage_inst_dmem_U14154 ( .A1(MEM_stage_inst_dmem_n16409), .A2(MEM_stage_inst_dmem_n16408), .ZN(MEM_stage_inst_dmem_n11117) );
NAND2_X1 MEM_stage_inst_dmem_U14153 ( .A1(MEM_stage_inst_dmem_n16789), .A2(MEM_stage_inst_dmem_n16413), .ZN(MEM_stage_inst_dmem_n16408) );
NAND2_X1 MEM_stage_inst_dmem_U14152 ( .A1(MEM_stage_inst_dmem_ram_1842), .A2(MEM_stage_inst_dmem_n16412), .ZN(MEM_stage_inst_dmem_n16409) );
NAND2_X1 MEM_stage_inst_dmem_U14151 ( .A1(MEM_stage_inst_dmem_n16407), .A2(MEM_stage_inst_dmem_n16406), .ZN(MEM_stage_inst_dmem_n11118) );
NAND2_X1 MEM_stage_inst_dmem_U14150 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n16413), .ZN(MEM_stage_inst_dmem_n16406) );
NAND2_X1 MEM_stage_inst_dmem_U14149 ( .A1(MEM_stage_inst_dmem_ram_1843), .A2(MEM_stage_inst_dmem_n16412), .ZN(MEM_stage_inst_dmem_n16407) );
NAND2_X1 MEM_stage_inst_dmem_U14148 ( .A1(MEM_stage_inst_dmem_n16405), .A2(MEM_stage_inst_dmem_n16404), .ZN(MEM_stage_inst_dmem_n11119) );
NAND2_X1 MEM_stage_inst_dmem_U14147 ( .A1(MEM_stage_inst_dmem_n16784), .A2(MEM_stage_inst_dmem_n16413), .ZN(MEM_stage_inst_dmem_n16404) );
NAND2_X1 MEM_stage_inst_dmem_U14146 ( .A1(MEM_stage_inst_dmem_ram_1844), .A2(MEM_stage_inst_dmem_n16412), .ZN(MEM_stage_inst_dmem_n16405) );
NAND2_X1 MEM_stage_inst_dmem_U14145 ( .A1(MEM_stage_inst_dmem_n16403), .A2(MEM_stage_inst_dmem_n16402), .ZN(MEM_stage_inst_dmem_n11120) );
NAND2_X1 MEM_stage_inst_dmem_U14144 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n16413), .ZN(MEM_stage_inst_dmem_n16402) );
NAND2_X1 MEM_stage_inst_dmem_U14143 ( .A1(MEM_stage_inst_dmem_ram_1845), .A2(MEM_stage_inst_dmem_n16412), .ZN(MEM_stage_inst_dmem_n16403) );
NAND2_X1 MEM_stage_inst_dmem_U14142 ( .A1(MEM_stage_inst_dmem_n16401), .A2(MEM_stage_inst_dmem_n16400), .ZN(MEM_stage_inst_dmem_n11121) );
NAND2_X1 MEM_stage_inst_dmem_U14141 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n16413), .ZN(MEM_stage_inst_dmem_n16400) );
NAND2_X1 MEM_stage_inst_dmem_U14140 ( .A1(MEM_stage_inst_dmem_ram_1846), .A2(MEM_stage_inst_dmem_n16412), .ZN(MEM_stage_inst_dmem_n16401) );
NAND2_X1 MEM_stage_inst_dmem_U14139 ( .A1(MEM_stage_inst_dmem_n16399), .A2(MEM_stage_inst_dmem_n16398), .ZN(MEM_stage_inst_dmem_n11122) );
NAND2_X1 MEM_stage_inst_dmem_U14138 ( .A1(MEM_stage_inst_dmem_n16777), .A2(MEM_stage_inst_dmem_n16413), .ZN(MEM_stage_inst_dmem_n16398) );
NAND2_X1 MEM_stage_inst_dmem_U14137 ( .A1(MEM_stage_inst_dmem_ram_1847), .A2(MEM_stage_inst_dmem_n16412), .ZN(MEM_stage_inst_dmem_n16399) );
NAND2_X1 MEM_stage_inst_dmem_U14136 ( .A1(MEM_stage_inst_dmem_n16397), .A2(MEM_stage_inst_dmem_n16396), .ZN(MEM_stage_inst_dmem_n11123) );
NAND2_X1 MEM_stage_inst_dmem_U14135 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n16413), .ZN(MEM_stage_inst_dmem_n16396) );
NAND2_X1 MEM_stage_inst_dmem_U14134 ( .A1(MEM_stage_inst_dmem_ram_1848), .A2(MEM_stage_inst_dmem_n16412), .ZN(MEM_stage_inst_dmem_n16397) );
NAND2_X1 MEM_stage_inst_dmem_U14133 ( .A1(MEM_stage_inst_dmem_n16395), .A2(MEM_stage_inst_dmem_n16394), .ZN(MEM_stage_inst_dmem_n11124) );
NAND2_X1 MEM_stage_inst_dmem_U14132 ( .A1(MEM_stage_inst_dmem_n16772), .A2(MEM_stage_inst_dmem_n16413), .ZN(MEM_stage_inst_dmem_n16394) );
NAND2_X1 MEM_stage_inst_dmem_U14131 ( .A1(MEM_stage_inst_dmem_ram_1849), .A2(MEM_stage_inst_dmem_n16412), .ZN(MEM_stage_inst_dmem_n16395) );
NAND2_X1 MEM_stage_inst_dmem_U14130 ( .A1(MEM_stage_inst_dmem_n16393), .A2(MEM_stage_inst_dmem_n16392), .ZN(MEM_stage_inst_dmem_n11125) );
NAND2_X1 MEM_stage_inst_dmem_U14129 ( .A1(MEM_stage_inst_dmem_n16769), .A2(MEM_stage_inst_dmem_n16413), .ZN(MEM_stage_inst_dmem_n16392) );
NAND2_X1 MEM_stage_inst_dmem_U14128 ( .A1(MEM_stage_inst_dmem_ram_1850), .A2(MEM_stage_inst_dmem_n16412), .ZN(MEM_stage_inst_dmem_n16393) );
NAND2_X1 MEM_stage_inst_dmem_U14127 ( .A1(MEM_stage_inst_dmem_n16391), .A2(MEM_stage_inst_dmem_n16390), .ZN(MEM_stage_inst_dmem_n11126) );
NAND2_X1 MEM_stage_inst_dmem_U14126 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n16413), .ZN(MEM_stage_inst_dmem_n16390) );
NAND2_X1 MEM_stage_inst_dmem_U14125 ( .A1(MEM_stage_inst_dmem_ram_1851), .A2(MEM_stage_inst_dmem_n16412), .ZN(MEM_stage_inst_dmem_n16391) );
NAND2_X1 MEM_stage_inst_dmem_U14124 ( .A1(MEM_stage_inst_dmem_n16389), .A2(MEM_stage_inst_dmem_n16388), .ZN(MEM_stage_inst_dmem_n11127) );
NAND2_X1 MEM_stage_inst_dmem_U14123 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n16413), .ZN(MEM_stage_inst_dmem_n16388) );
NAND2_X1 MEM_stage_inst_dmem_U14122 ( .A1(MEM_stage_inst_dmem_ram_1852), .A2(MEM_stage_inst_dmem_n16412), .ZN(MEM_stage_inst_dmem_n16389) );
NAND2_X1 MEM_stage_inst_dmem_U14121 ( .A1(MEM_stage_inst_dmem_n16387), .A2(MEM_stage_inst_dmem_n16386), .ZN(MEM_stage_inst_dmem_n11128) );
NAND2_X1 MEM_stage_inst_dmem_U14120 ( .A1(MEM_stage_inst_dmem_n15116), .A2(MEM_stage_inst_dmem_n16413), .ZN(MEM_stage_inst_dmem_n16386) );
NAND2_X1 MEM_stage_inst_dmem_U14119 ( .A1(MEM_stage_inst_dmem_ram_1853), .A2(MEM_stage_inst_dmem_n16412), .ZN(MEM_stage_inst_dmem_n16387) );
NAND2_X1 MEM_stage_inst_dmem_U14118 ( .A1(MEM_stage_inst_dmem_n16385), .A2(MEM_stage_inst_dmem_n16384), .ZN(MEM_stage_inst_dmem_n11129) );
NAND2_X1 MEM_stage_inst_dmem_U14117 ( .A1(MEM_stage_inst_dmem_n15113), .A2(MEM_stage_inst_dmem_n16413), .ZN(MEM_stage_inst_dmem_n16384) );
NAND2_X1 MEM_stage_inst_dmem_U14116 ( .A1(MEM_stage_inst_dmem_ram_1854), .A2(MEM_stage_inst_dmem_n16412), .ZN(MEM_stage_inst_dmem_n16385) );
NAND2_X1 MEM_stage_inst_dmem_U14115 ( .A1(MEM_stage_inst_dmem_n16383), .A2(MEM_stage_inst_dmem_n16382), .ZN(MEM_stage_inst_dmem_n11130) );
NAND2_X1 MEM_stage_inst_dmem_U14114 ( .A1(MEM_stage_inst_dmem_n16758), .A2(MEM_stage_inst_dmem_n16413), .ZN(MEM_stage_inst_dmem_n16382) );
INV_X1 MEM_stage_inst_dmem_U14113 ( .A(MEM_stage_inst_dmem_n16412), .ZN(MEM_stage_inst_dmem_n16413) );
NAND2_X1 MEM_stage_inst_dmem_U14112 ( .A1(MEM_stage_inst_dmem_ram_1855), .A2(MEM_stage_inst_dmem_n16412), .ZN(MEM_stage_inst_dmem_n16383) );
NAND2_X1 MEM_stage_inst_dmem_U14111 ( .A1(MEM_stage_inst_dmem_n21359), .A2(MEM_stage_inst_dmem_n16484), .ZN(MEM_stage_inst_dmem_n16412) );
NAND2_X1 MEM_stage_inst_dmem_U14110 ( .A1(MEM_stage_inst_dmem_n16381), .A2(MEM_stage_inst_dmem_n16380), .ZN(MEM_stage_inst_dmem_n11131) );
NAND2_X1 MEM_stage_inst_dmem_U14109 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n16379), .ZN(MEM_stage_inst_dmem_n16380) );
NAND2_X1 MEM_stage_inst_dmem_U14108 ( .A1(MEM_stage_inst_dmem_ram_1856), .A2(MEM_stage_inst_dmem_n16378), .ZN(MEM_stage_inst_dmem_n16381) );
NAND2_X1 MEM_stage_inst_dmem_U14107 ( .A1(MEM_stage_inst_dmem_n16377), .A2(MEM_stage_inst_dmem_n16376), .ZN(MEM_stage_inst_dmem_n11132) );
NAND2_X1 MEM_stage_inst_dmem_U14106 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n16379), .ZN(MEM_stage_inst_dmem_n16376) );
NAND2_X1 MEM_stage_inst_dmem_U14105 ( .A1(MEM_stage_inst_dmem_ram_1857), .A2(MEM_stage_inst_dmem_n16378), .ZN(MEM_stage_inst_dmem_n16377) );
NAND2_X1 MEM_stage_inst_dmem_U14104 ( .A1(MEM_stage_inst_dmem_n16375), .A2(MEM_stage_inst_dmem_n16374), .ZN(MEM_stage_inst_dmem_n11133) );
NAND2_X1 MEM_stage_inst_dmem_U14103 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n16379), .ZN(MEM_stage_inst_dmem_n16374) );
NAND2_X1 MEM_stage_inst_dmem_U14102 ( .A1(MEM_stage_inst_dmem_ram_1858), .A2(MEM_stage_inst_dmem_n16378), .ZN(MEM_stage_inst_dmem_n16375) );
NAND2_X1 MEM_stage_inst_dmem_U14101 ( .A1(MEM_stage_inst_dmem_n16372), .A2(MEM_stage_inst_dmem_n16371), .ZN(MEM_stage_inst_dmem_n11134) );
NAND2_X1 MEM_stage_inst_dmem_U14100 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n16379), .ZN(MEM_stage_inst_dmem_n16371) );
NAND2_X1 MEM_stage_inst_dmem_U14099 ( .A1(MEM_stage_inst_dmem_ram_1859), .A2(MEM_stage_inst_dmem_n16378), .ZN(MEM_stage_inst_dmem_n16372) );
NAND2_X1 MEM_stage_inst_dmem_U14098 ( .A1(MEM_stage_inst_dmem_n16370), .A2(MEM_stage_inst_dmem_n16369), .ZN(MEM_stage_inst_dmem_n11135) );
NAND2_X1 MEM_stage_inst_dmem_U14097 ( .A1(MEM_stage_inst_dmem_n16368), .A2(MEM_stage_inst_dmem_n16379), .ZN(MEM_stage_inst_dmem_n16369) );
NAND2_X1 MEM_stage_inst_dmem_U14096 ( .A1(MEM_stage_inst_dmem_ram_1860), .A2(MEM_stage_inst_dmem_n16378), .ZN(MEM_stage_inst_dmem_n16370) );
NAND2_X1 MEM_stage_inst_dmem_U14095 ( .A1(MEM_stage_inst_dmem_n16367), .A2(MEM_stage_inst_dmem_n16366), .ZN(MEM_stage_inst_dmem_n11136) );
NAND2_X1 MEM_stage_inst_dmem_U14094 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n16379), .ZN(MEM_stage_inst_dmem_n16366) );
NAND2_X1 MEM_stage_inst_dmem_U14093 ( .A1(MEM_stage_inst_dmem_ram_1861), .A2(MEM_stage_inst_dmem_n16378), .ZN(MEM_stage_inst_dmem_n16367) );
NAND2_X1 MEM_stage_inst_dmem_U14092 ( .A1(MEM_stage_inst_dmem_n16365), .A2(MEM_stage_inst_dmem_n16364), .ZN(MEM_stage_inst_dmem_n11137) );
NAND2_X1 MEM_stage_inst_dmem_U14091 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n16379), .ZN(MEM_stage_inst_dmem_n16364) );
NAND2_X1 MEM_stage_inst_dmem_U14090 ( .A1(MEM_stage_inst_dmem_ram_1862), .A2(MEM_stage_inst_dmem_n16378), .ZN(MEM_stage_inst_dmem_n16365) );
NAND2_X1 MEM_stage_inst_dmem_U14089 ( .A1(MEM_stage_inst_dmem_n16363), .A2(MEM_stage_inst_dmem_n16362), .ZN(MEM_stage_inst_dmem_n11138) );
NAND2_X1 MEM_stage_inst_dmem_U14088 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n16379), .ZN(MEM_stage_inst_dmem_n16362) );
NAND2_X1 MEM_stage_inst_dmem_U14087 ( .A1(MEM_stage_inst_dmem_ram_1863), .A2(MEM_stage_inst_dmem_n16378), .ZN(MEM_stage_inst_dmem_n16363) );
NAND2_X1 MEM_stage_inst_dmem_U14086 ( .A1(MEM_stage_inst_dmem_n16360), .A2(MEM_stage_inst_dmem_n16359), .ZN(MEM_stage_inst_dmem_n11139) );
NAND2_X1 MEM_stage_inst_dmem_U14085 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n16379), .ZN(MEM_stage_inst_dmem_n16359) );
NAND2_X1 MEM_stage_inst_dmem_U14084 ( .A1(MEM_stage_inst_dmem_ram_1864), .A2(MEM_stage_inst_dmem_n16378), .ZN(MEM_stage_inst_dmem_n16360) );
NAND2_X1 MEM_stage_inst_dmem_U14083 ( .A1(MEM_stage_inst_dmem_n16358), .A2(MEM_stage_inst_dmem_n16357), .ZN(MEM_stage_inst_dmem_n11140) );
NAND2_X1 MEM_stage_inst_dmem_U14082 ( .A1(MEM_stage_inst_dmem_n20524), .A2(MEM_stage_inst_dmem_n16379), .ZN(MEM_stage_inst_dmem_n16357) );
NAND2_X1 MEM_stage_inst_dmem_U14081 ( .A1(MEM_stage_inst_dmem_ram_1865), .A2(MEM_stage_inst_dmem_n16378), .ZN(MEM_stage_inst_dmem_n16358) );
NAND2_X1 MEM_stage_inst_dmem_U14080 ( .A1(MEM_stage_inst_dmem_n16356), .A2(MEM_stage_inst_dmem_n16355), .ZN(MEM_stage_inst_dmem_n11141) );
NAND2_X1 MEM_stage_inst_dmem_U14079 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n16379), .ZN(MEM_stage_inst_dmem_n16355) );
NAND2_X1 MEM_stage_inst_dmem_U14078 ( .A1(MEM_stage_inst_dmem_ram_1866), .A2(MEM_stage_inst_dmem_n16378), .ZN(MEM_stage_inst_dmem_n16356) );
NAND2_X1 MEM_stage_inst_dmem_U14077 ( .A1(MEM_stage_inst_dmem_n16353), .A2(MEM_stage_inst_dmem_n16352), .ZN(MEM_stage_inst_dmem_n11142) );
NAND2_X1 MEM_stage_inst_dmem_U14076 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n16379), .ZN(MEM_stage_inst_dmem_n16352) );
NAND2_X1 MEM_stage_inst_dmem_U14075 ( .A1(MEM_stage_inst_dmem_ram_1867), .A2(MEM_stage_inst_dmem_n16378), .ZN(MEM_stage_inst_dmem_n16353) );
NAND2_X1 MEM_stage_inst_dmem_U14074 ( .A1(MEM_stage_inst_dmem_n16351), .A2(MEM_stage_inst_dmem_n16350), .ZN(MEM_stage_inst_dmem_n11143) );
NAND2_X1 MEM_stage_inst_dmem_U14073 ( .A1(MEM_stage_inst_dmem_n18861), .A2(MEM_stage_inst_dmem_n16379), .ZN(MEM_stage_inst_dmem_n16350) );
NAND2_X1 MEM_stage_inst_dmem_U14072 ( .A1(MEM_stage_inst_dmem_ram_1868), .A2(MEM_stage_inst_dmem_n16378), .ZN(MEM_stage_inst_dmem_n16351) );
NAND2_X1 MEM_stage_inst_dmem_U14071 ( .A1(MEM_stage_inst_dmem_n16349), .A2(MEM_stage_inst_dmem_n16348), .ZN(MEM_stage_inst_dmem_n11144) );
NAND2_X1 MEM_stage_inst_dmem_U14070 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n16379), .ZN(MEM_stage_inst_dmem_n16348) );
NAND2_X1 MEM_stage_inst_dmem_U14069 ( .A1(MEM_stage_inst_dmem_ram_1869), .A2(MEM_stage_inst_dmem_n16378), .ZN(MEM_stage_inst_dmem_n16349) );
NAND2_X1 MEM_stage_inst_dmem_U14068 ( .A1(MEM_stage_inst_dmem_n16347), .A2(MEM_stage_inst_dmem_n16346), .ZN(MEM_stage_inst_dmem_n11145) );
NAND2_X1 MEM_stage_inst_dmem_U14067 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n16379), .ZN(MEM_stage_inst_dmem_n16346) );
NAND2_X1 MEM_stage_inst_dmem_U14066 ( .A1(MEM_stage_inst_dmem_ram_1870), .A2(MEM_stage_inst_dmem_n16378), .ZN(MEM_stage_inst_dmem_n16347) );
NAND2_X1 MEM_stage_inst_dmem_U14065 ( .A1(MEM_stage_inst_dmem_n16345), .A2(MEM_stage_inst_dmem_n16344), .ZN(MEM_stage_inst_dmem_n11146) );
NAND2_X1 MEM_stage_inst_dmem_U14064 ( .A1(MEM_stage_inst_dmem_n15110), .A2(MEM_stage_inst_dmem_n16379), .ZN(MEM_stage_inst_dmem_n16344) );
INV_X1 MEM_stage_inst_dmem_U14063 ( .A(MEM_stage_inst_dmem_n16378), .ZN(MEM_stage_inst_dmem_n16379) );
NAND2_X1 MEM_stage_inst_dmem_U14062 ( .A1(MEM_stage_inst_dmem_ram_1871), .A2(MEM_stage_inst_dmem_n16378), .ZN(MEM_stage_inst_dmem_n16345) );
NAND2_X1 MEM_stage_inst_dmem_U14061 ( .A1(MEM_stage_inst_dmem_n21319), .A2(MEM_stage_inst_dmem_n16484), .ZN(MEM_stage_inst_dmem_n16378) );
NAND2_X1 MEM_stage_inst_dmem_U14060 ( .A1(MEM_stage_inst_dmem_n16342), .A2(MEM_stage_inst_dmem_n16341), .ZN(MEM_stage_inst_dmem_n11147) );
NAND2_X1 MEM_stage_inst_dmem_U14059 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n16340), .ZN(MEM_stage_inst_dmem_n16341) );
NAND2_X1 MEM_stage_inst_dmem_U14058 ( .A1(MEM_stage_inst_dmem_ram_1872), .A2(MEM_stage_inst_dmem_n16339), .ZN(MEM_stage_inst_dmem_n16342) );
NAND2_X1 MEM_stage_inst_dmem_U14057 ( .A1(MEM_stage_inst_dmem_n16338), .A2(MEM_stage_inst_dmem_n16337), .ZN(MEM_stage_inst_dmem_n11148) );
NAND2_X1 MEM_stage_inst_dmem_U14056 ( .A1(MEM_stage_inst_dmem_n109), .A2(MEM_stage_inst_dmem_n16340), .ZN(MEM_stage_inst_dmem_n16337) );
NAND2_X1 MEM_stage_inst_dmem_U14055 ( .A1(MEM_stage_inst_dmem_ram_1873), .A2(MEM_stage_inst_dmem_n16339), .ZN(MEM_stage_inst_dmem_n16338) );
NAND2_X1 MEM_stage_inst_dmem_U14054 ( .A1(MEM_stage_inst_dmem_n16336), .A2(MEM_stage_inst_dmem_n16335), .ZN(MEM_stage_inst_dmem_n11149) );
NAND2_X1 MEM_stage_inst_dmem_U14053 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n16340), .ZN(MEM_stage_inst_dmem_n16335) );
NAND2_X1 MEM_stage_inst_dmem_U14052 ( .A1(MEM_stage_inst_dmem_ram_1874), .A2(MEM_stage_inst_dmem_n16339), .ZN(MEM_stage_inst_dmem_n16336) );
NAND2_X1 MEM_stage_inst_dmem_U14051 ( .A1(MEM_stage_inst_dmem_n16334), .A2(MEM_stage_inst_dmem_n16333), .ZN(MEM_stage_inst_dmem_n11150) );
NAND2_X1 MEM_stage_inst_dmem_U14050 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n16340), .ZN(MEM_stage_inst_dmem_n16333) );
NAND2_X1 MEM_stage_inst_dmem_U14049 ( .A1(MEM_stage_inst_dmem_ram_1875), .A2(MEM_stage_inst_dmem_n16339), .ZN(MEM_stage_inst_dmem_n16334) );
NAND2_X1 MEM_stage_inst_dmem_U14048 ( .A1(MEM_stage_inst_dmem_n16332), .A2(MEM_stage_inst_dmem_n16331), .ZN(MEM_stage_inst_dmem_n11151) );
NAND2_X1 MEM_stage_inst_dmem_U14047 ( .A1(MEM_stage_inst_dmem_n16368), .A2(MEM_stage_inst_dmem_n16340), .ZN(MEM_stage_inst_dmem_n16331) );
NAND2_X1 MEM_stage_inst_dmem_U14046 ( .A1(MEM_stage_inst_dmem_ram_1876), .A2(MEM_stage_inst_dmem_n16339), .ZN(MEM_stage_inst_dmem_n16332) );
NAND2_X1 MEM_stage_inst_dmem_U14045 ( .A1(MEM_stage_inst_dmem_n16330), .A2(MEM_stage_inst_dmem_n16329), .ZN(MEM_stage_inst_dmem_n11152) );
NAND2_X1 MEM_stage_inst_dmem_U14044 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n16340), .ZN(MEM_stage_inst_dmem_n16329) );
NAND2_X1 MEM_stage_inst_dmem_U14043 ( .A1(MEM_stage_inst_dmem_ram_1877), .A2(MEM_stage_inst_dmem_n16339), .ZN(MEM_stage_inst_dmem_n16330) );
NAND2_X1 MEM_stage_inst_dmem_U14042 ( .A1(MEM_stage_inst_dmem_n16328), .A2(MEM_stage_inst_dmem_n16327), .ZN(MEM_stage_inst_dmem_n11153) );
NAND2_X1 MEM_stage_inst_dmem_U14041 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n16340), .ZN(MEM_stage_inst_dmem_n16327) );
NAND2_X1 MEM_stage_inst_dmem_U14040 ( .A1(MEM_stage_inst_dmem_ram_1878), .A2(MEM_stage_inst_dmem_n16339), .ZN(MEM_stage_inst_dmem_n16328) );
NAND2_X1 MEM_stage_inst_dmem_U14039 ( .A1(MEM_stage_inst_dmem_n16326), .A2(MEM_stage_inst_dmem_n16325), .ZN(MEM_stage_inst_dmem_n11154) );
NAND2_X1 MEM_stage_inst_dmem_U14038 ( .A1(MEM_stage_inst_dmem_n112), .A2(MEM_stage_inst_dmem_n16340), .ZN(MEM_stage_inst_dmem_n16325) );
NAND2_X1 MEM_stage_inst_dmem_U14037 ( .A1(MEM_stage_inst_dmem_ram_1879), .A2(MEM_stage_inst_dmem_n16339), .ZN(MEM_stage_inst_dmem_n16326) );
NAND2_X1 MEM_stage_inst_dmem_U14036 ( .A1(MEM_stage_inst_dmem_n16324), .A2(MEM_stage_inst_dmem_n16323), .ZN(MEM_stage_inst_dmem_n11155) );
NAND2_X1 MEM_stage_inst_dmem_U14035 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n16340), .ZN(MEM_stage_inst_dmem_n16323) );
NAND2_X1 MEM_stage_inst_dmem_U14034 ( .A1(MEM_stage_inst_dmem_ram_1880), .A2(MEM_stage_inst_dmem_n16339), .ZN(MEM_stage_inst_dmem_n16324) );
NAND2_X1 MEM_stage_inst_dmem_U14033 ( .A1(MEM_stage_inst_dmem_n16322), .A2(MEM_stage_inst_dmem_n16321), .ZN(MEM_stage_inst_dmem_n11156) );
NAND2_X1 MEM_stage_inst_dmem_U14032 ( .A1(EX_pipeline_reg_out_14), .A2(MEM_stage_inst_dmem_n16340), .ZN(MEM_stage_inst_dmem_n16321) );
NAND2_X1 MEM_stage_inst_dmem_U14031 ( .A1(MEM_stage_inst_dmem_ram_1881), .A2(MEM_stage_inst_dmem_n16339), .ZN(MEM_stage_inst_dmem_n16322) );
NAND2_X1 MEM_stage_inst_dmem_U14030 ( .A1(MEM_stage_inst_dmem_n16320), .A2(MEM_stage_inst_dmem_n16319), .ZN(MEM_stage_inst_dmem_n11157) );
NAND2_X1 MEM_stage_inst_dmem_U14029 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n16340), .ZN(MEM_stage_inst_dmem_n16319) );
NAND2_X1 MEM_stage_inst_dmem_U14028 ( .A1(MEM_stage_inst_dmem_ram_1882), .A2(MEM_stage_inst_dmem_n16339), .ZN(MEM_stage_inst_dmem_n16320) );
NAND2_X1 MEM_stage_inst_dmem_U14027 ( .A1(MEM_stage_inst_dmem_n16318), .A2(MEM_stage_inst_dmem_n16317), .ZN(MEM_stage_inst_dmem_n11158) );
NAND2_X1 MEM_stage_inst_dmem_U14026 ( .A1(MEM_stage_inst_dmem_n18864), .A2(MEM_stage_inst_dmem_n16340), .ZN(MEM_stage_inst_dmem_n16317) );
NAND2_X1 MEM_stage_inst_dmem_U14025 ( .A1(MEM_stage_inst_dmem_ram_1883), .A2(MEM_stage_inst_dmem_n16339), .ZN(MEM_stage_inst_dmem_n16318) );
NAND2_X1 MEM_stage_inst_dmem_U14024 ( .A1(MEM_stage_inst_dmem_n16316), .A2(MEM_stage_inst_dmem_n16315), .ZN(MEM_stage_inst_dmem_n11159) );
NAND2_X1 MEM_stage_inst_dmem_U14023 ( .A1(EX_pipeline_reg_out_17), .A2(MEM_stage_inst_dmem_n16340), .ZN(MEM_stage_inst_dmem_n16315) );
NAND2_X1 MEM_stage_inst_dmem_U14022 ( .A1(MEM_stage_inst_dmem_ram_1884), .A2(MEM_stage_inst_dmem_n16339), .ZN(MEM_stage_inst_dmem_n16316) );
NAND2_X1 MEM_stage_inst_dmem_U14021 ( .A1(MEM_stage_inst_dmem_n16314), .A2(MEM_stage_inst_dmem_n16313), .ZN(MEM_stage_inst_dmem_n11160) );
NAND2_X1 MEM_stage_inst_dmem_U14020 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n16340), .ZN(MEM_stage_inst_dmem_n16313) );
NAND2_X1 MEM_stage_inst_dmem_U14019 ( .A1(MEM_stage_inst_dmem_ram_1885), .A2(MEM_stage_inst_dmem_n16339), .ZN(MEM_stage_inst_dmem_n16314) );
NAND2_X1 MEM_stage_inst_dmem_U14018 ( .A1(MEM_stage_inst_dmem_n16312), .A2(MEM_stage_inst_dmem_n16311), .ZN(MEM_stage_inst_dmem_n11161) );
NAND2_X1 MEM_stage_inst_dmem_U14017 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n16340), .ZN(MEM_stage_inst_dmem_n16311) );
NAND2_X1 MEM_stage_inst_dmem_U14016 ( .A1(MEM_stage_inst_dmem_ram_1886), .A2(MEM_stage_inst_dmem_n16339), .ZN(MEM_stage_inst_dmem_n16312) );
NAND2_X1 MEM_stage_inst_dmem_U14015 ( .A1(MEM_stage_inst_dmem_n16310), .A2(MEM_stage_inst_dmem_n16309), .ZN(MEM_stage_inst_dmem_n11162) );
NAND2_X1 MEM_stage_inst_dmem_U14014 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n16340), .ZN(MEM_stage_inst_dmem_n16309) );
NAND2_X1 MEM_stage_inst_dmem_U14013 ( .A1(MEM_stage_inst_dmem_ram_1887), .A2(MEM_stage_inst_dmem_n16339), .ZN(MEM_stage_inst_dmem_n16310) );
NAND2_X1 MEM_stage_inst_dmem_U14012 ( .A1(MEM_stage_inst_dmem_n21284), .A2(MEM_stage_inst_dmem_n16484), .ZN(MEM_stage_inst_dmem_n16339) );
NAND2_X1 MEM_stage_inst_dmem_U14011 ( .A1(MEM_stage_inst_dmem_n16308), .A2(MEM_stage_inst_dmem_n16307), .ZN(MEM_stage_inst_dmem_n11163) );
NAND2_X1 MEM_stage_inst_dmem_U14010 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n16306), .ZN(MEM_stage_inst_dmem_n16307) );
NAND2_X1 MEM_stage_inst_dmem_U14009 ( .A1(MEM_stage_inst_dmem_ram_1888), .A2(MEM_stage_inst_dmem_n16305), .ZN(MEM_stage_inst_dmem_n16308) );
NAND2_X1 MEM_stage_inst_dmem_U14008 ( .A1(MEM_stage_inst_dmem_n16304), .A2(MEM_stage_inst_dmem_n16303), .ZN(MEM_stage_inst_dmem_n11164) );
NAND2_X1 MEM_stage_inst_dmem_U14007 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n16306), .ZN(MEM_stage_inst_dmem_n16303) );
NAND2_X1 MEM_stage_inst_dmem_U14006 ( .A1(MEM_stage_inst_dmem_ram_1889), .A2(MEM_stage_inst_dmem_n16305), .ZN(MEM_stage_inst_dmem_n16304) );
NAND2_X1 MEM_stage_inst_dmem_U14005 ( .A1(MEM_stage_inst_dmem_n16302), .A2(MEM_stage_inst_dmem_n16301), .ZN(MEM_stage_inst_dmem_n11165) );
NAND2_X1 MEM_stage_inst_dmem_U14004 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n16306), .ZN(MEM_stage_inst_dmem_n16301) );
NAND2_X1 MEM_stage_inst_dmem_U14003 ( .A1(MEM_stage_inst_dmem_ram_1890), .A2(MEM_stage_inst_dmem_n16305), .ZN(MEM_stage_inst_dmem_n16302) );
NAND2_X1 MEM_stage_inst_dmem_U14002 ( .A1(MEM_stage_inst_dmem_n16300), .A2(MEM_stage_inst_dmem_n16299), .ZN(MEM_stage_inst_dmem_n11166) );
NAND2_X1 MEM_stage_inst_dmem_U14001 ( .A1(MEM_stage_inst_dmem_n13064), .A2(MEM_stage_inst_dmem_n16306), .ZN(MEM_stage_inst_dmem_n16299) );
NAND2_X1 MEM_stage_inst_dmem_U14000 ( .A1(MEM_stage_inst_dmem_ram_1891), .A2(MEM_stage_inst_dmem_n16305), .ZN(MEM_stage_inst_dmem_n16300) );
NAND2_X1 MEM_stage_inst_dmem_U13999 ( .A1(MEM_stage_inst_dmem_n16298), .A2(MEM_stage_inst_dmem_n16297), .ZN(MEM_stage_inst_dmem_n11167) );
NAND2_X1 MEM_stage_inst_dmem_U13998 ( .A1(MEM_stage_inst_dmem_n16368), .A2(MEM_stage_inst_dmem_n16306), .ZN(MEM_stage_inst_dmem_n16297) );
NAND2_X1 MEM_stage_inst_dmem_U13997 ( .A1(MEM_stage_inst_dmem_ram_1892), .A2(MEM_stage_inst_dmem_n16305), .ZN(MEM_stage_inst_dmem_n16298) );
NAND2_X1 MEM_stage_inst_dmem_U13996 ( .A1(MEM_stage_inst_dmem_n16296), .A2(MEM_stage_inst_dmem_n16295), .ZN(MEM_stage_inst_dmem_n11168) );
NAND2_X1 MEM_stage_inst_dmem_U13995 ( .A1(MEM_stage_inst_dmem_n13059), .A2(MEM_stage_inst_dmem_n16306), .ZN(MEM_stage_inst_dmem_n16295) );
NAND2_X1 MEM_stage_inst_dmem_U13994 ( .A1(MEM_stage_inst_dmem_ram_1893), .A2(MEM_stage_inst_dmem_n16305), .ZN(MEM_stage_inst_dmem_n16296) );
NAND2_X1 MEM_stage_inst_dmem_U13993 ( .A1(MEM_stage_inst_dmem_n16294), .A2(MEM_stage_inst_dmem_n16293), .ZN(MEM_stage_inst_dmem_n11169) );
NAND2_X1 MEM_stage_inst_dmem_U13992 ( .A1(MEM_stage_inst_dmem_n13056), .A2(MEM_stage_inst_dmem_n16306), .ZN(MEM_stage_inst_dmem_n16293) );
NAND2_X1 MEM_stage_inst_dmem_U13991 ( .A1(MEM_stage_inst_dmem_ram_1894), .A2(MEM_stage_inst_dmem_n16305), .ZN(MEM_stage_inst_dmem_n16294) );
NAND2_X1 MEM_stage_inst_dmem_U13990 ( .A1(MEM_stage_inst_dmem_n16292), .A2(MEM_stage_inst_dmem_n16291), .ZN(MEM_stage_inst_dmem_n11170) );
NAND2_X1 MEM_stage_inst_dmem_U13989 ( .A1(MEM_stage_inst_dmem_n16361), .A2(MEM_stage_inst_dmem_n16306), .ZN(MEM_stage_inst_dmem_n16291) );
NAND2_X1 MEM_stage_inst_dmem_U13988 ( .A1(MEM_stage_inst_dmem_ram_1895), .A2(MEM_stage_inst_dmem_n16305), .ZN(MEM_stage_inst_dmem_n16292) );
NAND2_X1 MEM_stage_inst_dmem_U13987 ( .A1(MEM_stage_inst_dmem_n16290), .A2(MEM_stage_inst_dmem_n16289), .ZN(MEM_stage_inst_dmem_n11171) );
NAND2_X1 MEM_stage_inst_dmem_U13986 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n16306), .ZN(MEM_stage_inst_dmem_n16289) );
NAND2_X1 MEM_stage_inst_dmem_U13985 ( .A1(MEM_stage_inst_dmem_ram_1896), .A2(MEM_stage_inst_dmem_n16305), .ZN(MEM_stage_inst_dmem_n16290) );
NAND2_X1 MEM_stage_inst_dmem_U13984 ( .A1(MEM_stage_inst_dmem_n16288), .A2(MEM_stage_inst_dmem_n16287), .ZN(MEM_stage_inst_dmem_n11172) );
NAND2_X1 MEM_stage_inst_dmem_U13983 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n16306), .ZN(MEM_stage_inst_dmem_n16287) );
NAND2_X1 MEM_stage_inst_dmem_U13982 ( .A1(MEM_stage_inst_dmem_ram_1897), .A2(MEM_stage_inst_dmem_n16305), .ZN(MEM_stage_inst_dmem_n16288) );
NAND2_X1 MEM_stage_inst_dmem_U13981 ( .A1(MEM_stage_inst_dmem_n16286), .A2(MEM_stage_inst_dmem_n16285), .ZN(MEM_stage_inst_dmem_n11173) );
NAND2_X1 MEM_stage_inst_dmem_U13980 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n16306), .ZN(MEM_stage_inst_dmem_n16285) );
NAND2_X1 MEM_stage_inst_dmem_U13979 ( .A1(MEM_stage_inst_dmem_ram_1898), .A2(MEM_stage_inst_dmem_n16305), .ZN(MEM_stage_inst_dmem_n16286) );
NAND2_X1 MEM_stage_inst_dmem_U13978 ( .A1(MEM_stage_inst_dmem_n16284), .A2(MEM_stage_inst_dmem_n16283), .ZN(MEM_stage_inst_dmem_n11174) );
NAND2_X1 MEM_stage_inst_dmem_U13977 ( .A1(EX_pipeline_reg_out_16), .A2(MEM_stage_inst_dmem_n16306), .ZN(MEM_stage_inst_dmem_n16283) );
NAND2_X1 MEM_stage_inst_dmem_U13976 ( .A1(MEM_stage_inst_dmem_ram_1899), .A2(MEM_stage_inst_dmem_n16305), .ZN(MEM_stage_inst_dmem_n16284) );
NAND2_X1 MEM_stage_inst_dmem_U13975 ( .A1(MEM_stage_inst_dmem_n16282), .A2(MEM_stage_inst_dmem_n16281), .ZN(MEM_stage_inst_dmem_n11175) );
NAND2_X1 MEM_stage_inst_dmem_U13974 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n16306), .ZN(MEM_stage_inst_dmem_n16281) );
NAND2_X1 MEM_stage_inst_dmem_U13973 ( .A1(MEM_stage_inst_dmem_ram_1900), .A2(MEM_stage_inst_dmem_n16305), .ZN(MEM_stage_inst_dmem_n16282) );
NAND2_X1 MEM_stage_inst_dmem_U13972 ( .A1(MEM_stage_inst_dmem_n16280), .A2(MEM_stage_inst_dmem_n16279), .ZN(MEM_stage_inst_dmem_n11176) );
NAND2_X1 MEM_stage_inst_dmem_U13971 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n16306), .ZN(MEM_stage_inst_dmem_n16279) );
NAND2_X1 MEM_stage_inst_dmem_U13970 ( .A1(MEM_stage_inst_dmem_ram_1901), .A2(MEM_stage_inst_dmem_n16305), .ZN(MEM_stage_inst_dmem_n16280) );
NAND2_X1 MEM_stage_inst_dmem_U13969 ( .A1(MEM_stage_inst_dmem_n16278), .A2(MEM_stage_inst_dmem_n16277), .ZN(MEM_stage_inst_dmem_n11177) );
NAND2_X1 MEM_stage_inst_dmem_U13968 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n16306), .ZN(MEM_stage_inst_dmem_n16277) );
NAND2_X1 MEM_stage_inst_dmem_U13967 ( .A1(MEM_stage_inst_dmem_ram_1902), .A2(MEM_stage_inst_dmem_n16305), .ZN(MEM_stage_inst_dmem_n16278) );
NAND2_X1 MEM_stage_inst_dmem_U13966 ( .A1(MEM_stage_inst_dmem_n16276), .A2(MEM_stage_inst_dmem_n16275), .ZN(MEM_stage_inst_dmem_n11178) );
NAND2_X1 MEM_stage_inst_dmem_U13965 ( .A1(MEM_stage_inst_dmem_n16343), .A2(MEM_stage_inst_dmem_n16306), .ZN(MEM_stage_inst_dmem_n16275) );
INV_X1 MEM_stage_inst_dmem_U13964 ( .A(MEM_stage_inst_dmem_n16305), .ZN(MEM_stage_inst_dmem_n16306) );
NAND2_X1 MEM_stage_inst_dmem_U13963 ( .A1(MEM_stage_inst_dmem_ram_1903), .A2(MEM_stage_inst_dmem_n16305), .ZN(MEM_stage_inst_dmem_n16276) );
NAND2_X1 MEM_stage_inst_dmem_U13962 ( .A1(MEM_stage_inst_dmem_n21249), .A2(MEM_stage_inst_dmem_n16484), .ZN(MEM_stage_inst_dmem_n16305) );
NAND2_X1 MEM_stage_inst_dmem_U13961 ( .A1(MEM_stage_inst_dmem_n16274), .A2(MEM_stage_inst_dmem_n16273), .ZN(MEM_stage_inst_dmem_n11179) );
NAND2_X1 MEM_stage_inst_dmem_U13960 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n16272), .ZN(MEM_stage_inst_dmem_n16273) );
NAND2_X1 MEM_stage_inst_dmem_U13959 ( .A1(MEM_stage_inst_dmem_ram_1904), .A2(MEM_stage_inst_dmem_n16271), .ZN(MEM_stage_inst_dmem_n16274) );
NAND2_X1 MEM_stage_inst_dmem_U13958 ( .A1(MEM_stage_inst_dmem_n16270), .A2(MEM_stage_inst_dmem_n16269), .ZN(MEM_stage_inst_dmem_n11180) );
NAND2_X1 MEM_stage_inst_dmem_U13957 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n16272), .ZN(MEM_stage_inst_dmem_n16269) );
NAND2_X1 MEM_stage_inst_dmem_U13956 ( .A1(MEM_stage_inst_dmem_ram_1905), .A2(MEM_stage_inst_dmem_n16271), .ZN(MEM_stage_inst_dmem_n16270) );
NAND2_X1 MEM_stage_inst_dmem_U13955 ( .A1(MEM_stage_inst_dmem_n16268), .A2(MEM_stage_inst_dmem_n16267), .ZN(MEM_stage_inst_dmem_n11181) );
NAND2_X1 MEM_stage_inst_dmem_U13954 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n16272), .ZN(MEM_stage_inst_dmem_n16267) );
NAND2_X1 MEM_stage_inst_dmem_U13953 ( .A1(MEM_stage_inst_dmem_ram_1906), .A2(MEM_stage_inst_dmem_n16271), .ZN(MEM_stage_inst_dmem_n16268) );
NAND2_X1 MEM_stage_inst_dmem_U13952 ( .A1(MEM_stage_inst_dmem_n16266), .A2(MEM_stage_inst_dmem_n16265), .ZN(MEM_stage_inst_dmem_n11182) );
NAND2_X1 MEM_stage_inst_dmem_U13951 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n16272), .ZN(MEM_stage_inst_dmem_n16265) );
NAND2_X1 MEM_stage_inst_dmem_U13950 ( .A1(MEM_stage_inst_dmem_ram_1907), .A2(MEM_stage_inst_dmem_n16271), .ZN(MEM_stage_inst_dmem_n16266) );
NAND2_X1 MEM_stage_inst_dmem_U13949 ( .A1(MEM_stage_inst_dmem_n16264), .A2(MEM_stage_inst_dmem_n16263), .ZN(MEM_stage_inst_dmem_n11183) );
NAND2_X1 MEM_stage_inst_dmem_U13948 ( .A1(MEM_stage_inst_dmem_n16368), .A2(MEM_stage_inst_dmem_n16272), .ZN(MEM_stage_inst_dmem_n16263) );
NAND2_X1 MEM_stage_inst_dmem_U13947 ( .A1(MEM_stage_inst_dmem_ram_1908), .A2(MEM_stage_inst_dmem_n16271), .ZN(MEM_stage_inst_dmem_n16264) );
NAND2_X1 MEM_stage_inst_dmem_U13946 ( .A1(MEM_stage_inst_dmem_n16262), .A2(MEM_stage_inst_dmem_n16261), .ZN(MEM_stage_inst_dmem_n11184) );
NAND2_X1 MEM_stage_inst_dmem_U13945 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n16272), .ZN(MEM_stage_inst_dmem_n16261) );
NAND2_X1 MEM_stage_inst_dmem_U13944 ( .A1(MEM_stage_inst_dmem_ram_1909), .A2(MEM_stage_inst_dmem_n16271), .ZN(MEM_stage_inst_dmem_n16262) );
NAND2_X1 MEM_stage_inst_dmem_U13943 ( .A1(MEM_stage_inst_dmem_n16260), .A2(MEM_stage_inst_dmem_n16259), .ZN(MEM_stage_inst_dmem_n11185) );
NAND2_X1 MEM_stage_inst_dmem_U13942 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n16272), .ZN(MEM_stage_inst_dmem_n16259) );
NAND2_X1 MEM_stage_inst_dmem_U13941 ( .A1(MEM_stage_inst_dmem_ram_1910), .A2(MEM_stage_inst_dmem_n16271), .ZN(MEM_stage_inst_dmem_n16260) );
NAND2_X1 MEM_stage_inst_dmem_U13940 ( .A1(MEM_stage_inst_dmem_n16258), .A2(MEM_stage_inst_dmem_n16257), .ZN(MEM_stage_inst_dmem_n11186) );
NAND2_X1 MEM_stage_inst_dmem_U13939 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n16272), .ZN(MEM_stage_inst_dmem_n16257) );
NAND2_X1 MEM_stage_inst_dmem_U13938 ( .A1(MEM_stage_inst_dmem_ram_1911), .A2(MEM_stage_inst_dmem_n16271), .ZN(MEM_stage_inst_dmem_n16258) );
NAND2_X1 MEM_stage_inst_dmem_U13937 ( .A1(MEM_stage_inst_dmem_n16256), .A2(MEM_stage_inst_dmem_n16255), .ZN(MEM_stage_inst_dmem_n11187) );
NAND2_X1 MEM_stage_inst_dmem_U13936 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n16272), .ZN(MEM_stage_inst_dmem_n16255) );
NAND2_X1 MEM_stage_inst_dmem_U13935 ( .A1(MEM_stage_inst_dmem_ram_1912), .A2(MEM_stage_inst_dmem_n16271), .ZN(MEM_stage_inst_dmem_n16256) );
NAND2_X1 MEM_stage_inst_dmem_U13934 ( .A1(MEM_stage_inst_dmem_n16254), .A2(MEM_stage_inst_dmem_n16253), .ZN(MEM_stage_inst_dmem_n11188) );
NAND2_X1 MEM_stage_inst_dmem_U13933 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n16272), .ZN(MEM_stage_inst_dmem_n16253) );
NAND2_X1 MEM_stage_inst_dmem_U13932 ( .A1(MEM_stage_inst_dmem_ram_1913), .A2(MEM_stage_inst_dmem_n16271), .ZN(MEM_stage_inst_dmem_n16254) );
NAND2_X1 MEM_stage_inst_dmem_U13931 ( .A1(MEM_stage_inst_dmem_n16252), .A2(MEM_stage_inst_dmem_n16251), .ZN(MEM_stage_inst_dmem_n11189) );
NAND2_X1 MEM_stage_inst_dmem_U13930 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n16272), .ZN(MEM_stage_inst_dmem_n16251) );
NAND2_X1 MEM_stage_inst_dmem_U13929 ( .A1(MEM_stage_inst_dmem_ram_1914), .A2(MEM_stage_inst_dmem_n16271), .ZN(MEM_stage_inst_dmem_n16252) );
NAND2_X1 MEM_stage_inst_dmem_U13928 ( .A1(MEM_stage_inst_dmem_n16250), .A2(MEM_stage_inst_dmem_n16249), .ZN(MEM_stage_inst_dmem_n11190) );
NAND2_X1 MEM_stage_inst_dmem_U13927 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n16272), .ZN(MEM_stage_inst_dmem_n16249) );
NAND2_X1 MEM_stage_inst_dmem_U13926 ( .A1(MEM_stage_inst_dmem_ram_1915), .A2(MEM_stage_inst_dmem_n16271), .ZN(MEM_stage_inst_dmem_n16250) );
NAND2_X1 MEM_stage_inst_dmem_U13925 ( .A1(MEM_stage_inst_dmem_n16248), .A2(MEM_stage_inst_dmem_n16247), .ZN(MEM_stage_inst_dmem_n11191) );
NAND2_X1 MEM_stage_inst_dmem_U13924 ( .A1(MEM_stage_inst_dmem_n13041), .A2(MEM_stage_inst_dmem_n16272), .ZN(MEM_stage_inst_dmem_n16247) );
NAND2_X1 MEM_stage_inst_dmem_U13923 ( .A1(MEM_stage_inst_dmem_ram_1916), .A2(MEM_stage_inst_dmem_n16271), .ZN(MEM_stage_inst_dmem_n16248) );
NAND2_X1 MEM_stage_inst_dmem_U13922 ( .A1(MEM_stage_inst_dmem_n16246), .A2(MEM_stage_inst_dmem_n16245), .ZN(MEM_stage_inst_dmem_n11192) );
NAND2_X1 MEM_stage_inst_dmem_U13921 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n16272), .ZN(MEM_stage_inst_dmem_n16245) );
NAND2_X1 MEM_stage_inst_dmem_U13920 ( .A1(MEM_stage_inst_dmem_ram_1917), .A2(MEM_stage_inst_dmem_n16271), .ZN(MEM_stage_inst_dmem_n16246) );
NAND2_X1 MEM_stage_inst_dmem_U13919 ( .A1(MEM_stage_inst_dmem_n16244), .A2(MEM_stage_inst_dmem_n16243), .ZN(MEM_stage_inst_dmem_n11193) );
NAND2_X1 MEM_stage_inst_dmem_U13918 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n16272), .ZN(MEM_stage_inst_dmem_n16243) );
NAND2_X1 MEM_stage_inst_dmem_U13917 ( .A1(MEM_stage_inst_dmem_ram_1918), .A2(MEM_stage_inst_dmem_n16271), .ZN(MEM_stage_inst_dmem_n16244) );
NAND2_X1 MEM_stage_inst_dmem_U13916 ( .A1(MEM_stage_inst_dmem_n16242), .A2(MEM_stage_inst_dmem_n16241), .ZN(MEM_stage_inst_dmem_n11194) );
NAND2_X1 MEM_stage_inst_dmem_U13915 ( .A1(MEM_stage_inst_dmem_n14693), .A2(MEM_stage_inst_dmem_n16272), .ZN(MEM_stage_inst_dmem_n16241) );
INV_X1 MEM_stage_inst_dmem_U13914 ( .A(MEM_stage_inst_dmem_n16271), .ZN(MEM_stage_inst_dmem_n16272) );
NAND2_X1 MEM_stage_inst_dmem_U13913 ( .A1(MEM_stage_inst_dmem_ram_1919), .A2(MEM_stage_inst_dmem_n16271), .ZN(MEM_stage_inst_dmem_n16242) );
NAND2_X1 MEM_stage_inst_dmem_U13912 ( .A1(MEM_stage_inst_dmem_n21214), .A2(MEM_stage_inst_dmem_n16484), .ZN(MEM_stage_inst_dmem_n16271) );
NAND2_X1 MEM_stage_inst_dmem_U13911 ( .A1(MEM_stage_inst_dmem_n16240), .A2(MEM_stage_inst_dmem_n16239), .ZN(MEM_stage_inst_dmem_n11195) );
NAND2_X1 MEM_stage_inst_dmem_U13910 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n16238), .ZN(MEM_stage_inst_dmem_n16239) );
NAND2_X1 MEM_stage_inst_dmem_U13909 ( .A1(MEM_stage_inst_dmem_ram_1920), .A2(MEM_stage_inst_dmem_n16237), .ZN(MEM_stage_inst_dmem_n16240) );
NAND2_X1 MEM_stage_inst_dmem_U13908 ( .A1(MEM_stage_inst_dmem_n16236), .A2(MEM_stage_inst_dmem_n16235), .ZN(MEM_stage_inst_dmem_n11196) );
NAND2_X1 MEM_stage_inst_dmem_U13907 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n16238), .ZN(MEM_stage_inst_dmem_n16235) );
NAND2_X1 MEM_stage_inst_dmem_U13906 ( .A1(MEM_stage_inst_dmem_ram_1921), .A2(MEM_stage_inst_dmem_n16237), .ZN(MEM_stage_inst_dmem_n16236) );
NAND2_X1 MEM_stage_inst_dmem_U13905 ( .A1(MEM_stage_inst_dmem_n16234), .A2(MEM_stage_inst_dmem_n16233), .ZN(MEM_stage_inst_dmem_n11197) );
NAND2_X1 MEM_stage_inst_dmem_U13904 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n16238), .ZN(MEM_stage_inst_dmem_n16233) );
NAND2_X1 MEM_stage_inst_dmem_U13903 ( .A1(MEM_stage_inst_dmem_ram_1922), .A2(MEM_stage_inst_dmem_n16237), .ZN(MEM_stage_inst_dmem_n16234) );
NAND2_X1 MEM_stage_inst_dmem_U13902 ( .A1(MEM_stage_inst_dmem_n16232), .A2(MEM_stage_inst_dmem_n16231), .ZN(MEM_stage_inst_dmem_n11198) );
NAND2_X1 MEM_stage_inst_dmem_U13901 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n16238), .ZN(MEM_stage_inst_dmem_n16231) );
NAND2_X1 MEM_stage_inst_dmem_U13900 ( .A1(MEM_stage_inst_dmem_ram_1923), .A2(MEM_stage_inst_dmem_n16237), .ZN(MEM_stage_inst_dmem_n16232) );
NAND2_X1 MEM_stage_inst_dmem_U13899 ( .A1(MEM_stage_inst_dmem_n16230), .A2(MEM_stage_inst_dmem_n16229), .ZN(MEM_stage_inst_dmem_n11199) );
NAND2_X1 MEM_stage_inst_dmem_U13898 ( .A1(MEM_stage_inst_dmem_n16368), .A2(MEM_stage_inst_dmem_n16238), .ZN(MEM_stage_inst_dmem_n16229) );
NAND2_X1 MEM_stage_inst_dmem_U13897 ( .A1(MEM_stage_inst_dmem_ram_1924), .A2(MEM_stage_inst_dmem_n16237), .ZN(MEM_stage_inst_dmem_n16230) );
NAND2_X1 MEM_stage_inst_dmem_U13896 ( .A1(MEM_stage_inst_dmem_n16228), .A2(MEM_stage_inst_dmem_n16227), .ZN(MEM_stage_inst_dmem_n11200) );
NAND2_X1 MEM_stage_inst_dmem_U13895 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n16238), .ZN(MEM_stage_inst_dmem_n16227) );
NAND2_X1 MEM_stage_inst_dmem_U13894 ( .A1(MEM_stage_inst_dmem_ram_1925), .A2(MEM_stage_inst_dmem_n16237), .ZN(MEM_stage_inst_dmem_n16228) );
NAND2_X1 MEM_stage_inst_dmem_U13893 ( .A1(MEM_stage_inst_dmem_n16226), .A2(MEM_stage_inst_dmem_n16225), .ZN(MEM_stage_inst_dmem_n11201) );
NAND2_X1 MEM_stage_inst_dmem_U13892 ( .A1(MEM_stage_inst_dmem_n14717), .A2(MEM_stage_inst_dmem_n16238), .ZN(MEM_stage_inst_dmem_n16225) );
NAND2_X1 MEM_stage_inst_dmem_U13891 ( .A1(MEM_stage_inst_dmem_ram_1926), .A2(MEM_stage_inst_dmem_n16237), .ZN(MEM_stage_inst_dmem_n16226) );
NAND2_X1 MEM_stage_inst_dmem_U13890 ( .A1(MEM_stage_inst_dmem_n16224), .A2(MEM_stage_inst_dmem_n16223), .ZN(MEM_stage_inst_dmem_n11202) );
NAND2_X1 MEM_stage_inst_dmem_U13889 ( .A1(MEM_stage_inst_dmem_n112), .A2(MEM_stage_inst_dmem_n16238), .ZN(MEM_stage_inst_dmem_n16223) );
NAND2_X1 MEM_stage_inst_dmem_U13888 ( .A1(MEM_stage_inst_dmem_ram_1927), .A2(MEM_stage_inst_dmem_n16237), .ZN(MEM_stage_inst_dmem_n16224) );
NAND2_X1 MEM_stage_inst_dmem_U13887 ( .A1(MEM_stage_inst_dmem_n16222), .A2(MEM_stage_inst_dmem_n16221), .ZN(MEM_stage_inst_dmem_n11203) );
NAND2_X1 MEM_stage_inst_dmem_U13886 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n16238), .ZN(MEM_stage_inst_dmem_n16221) );
NAND2_X1 MEM_stage_inst_dmem_U13885 ( .A1(MEM_stage_inst_dmem_ram_1928), .A2(MEM_stage_inst_dmem_n16237), .ZN(MEM_stage_inst_dmem_n16222) );
NAND2_X1 MEM_stage_inst_dmem_U13884 ( .A1(MEM_stage_inst_dmem_n16220), .A2(MEM_stage_inst_dmem_n16219), .ZN(MEM_stage_inst_dmem_n11204) );
NAND2_X1 MEM_stage_inst_dmem_U13883 ( .A1(MEM_stage_inst_dmem_n19251), .A2(MEM_stage_inst_dmem_n16238), .ZN(MEM_stage_inst_dmem_n16219) );
NAND2_X1 MEM_stage_inst_dmem_U13882 ( .A1(MEM_stage_inst_dmem_ram_1929), .A2(MEM_stage_inst_dmem_n16237), .ZN(MEM_stage_inst_dmem_n16220) );
NAND2_X1 MEM_stage_inst_dmem_U13881 ( .A1(MEM_stage_inst_dmem_n16218), .A2(MEM_stage_inst_dmem_n16217), .ZN(MEM_stage_inst_dmem_n11205) );
NAND2_X1 MEM_stage_inst_dmem_U13880 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n16238), .ZN(MEM_stage_inst_dmem_n16217) );
NAND2_X1 MEM_stage_inst_dmem_U13879 ( .A1(MEM_stage_inst_dmem_ram_1930), .A2(MEM_stage_inst_dmem_n16237), .ZN(MEM_stage_inst_dmem_n16218) );
NAND2_X1 MEM_stage_inst_dmem_U13878 ( .A1(MEM_stage_inst_dmem_n16216), .A2(MEM_stage_inst_dmem_n16215), .ZN(MEM_stage_inst_dmem_n11206) );
NAND2_X1 MEM_stage_inst_dmem_U13877 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n16238), .ZN(MEM_stage_inst_dmem_n16215) );
NAND2_X1 MEM_stage_inst_dmem_U13876 ( .A1(MEM_stage_inst_dmem_ram_1931), .A2(MEM_stage_inst_dmem_n16237), .ZN(MEM_stage_inst_dmem_n16216) );
NAND2_X1 MEM_stage_inst_dmem_U13875 ( .A1(MEM_stage_inst_dmem_n16214), .A2(MEM_stage_inst_dmem_n16213), .ZN(MEM_stage_inst_dmem_n11207) );
NAND2_X1 MEM_stage_inst_dmem_U13874 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n16238), .ZN(MEM_stage_inst_dmem_n16213) );
NAND2_X1 MEM_stage_inst_dmem_U13873 ( .A1(MEM_stage_inst_dmem_ram_1932), .A2(MEM_stage_inst_dmem_n16237), .ZN(MEM_stage_inst_dmem_n16214) );
NAND2_X1 MEM_stage_inst_dmem_U13872 ( .A1(MEM_stage_inst_dmem_n16212), .A2(MEM_stage_inst_dmem_n16211), .ZN(MEM_stage_inst_dmem_n11208) );
NAND2_X1 MEM_stage_inst_dmem_U13871 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n16238), .ZN(MEM_stage_inst_dmem_n16211) );
NAND2_X1 MEM_stage_inst_dmem_U13870 ( .A1(MEM_stage_inst_dmem_ram_1933), .A2(MEM_stage_inst_dmem_n16237), .ZN(MEM_stage_inst_dmem_n16212) );
NAND2_X1 MEM_stage_inst_dmem_U13869 ( .A1(MEM_stage_inst_dmem_n16210), .A2(MEM_stage_inst_dmem_n16209), .ZN(MEM_stage_inst_dmem_n11209) );
NAND2_X1 MEM_stage_inst_dmem_U13868 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n16238), .ZN(MEM_stage_inst_dmem_n16209) );
NAND2_X1 MEM_stage_inst_dmem_U13867 ( .A1(MEM_stage_inst_dmem_ram_1934), .A2(MEM_stage_inst_dmem_n16237), .ZN(MEM_stage_inst_dmem_n16210) );
NAND2_X1 MEM_stage_inst_dmem_U13866 ( .A1(MEM_stage_inst_dmem_n16208), .A2(MEM_stage_inst_dmem_n16207), .ZN(MEM_stage_inst_dmem_n11210) );
NAND2_X1 MEM_stage_inst_dmem_U13865 ( .A1(MEM_stage_inst_dmem_n15110), .A2(MEM_stage_inst_dmem_n16238), .ZN(MEM_stage_inst_dmem_n16207) );
INV_X1 MEM_stage_inst_dmem_U13864 ( .A(MEM_stage_inst_dmem_n16237), .ZN(MEM_stage_inst_dmem_n16238) );
NAND2_X1 MEM_stage_inst_dmem_U13863 ( .A1(MEM_stage_inst_dmem_ram_1935), .A2(MEM_stage_inst_dmem_n16237), .ZN(MEM_stage_inst_dmem_n16208) );
NAND2_X1 MEM_stage_inst_dmem_U13862 ( .A1(MEM_stage_inst_dmem_n21179), .A2(MEM_stage_inst_dmem_n16484), .ZN(MEM_stage_inst_dmem_n16237) );
NAND2_X1 MEM_stage_inst_dmem_U13861 ( .A1(MEM_stage_inst_dmem_n16206), .A2(MEM_stage_inst_dmem_n16205), .ZN(MEM_stage_inst_dmem_n11211) );
NAND2_X1 MEM_stage_inst_dmem_U13860 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n16204), .ZN(MEM_stage_inst_dmem_n16205) );
NAND2_X1 MEM_stage_inst_dmem_U13859 ( .A1(MEM_stage_inst_dmem_ram_1936), .A2(MEM_stage_inst_dmem_n16203), .ZN(MEM_stage_inst_dmem_n16206) );
NAND2_X1 MEM_stage_inst_dmem_U13858 ( .A1(MEM_stage_inst_dmem_n16202), .A2(MEM_stage_inst_dmem_n16201), .ZN(MEM_stage_inst_dmem_n11212) );
NAND2_X1 MEM_stage_inst_dmem_U13857 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n16204), .ZN(MEM_stage_inst_dmem_n16201) );
NAND2_X1 MEM_stage_inst_dmem_U13856 ( .A1(MEM_stage_inst_dmem_ram_1937), .A2(MEM_stage_inst_dmem_n16203), .ZN(MEM_stage_inst_dmem_n16202) );
NAND2_X1 MEM_stage_inst_dmem_U13855 ( .A1(MEM_stage_inst_dmem_n16200), .A2(MEM_stage_inst_dmem_n16199), .ZN(MEM_stage_inst_dmem_n11213) );
NAND2_X1 MEM_stage_inst_dmem_U13854 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n16204), .ZN(MEM_stage_inst_dmem_n16199) );
NAND2_X1 MEM_stage_inst_dmem_U13853 ( .A1(MEM_stage_inst_dmem_ram_1938), .A2(MEM_stage_inst_dmem_n16203), .ZN(MEM_stage_inst_dmem_n16200) );
NAND2_X1 MEM_stage_inst_dmem_U13852 ( .A1(MEM_stage_inst_dmem_n16198), .A2(MEM_stage_inst_dmem_n16197), .ZN(MEM_stage_inst_dmem_n11214) );
NAND2_X1 MEM_stage_inst_dmem_U13851 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n16204), .ZN(MEM_stage_inst_dmem_n16197) );
NAND2_X1 MEM_stage_inst_dmem_U13850 ( .A1(MEM_stage_inst_dmem_ram_1939), .A2(MEM_stage_inst_dmem_n16203), .ZN(MEM_stage_inst_dmem_n16198) );
NAND2_X1 MEM_stage_inst_dmem_U13849 ( .A1(MEM_stage_inst_dmem_n16196), .A2(MEM_stage_inst_dmem_n16195), .ZN(MEM_stage_inst_dmem_n11215) );
NAND2_X1 MEM_stage_inst_dmem_U13848 ( .A1(MEM_stage_inst_dmem_n16368), .A2(MEM_stage_inst_dmem_n16204), .ZN(MEM_stage_inst_dmem_n16195) );
NAND2_X1 MEM_stage_inst_dmem_U13847 ( .A1(MEM_stage_inst_dmem_ram_1940), .A2(MEM_stage_inst_dmem_n16203), .ZN(MEM_stage_inst_dmem_n16196) );
NAND2_X1 MEM_stage_inst_dmem_U13846 ( .A1(MEM_stage_inst_dmem_n16194), .A2(MEM_stage_inst_dmem_n16193), .ZN(MEM_stage_inst_dmem_n11216) );
NAND2_X1 MEM_stage_inst_dmem_U13845 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n16204), .ZN(MEM_stage_inst_dmem_n16193) );
NAND2_X1 MEM_stage_inst_dmem_U13844 ( .A1(MEM_stage_inst_dmem_ram_1941), .A2(MEM_stage_inst_dmem_n16203), .ZN(MEM_stage_inst_dmem_n16194) );
NAND2_X1 MEM_stage_inst_dmem_U13843 ( .A1(MEM_stage_inst_dmem_n16192), .A2(MEM_stage_inst_dmem_n16191), .ZN(MEM_stage_inst_dmem_n11217) );
NAND2_X1 MEM_stage_inst_dmem_U13842 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n16204), .ZN(MEM_stage_inst_dmem_n16191) );
NAND2_X1 MEM_stage_inst_dmem_U13841 ( .A1(MEM_stage_inst_dmem_ram_1942), .A2(MEM_stage_inst_dmem_n16203), .ZN(MEM_stage_inst_dmem_n16192) );
NAND2_X1 MEM_stage_inst_dmem_U13840 ( .A1(MEM_stage_inst_dmem_n16190), .A2(MEM_stage_inst_dmem_n16189), .ZN(MEM_stage_inst_dmem_n11218) );
NAND2_X1 MEM_stage_inst_dmem_U13839 ( .A1(MEM_stage_inst_dmem_n16361), .A2(MEM_stage_inst_dmem_n16204), .ZN(MEM_stage_inst_dmem_n16189) );
NAND2_X1 MEM_stage_inst_dmem_U13838 ( .A1(MEM_stage_inst_dmem_ram_1943), .A2(MEM_stage_inst_dmem_n16203), .ZN(MEM_stage_inst_dmem_n16190) );
NAND2_X1 MEM_stage_inst_dmem_U13837 ( .A1(MEM_stage_inst_dmem_n16188), .A2(MEM_stage_inst_dmem_n16187), .ZN(MEM_stage_inst_dmem_n11219) );
NAND2_X1 MEM_stage_inst_dmem_U13836 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n16204), .ZN(MEM_stage_inst_dmem_n16187) );
NAND2_X1 MEM_stage_inst_dmem_U13835 ( .A1(MEM_stage_inst_dmem_ram_1944), .A2(MEM_stage_inst_dmem_n16203), .ZN(MEM_stage_inst_dmem_n16188) );
NAND2_X1 MEM_stage_inst_dmem_U13834 ( .A1(MEM_stage_inst_dmem_n16186), .A2(MEM_stage_inst_dmem_n16185), .ZN(MEM_stage_inst_dmem_n11220) );
NAND2_X1 MEM_stage_inst_dmem_U13833 ( .A1(MEM_stage_inst_dmem_n16772), .A2(MEM_stage_inst_dmem_n16204), .ZN(MEM_stage_inst_dmem_n16185) );
NAND2_X1 MEM_stage_inst_dmem_U13832 ( .A1(MEM_stage_inst_dmem_ram_1945), .A2(MEM_stage_inst_dmem_n16203), .ZN(MEM_stage_inst_dmem_n16186) );
NAND2_X1 MEM_stage_inst_dmem_U13831 ( .A1(MEM_stage_inst_dmem_n16184), .A2(MEM_stage_inst_dmem_n16183), .ZN(MEM_stage_inst_dmem_n11221) );
NAND2_X1 MEM_stage_inst_dmem_U13830 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n16204), .ZN(MEM_stage_inst_dmem_n16183) );
NAND2_X1 MEM_stage_inst_dmem_U13829 ( .A1(MEM_stage_inst_dmem_ram_1946), .A2(MEM_stage_inst_dmem_n16203), .ZN(MEM_stage_inst_dmem_n16184) );
NAND2_X1 MEM_stage_inst_dmem_U13828 ( .A1(MEM_stage_inst_dmem_n16182), .A2(MEM_stage_inst_dmem_n16181), .ZN(MEM_stage_inst_dmem_n11222) );
NAND2_X1 MEM_stage_inst_dmem_U13827 ( .A1(MEM_stage_inst_dmem_n20518), .A2(MEM_stage_inst_dmem_n16204), .ZN(MEM_stage_inst_dmem_n16181) );
NAND2_X1 MEM_stage_inst_dmem_U13826 ( .A1(MEM_stage_inst_dmem_ram_1947), .A2(MEM_stage_inst_dmem_n16203), .ZN(MEM_stage_inst_dmem_n16182) );
NAND2_X1 MEM_stage_inst_dmem_U13825 ( .A1(MEM_stage_inst_dmem_n16180), .A2(MEM_stage_inst_dmem_n16179), .ZN(MEM_stage_inst_dmem_n11223) );
NAND2_X1 MEM_stage_inst_dmem_U13824 ( .A1(MEM_stage_inst_dmem_n20515), .A2(MEM_stage_inst_dmem_n16204), .ZN(MEM_stage_inst_dmem_n16179) );
NAND2_X1 MEM_stage_inst_dmem_U13823 ( .A1(MEM_stage_inst_dmem_ram_1948), .A2(MEM_stage_inst_dmem_n16203), .ZN(MEM_stage_inst_dmem_n16180) );
NAND2_X1 MEM_stage_inst_dmem_U13822 ( .A1(MEM_stage_inst_dmem_n16178), .A2(MEM_stage_inst_dmem_n16177), .ZN(MEM_stage_inst_dmem_n11224) );
NAND2_X1 MEM_stage_inst_dmem_U13821 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n16204), .ZN(MEM_stage_inst_dmem_n16177) );
NAND2_X1 MEM_stage_inst_dmem_U13820 ( .A1(MEM_stage_inst_dmem_ram_1949), .A2(MEM_stage_inst_dmem_n16203), .ZN(MEM_stage_inst_dmem_n16178) );
NAND2_X1 MEM_stage_inst_dmem_U13819 ( .A1(MEM_stage_inst_dmem_n16176), .A2(MEM_stage_inst_dmem_n16175), .ZN(MEM_stage_inst_dmem_n11225) );
NAND2_X1 MEM_stage_inst_dmem_U13818 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n16204), .ZN(MEM_stage_inst_dmem_n16175) );
NAND2_X1 MEM_stage_inst_dmem_U13817 ( .A1(MEM_stage_inst_dmem_ram_1950), .A2(MEM_stage_inst_dmem_n16203), .ZN(MEM_stage_inst_dmem_n16176) );
NAND2_X1 MEM_stage_inst_dmem_U13816 ( .A1(MEM_stage_inst_dmem_n16174), .A2(MEM_stage_inst_dmem_n16173), .ZN(MEM_stage_inst_dmem_n11226) );
NAND2_X1 MEM_stage_inst_dmem_U13815 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n16204), .ZN(MEM_stage_inst_dmem_n16173) );
INV_X1 MEM_stage_inst_dmem_U13814 ( .A(MEM_stage_inst_dmem_n16203), .ZN(MEM_stage_inst_dmem_n16204) );
NAND2_X1 MEM_stage_inst_dmem_U13813 ( .A1(MEM_stage_inst_dmem_ram_1951), .A2(MEM_stage_inst_dmem_n16203), .ZN(MEM_stage_inst_dmem_n16174) );
NAND2_X1 MEM_stage_inst_dmem_U13812 ( .A1(MEM_stage_inst_dmem_n21144), .A2(MEM_stage_inst_dmem_n16484), .ZN(MEM_stage_inst_dmem_n16203) );
NAND2_X1 MEM_stage_inst_dmem_U13811 ( .A1(MEM_stage_inst_dmem_n16172), .A2(MEM_stage_inst_dmem_n16171), .ZN(MEM_stage_inst_dmem_n11227) );
NAND2_X1 MEM_stage_inst_dmem_U13810 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n16170), .ZN(MEM_stage_inst_dmem_n16171) );
NAND2_X1 MEM_stage_inst_dmem_U13809 ( .A1(MEM_stage_inst_dmem_ram_1952), .A2(MEM_stage_inst_dmem_n16169), .ZN(MEM_stage_inst_dmem_n16172) );
NAND2_X1 MEM_stage_inst_dmem_U13808 ( .A1(MEM_stage_inst_dmem_n16168), .A2(MEM_stage_inst_dmem_n16167), .ZN(MEM_stage_inst_dmem_n11228) );
NAND2_X1 MEM_stage_inst_dmem_U13807 ( .A1(MEM_stage_inst_dmem_n20547), .A2(MEM_stage_inst_dmem_n16170), .ZN(MEM_stage_inst_dmem_n16167) );
NAND2_X1 MEM_stage_inst_dmem_U13806 ( .A1(MEM_stage_inst_dmem_ram_1953), .A2(MEM_stage_inst_dmem_n16169), .ZN(MEM_stage_inst_dmem_n16168) );
NAND2_X1 MEM_stage_inst_dmem_U13805 ( .A1(MEM_stage_inst_dmem_n16166), .A2(MEM_stage_inst_dmem_n16165), .ZN(MEM_stage_inst_dmem_n11229) );
NAND2_X1 MEM_stage_inst_dmem_U13804 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n16170), .ZN(MEM_stage_inst_dmem_n16165) );
NAND2_X1 MEM_stage_inst_dmem_U13803 ( .A1(MEM_stage_inst_dmem_ram_1954), .A2(MEM_stage_inst_dmem_n16169), .ZN(MEM_stage_inst_dmem_n16166) );
NAND2_X1 MEM_stage_inst_dmem_U13802 ( .A1(MEM_stage_inst_dmem_n16164), .A2(MEM_stage_inst_dmem_n16163), .ZN(MEM_stage_inst_dmem_n11230) );
NAND2_X1 MEM_stage_inst_dmem_U13801 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n16170), .ZN(MEM_stage_inst_dmem_n16163) );
NAND2_X1 MEM_stage_inst_dmem_U13800 ( .A1(MEM_stage_inst_dmem_ram_1955), .A2(MEM_stage_inst_dmem_n16169), .ZN(MEM_stage_inst_dmem_n16164) );
NAND2_X1 MEM_stage_inst_dmem_U13799 ( .A1(MEM_stage_inst_dmem_n16162), .A2(MEM_stage_inst_dmem_n16161), .ZN(MEM_stage_inst_dmem_n11231) );
NAND2_X1 MEM_stage_inst_dmem_U13798 ( .A1(MEM_stage_inst_dmem_n16368), .A2(MEM_stage_inst_dmem_n16170), .ZN(MEM_stage_inst_dmem_n16161) );
NAND2_X1 MEM_stage_inst_dmem_U13797 ( .A1(MEM_stage_inst_dmem_ram_1956), .A2(MEM_stage_inst_dmem_n16169), .ZN(MEM_stage_inst_dmem_n16162) );
NAND2_X1 MEM_stage_inst_dmem_U13796 ( .A1(MEM_stage_inst_dmem_n16160), .A2(MEM_stage_inst_dmem_n16159), .ZN(MEM_stage_inst_dmem_n11232) );
NAND2_X1 MEM_stage_inst_dmem_U13795 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n16170), .ZN(MEM_stage_inst_dmem_n16159) );
NAND2_X1 MEM_stage_inst_dmem_U13794 ( .A1(MEM_stage_inst_dmem_ram_1957), .A2(MEM_stage_inst_dmem_n16169), .ZN(MEM_stage_inst_dmem_n16160) );
NAND2_X1 MEM_stage_inst_dmem_U13793 ( .A1(MEM_stage_inst_dmem_n16158), .A2(MEM_stage_inst_dmem_n16157), .ZN(MEM_stage_inst_dmem_n11233) );
NAND2_X1 MEM_stage_inst_dmem_U13792 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n16170), .ZN(MEM_stage_inst_dmem_n16157) );
NAND2_X1 MEM_stage_inst_dmem_U13791 ( .A1(MEM_stage_inst_dmem_ram_1958), .A2(MEM_stage_inst_dmem_n16169), .ZN(MEM_stage_inst_dmem_n16158) );
NAND2_X1 MEM_stage_inst_dmem_U13790 ( .A1(MEM_stage_inst_dmem_n16156), .A2(MEM_stage_inst_dmem_n16155), .ZN(MEM_stage_inst_dmem_n11234) );
NAND2_X1 MEM_stage_inst_dmem_U13789 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n16170), .ZN(MEM_stage_inst_dmem_n16155) );
NAND2_X1 MEM_stage_inst_dmem_U13788 ( .A1(MEM_stage_inst_dmem_ram_1959), .A2(MEM_stage_inst_dmem_n16169), .ZN(MEM_stage_inst_dmem_n16156) );
NAND2_X1 MEM_stage_inst_dmem_U13787 ( .A1(MEM_stage_inst_dmem_n16154), .A2(MEM_stage_inst_dmem_n16153), .ZN(MEM_stage_inst_dmem_n11235) );
NAND2_X1 MEM_stage_inst_dmem_U13786 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n16170), .ZN(MEM_stage_inst_dmem_n16153) );
NAND2_X1 MEM_stage_inst_dmem_U13785 ( .A1(MEM_stage_inst_dmem_ram_1960), .A2(MEM_stage_inst_dmem_n16169), .ZN(MEM_stage_inst_dmem_n16154) );
NAND2_X1 MEM_stage_inst_dmem_U13784 ( .A1(MEM_stage_inst_dmem_n16152), .A2(MEM_stage_inst_dmem_n16151), .ZN(MEM_stage_inst_dmem_n11236) );
NAND2_X1 MEM_stage_inst_dmem_U13783 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n16170), .ZN(MEM_stage_inst_dmem_n16151) );
NAND2_X1 MEM_stage_inst_dmem_U13782 ( .A1(MEM_stage_inst_dmem_ram_1961), .A2(MEM_stage_inst_dmem_n16169), .ZN(MEM_stage_inst_dmem_n16152) );
NAND2_X1 MEM_stage_inst_dmem_U13781 ( .A1(MEM_stage_inst_dmem_n16150), .A2(MEM_stage_inst_dmem_n16149), .ZN(MEM_stage_inst_dmem_n11237) );
NAND2_X1 MEM_stage_inst_dmem_U13780 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n16170), .ZN(MEM_stage_inst_dmem_n16149) );
NAND2_X1 MEM_stage_inst_dmem_U13779 ( .A1(MEM_stage_inst_dmem_ram_1962), .A2(MEM_stage_inst_dmem_n16169), .ZN(MEM_stage_inst_dmem_n16150) );
NAND2_X1 MEM_stage_inst_dmem_U13778 ( .A1(MEM_stage_inst_dmem_n16148), .A2(MEM_stage_inst_dmem_n16147), .ZN(MEM_stage_inst_dmem_n11238) );
NAND2_X1 MEM_stage_inst_dmem_U13777 ( .A1(MEM_stage_inst_dmem_n13044), .A2(MEM_stage_inst_dmem_n16170), .ZN(MEM_stage_inst_dmem_n16147) );
NAND2_X1 MEM_stage_inst_dmem_U13776 ( .A1(MEM_stage_inst_dmem_ram_1963), .A2(MEM_stage_inst_dmem_n16169), .ZN(MEM_stage_inst_dmem_n16148) );
NAND2_X1 MEM_stage_inst_dmem_U13775 ( .A1(MEM_stage_inst_dmem_n16146), .A2(MEM_stage_inst_dmem_n16145), .ZN(MEM_stage_inst_dmem_n11239) );
NAND2_X1 MEM_stage_inst_dmem_U13774 ( .A1(MEM_stage_inst_dmem_n13041), .A2(MEM_stage_inst_dmem_n16170), .ZN(MEM_stage_inst_dmem_n16145) );
NAND2_X1 MEM_stage_inst_dmem_U13773 ( .A1(MEM_stage_inst_dmem_ram_1964), .A2(MEM_stage_inst_dmem_n16169), .ZN(MEM_stage_inst_dmem_n16146) );
NAND2_X1 MEM_stage_inst_dmem_U13772 ( .A1(MEM_stage_inst_dmem_n16144), .A2(MEM_stage_inst_dmem_n16143), .ZN(MEM_stage_inst_dmem_n11240) );
NAND2_X1 MEM_stage_inst_dmem_U13771 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n16170), .ZN(MEM_stage_inst_dmem_n16143) );
NAND2_X1 MEM_stage_inst_dmem_U13770 ( .A1(MEM_stage_inst_dmem_ram_1965), .A2(MEM_stage_inst_dmem_n16169), .ZN(MEM_stage_inst_dmem_n16144) );
NAND2_X1 MEM_stage_inst_dmem_U13769 ( .A1(MEM_stage_inst_dmem_n16142), .A2(MEM_stage_inst_dmem_n16141), .ZN(MEM_stage_inst_dmem_n11241) );
NAND2_X1 MEM_stage_inst_dmem_U13768 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n16170), .ZN(MEM_stage_inst_dmem_n16141) );
NAND2_X1 MEM_stage_inst_dmem_U13767 ( .A1(MEM_stage_inst_dmem_ram_1966), .A2(MEM_stage_inst_dmem_n16169), .ZN(MEM_stage_inst_dmem_n16142) );
NAND2_X1 MEM_stage_inst_dmem_U13766 ( .A1(MEM_stage_inst_dmem_n16140), .A2(MEM_stage_inst_dmem_n16139), .ZN(MEM_stage_inst_dmem_n11242) );
NAND2_X1 MEM_stage_inst_dmem_U13765 ( .A1(MEM_stage_inst_dmem_n16343), .A2(MEM_stage_inst_dmem_n16170), .ZN(MEM_stage_inst_dmem_n16139) );
INV_X1 MEM_stage_inst_dmem_U13764 ( .A(MEM_stage_inst_dmem_n16169), .ZN(MEM_stage_inst_dmem_n16170) );
NAND2_X1 MEM_stage_inst_dmem_U13763 ( .A1(MEM_stage_inst_dmem_ram_1967), .A2(MEM_stage_inst_dmem_n16169), .ZN(MEM_stage_inst_dmem_n16140) );
NAND2_X1 MEM_stage_inst_dmem_U13762 ( .A1(MEM_stage_inst_dmem_n21109), .A2(MEM_stage_inst_dmem_n16484), .ZN(MEM_stage_inst_dmem_n16169) );
NAND2_X1 MEM_stage_inst_dmem_U13761 ( .A1(MEM_stage_inst_dmem_n16138), .A2(MEM_stage_inst_dmem_n16137), .ZN(MEM_stage_inst_dmem_n11243) );
NAND2_X1 MEM_stage_inst_dmem_U13760 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n16136), .ZN(MEM_stage_inst_dmem_n16137) );
NAND2_X1 MEM_stage_inst_dmem_U13759 ( .A1(MEM_stage_inst_dmem_ram_1968), .A2(MEM_stage_inst_dmem_n16135), .ZN(MEM_stage_inst_dmem_n16138) );
NAND2_X1 MEM_stage_inst_dmem_U13758 ( .A1(MEM_stage_inst_dmem_n16134), .A2(MEM_stage_inst_dmem_n16133), .ZN(MEM_stage_inst_dmem_n11244) );
NAND2_X1 MEM_stage_inst_dmem_U13757 ( .A1(MEM_stage_inst_dmem_n109), .A2(MEM_stage_inst_dmem_n16136), .ZN(MEM_stage_inst_dmem_n16133) );
NAND2_X1 MEM_stage_inst_dmem_U13756 ( .A1(MEM_stage_inst_dmem_ram_1969), .A2(MEM_stage_inst_dmem_n16135), .ZN(MEM_stage_inst_dmem_n16134) );
NAND2_X1 MEM_stage_inst_dmem_U13755 ( .A1(MEM_stage_inst_dmem_n16132), .A2(MEM_stage_inst_dmem_n16131), .ZN(MEM_stage_inst_dmem_n11245) );
NAND2_X1 MEM_stage_inst_dmem_U13754 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n16136), .ZN(MEM_stage_inst_dmem_n16131) );
NAND2_X1 MEM_stage_inst_dmem_U13753 ( .A1(MEM_stage_inst_dmem_ram_1970), .A2(MEM_stage_inst_dmem_n16135), .ZN(MEM_stage_inst_dmem_n16132) );
NAND2_X1 MEM_stage_inst_dmem_U13752 ( .A1(MEM_stage_inst_dmem_n16130), .A2(MEM_stage_inst_dmem_n16129), .ZN(MEM_stage_inst_dmem_n11246) );
NAND2_X1 MEM_stage_inst_dmem_U13751 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n16136), .ZN(MEM_stage_inst_dmem_n16129) );
NAND2_X1 MEM_stage_inst_dmem_U13750 ( .A1(MEM_stage_inst_dmem_ram_1971), .A2(MEM_stage_inst_dmem_n16135), .ZN(MEM_stage_inst_dmem_n16130) );
NAND2_X1 MEM_stage_inst_dmem_U13749 ( .A1(MEM_stage_inst_dmem_n16128), .A2(MEM_stage_inst_dmem_n16127), .ZN(MEM_stage_inst_dmem_n11247) );
NAND2_X1 MEM_stage_inst_dmem_U13748 ( .A1(MEM_stage_inst_dmem_n16368), .A2(MEM_stage_inst_dmem_n16136), .ZN(MEM_stage_inst_dmem_n16127) );
NAND2_X1 MEM_stage_inst_dmem_U13747 ( .A1(MEM_stage_inst_dmem_ram_1972), .A2(MEM_stage_inst_dmem_n16135), .ZN(MEM_stage_inst_dmem_n16128) );
NAND2_X1 MEM_stage_inst_dmem_U13746 ( .A1(MEM_stage_inst_dmem_n16126), .A2(MEM_stage_inst_dmem_n16125), .ZN(MEM_stage_inst_dmem_n11248) );
NAND2_X1 MEM_stage_inst_dmem_U13745 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n16136), .ZN(MEM_stage_inst_dmem_n16125) );
NAND2_X1 MEM_stage_inst_dmem_U13744 ( .A1(MEM_stage_inst_dmem_ram_1973), .A2(MEM_stage_inst_dmem_n16135), .ZN(MEM_stage_inst_dmem_n16126) );
NAND2_X1 MEM_stage_inst_dmem_U13743 ( .A1(MEM_stage_inst_dmem_n16124), .A2(MEM_stage_inst_dmem_n16123), .ZN(MEM_stage_inst_dmem_n11249) );
NAND2_X1 MEM_stage_inst_dmem_U13742 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n16136), .ZN(MEM_stage_inst_dmem_n16123) );
NAND2_X1 MEM_stage_inst_dmem_U13741 ( .A1(MEM_stage_inst_dmem_ram_1974), .A2(MEM_stage_inst_dmem_n16135), .ZN(MEM_stage_inst_dmem_n16124) );
NAND2_X1 MEM_stage_inst_dmem_U13740 ( .A1(MEM_stage_inst_dmem_n16122), .A2(MEM_stage_inst_dmem_n16121), .ZN(MEM_stage_inst_dmem_n11250) );
NAND2_X1 MEM_stage_inst_dmem_U13739 ( .A1(MEM_stage_inst_dmem_n16361), .A2(MEM_stage_inst_dmem_n16136), .ZN(MEM_stage_inst_dmem_n16121) );
NAND2_X1 MEM_stage_inst_dmem_U13738 ( .A1(MEM_stage_inst_dmem_ram_1975), .A2(MEM_stage_inst_dmem_n16135), .ZN(MEM_stage_inst_dmem_n16122) );
NAND2_X1 MEM_stage_inst_dmem_U13737 ( .A1(MEM_stage_inst_dmem_n16120), .A2(MEM_stage_inst_dmem_n16119), .ZN(MEM_stage_inst_dmem_n11251) );
NAND2_X1 MEM_stage_inst_dmem_U13736 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n16136), .ZN(MEM_stage_inst_dmem_n16119) );
NAND2_X1 MEM_stage_inst_dmem_U13735 ( .A1(MEM_stage_inst_dmem_ram_1976), .A2(MEM_stage_inst_dmem_n16135), .ZN(MEM_stage_inst_dmem_n16120) );
NAND2_X1 MEM_stage_inst_dmem_U13734 ( .A1(MEM_stage_inst_dmem_n16118), .A2(MEM_stage_inst_dmem_n16117), .ZN(MEM_stage_inst_dmem_n11252) );
NAND2_X1 MEM_stage_inst_dmem_U13733 ( .A1(MEM_stage_inst_dmem_n96), .A2(MEM_stage_inst_dmem_n16136), .ZN(MEM_stage_inst_dmem_n16117) );
NAND2_X1 MEM_stage_inst_dmem_U13732 ( .A1(MEM_stage_inst_dmem_ram_1977), .A2(MEM_stage_inst_dmem_n16135), .ZN(MEM_stage_inst_dmem_n16118) );
NAND2_X1 MEM_stage_inst_dmem_U13731 ( .A1(MEM_stage_inst_dmem_n16116), .A2(MEM_stage_inst_dmem_n16115), .ZN(MEM_stage_inst_dmem_n11253) );
NAND2_X1 MEM_stage_inst_dmem_U13730 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n16136), .ZN(MEM_stage_inst_dmem_n16115) );
NAND2_X1 MEM_stage_inst_dmem_U13729 ( .A1(MEM_stage_inst_dmem_ram_1978), .A2(MEM_stage_inst_dmem_n16135), .ZN(MEM_stage_inst_dmem_n16116) );
NAND2_X1 MEM_stage_inst_dmem_U13728 ( .A1(MEM_stage_inst_dmem_n16114), .A2(MEM_stage_inst_dmem_n16113), .ZN(MEM_stage_inst_dmem_n11254) );
NAND2_X1 MEM_stage_inst_dmem_U13727 ( .A1(MEM_stage_inst_dmem_n14705), .A2(MEM_stage_inst_dmem_n16136), .ZN(MEM_stage_inst_dmem_n16113) );
NAND2_X1 MEM_stage_inst_dmem_U13726 ( .A1(MEM_stage_inst_dmem_ram_1979), .A2(MEM_stage_inst_dmem_n16135), .ZN(MEM_stage_inst_dmem_n16114) );
NAND2_X1 MEM_stage_inst_dmem_U13725 ( .A1(MEM_stage_inst_dmem_n16112), .A2(MEM_stage_inst_dmem_n16111), .ZN(MEM_stage_inst_dmem_n11255) );
NAND2_X1 MEM_stage_inst_dmem_U13724 ( .A1(MEM_stage_inst_dmem_n14702), .A2(MEM_stage_inst_dmem_n16136), .ZN(MEM_stage_inst_dmem_n16111) );
NAND2_X1 MEM_stage_inst_dmem_U13723 ( .A1(MEM_stage_inst_dmem_ram_1980), .A2(MEM_stage_inst_dmem_n16135), .ZN(MEM_stage_inst_dmem_n16112) );
NAND2_X1 MEM_stage_inst_dmem_U13722 ( .A1(MEM_stage_inst_dmem_n16110), .A2(MEM_stage_inst_dmem_n16109), .ZN(MEM_stage_inst_dmem_n11256) );
NAND2_X1 MEM_stage_inst_dmem_U13721 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n16136), .ZN(MEM_stage_inst_dmem_n16109) );
NAND2_X1 MEM_stage_inst_dmem_U13720 ( .A1(MEM_stage_inst_dmem_ram_1981), .A2(MEM_stage_inst_dmem_n16135), .ZN(MEM_stage_inst_dmem_n16110) );
NAND2_X1 MEM_stage_inst_dmem_U13719 ( .A1(MEM_stage_inst_dmem_n16108), .A2(MEM_stage_inst_dmem_n16107), .ZN(MEM_stage_inst_dmem_n11257) );
NAND2_X1 MEM_stage_inst_dmem_U13718 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n16136), .ZN(MEM_stage_inst_dmem_n16107) );
NAND2_X1 MEM_stage_inst_dmem_U13717 ( .A1(MEM_stage_inst_dmem_ram_1982), .A2(MEM_stage_inst_dmem_n16135), .ZN(MEM_stage_inst_dmem_n16108) );
NAND2_X1 MEM_stage_inst_dmem_U13716 ( .A1(MEM_stage_inst_dmem_n16106), .A2(MEM_stage_inst_dmem_n16105), .ZN(MEM_stage_inst_dmem_n11258) );
NAND2_X1 MEM_stage_inst_dmem_U13715 ( .A1(MEM_stage_inst_dmem_n14693), .A2(MEM_stage_inst_dmem_n16136), .ZN(MEM_stage_inst_dmem_n16105) );
INV_X1 MEM_stage_inst_dmem_U13714 ( .A(MEM_stage_inst_dmem_n16135), .ZN(MEM_stage_inst_dmem_n16136) );
NAND2_X1 MEM_stage_inst_dmem_U13713 ( .A1(MEM_stage_inst_dmem_ram_1983), .A2(MEM_stage_inst_dmem_n16135), .ZN(MEM_stage_inst_dmem_n16106) );
NAND2_X1 MEM_stage_inst_dmem_U13712 ( .A1(MEM_stage_inst_dmem_n21074), .A2(MEM_stage_inst_dmem_n16484), .ZN(MEM_stage_inst_dmem_n16135) );
NAND2_X1 MEM_stage_inst_dmem_U13711 ( .A1(MEM_stage_inst_dmem_n16104), .A2(MEM_stage_inst_dmem_n16103), .ZN(MEM_stage_inst_dmem_n11259) );
NAND2_X1 MEM_stage_inst_dmem_U13710 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n16102), .ZN(MEM_stage_inst_dmem_n16103) );
NAND2_X1 MEM_stage_inst_dmem_U13709 ( .A1(MEM_stage_inst_dmem_ram_1984), .A2(MEM_stage_inst_dmem_n16101), .ZN(MEM_stage_inst_dmem_n16104) );
NAND2_X1 MEM_stage_inst_dmem_U13708 ( .A1(MEM_stage_inst_dmem_n16100), .A2(MEM_stage_inst_dmem_n16099), .ZN(MEM_stage_inst_dmem_n11260) );
NAND2_X1 MEM_stage_inst_dmem_U13707 ( .A1(EX_pipeline_reg_out_6), .A2(MEM_stage_inst_dmem_n16102), .ZN(MEM_stage_inst_dmem_n16099) );
NAND2_X1 MEM_stage_inst_dmem_U13706 ( .A1(MEM_stage_inst_dmem_ram_1985), .A2(MEM_stage_inst_dmem_n16101), .ZN(MEM_stage_inst_dmem_n16100) );
NAND2_X1 MEM_stage_inst_dmem_U13705 ( .A1(MEM_stage_inst_dmem_n16098), .A2(MEM_stage_inst_dmem_n16097), .ZN(MEM_stage_inst_dmem_n11261) );
NAND2_X1 MEM_stage_inst_dmem_U13704 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n16102), .ZN(MEM_stage_inst_dmem_n16097) );
NAND2_X1 MEM_stage_inst_dmem_U13703 ( .A1(MEM_stage_inst_dmem_ram_1986), .A2(MEM_stage_inst_dmem_n16101), .ZN(MEM_stage_inst_dmem_n16098) );
NAND2_X1 MEM_stage_inst_dmem_U13702 ( .A1(MEM_stage_inst_dmem_n16096), .A2(MEM_stage_inst_dmem_n16095), .ZN(MEM_stage_inst_dmem_n11262) );
NAND2_X1 MEM_stage_inst_dmem_U13701 ( .A1(MEM_stage_inst_dmem_n13064), .A2(MEM_stage_inst_dmem_n16102), .ZN(MEM_stage_inst_dmem_n16095) );
NAND2_X1 MEM_stage_inst_dmem_U13700 ( .A1(MEM_stage_inst_dmem_ram_1987), .A2(MEM_stage_inst_dmem_n16101), .ZN(MEM_stage_inst_dmem_n16096) );
NAND2_X1 MEM_stage_inst_dmem_U13699 ( .A1(MEM_stage_inst_dmem_n16094), .A2(MEM_stage_inst_dmem_n16093), .ZN(MEM_stage_inst_dmem_n11263) );
NAND2_X1 MEM_stage_inst_dmem_U13698 ( .A1(MEM_stage_inst_dmem_n16368), .A2(MEM_stage_inst_dmem_n16102), .ZN(MEM_stage_inst_dmem_n16093) );
NAND2_X1 MEM_stage_inst_dmem_U13697 ( .A1(MEM_stage_inst_dmem_ram_1988), .A2(MEM_stage_inst_dmem_n16101), .ZN(MEM_stage_inst_dmem_n16094) );
NAND2_X1 MEM_stage_inst_dmem_U13696 ( .A1(MEM_stage_inst_dmem_n16092), .A2(MEM_stage_inst_dmem_n16091), .ZN(MEM_stage_inst_dmem_n11264) );
NAND2_X1 MEM_stage_inst_dmem_U13695 ( .A1(MEM_stage_inst_dmem_n13059), .A2(MEM_stage_inst_dmem_n16102), .ZN(MEM_stage_inst_dmem_n16091) );
NAND2_X1 MEM_stage_inst_dmem_U13694 ( .A1(MEM_stage_inst_dmem_ram_1989), .A2(MEM_stage_inst_dmem_n16101), .ZN(MEM_stage_inst_dmem_n16092) );
NAND2_X1 MEM_stage_inst_dmem_U13693 ( .A1(MEM_stage_inst_dmem_n16090), .A2(MEM_stage_inst_dmem_n16089), .ZN(MEM_stage_inst_dmem_n11265) );
NAND2_X1 MEM_stage_inst_dmem_U13692 ( .A1(MEM_stage_inst_dmem_n13056), .A2(MEM_stage_inst_dmem_n16102), .ZN(MEM_stage_inst_dmem_n16089) );
NAND2_X1 MEM_stage_inst_dmem_U13691 ( .A1(MEM_stage_inst_dmem_ram_1990), .A2(MEM_stage_inst_dmem_n16101), .ZN(MEM_stage_inst_dmem_n16090) );
NAND2_X1 MEM_stage_inst_dmem_U13690 ( .A1(MEM_stage_inst_dmem_n16088), .A2(MEM_stage_inst_dmem_n16087), .ZN(MEM_stage_inst_dmem_n11266) );
NAND2_X1 MEM_stage_inst_dmem_U13689 ( .A1(MEM_stage_inst_dmem_n112), .A2(MEM_stage_inst_dmem_n16102), .ZN(MEM_stage_inst_dmem_n16087) );
NAND2_X1 MEM_stage_inst_dmem_U13688 ( .A1(MEM_stage_inst_dmem_ram_1991), .A2(MEM_stage_inst_dmem_n16101), .ZN(MEM_stage_inst_dmem_n16088) );
NAND2_X1 MEM_stage_inst_dmem_U13687 ( .A1(MEM_stage_inst_dmem_n16086), .A2(MEM_stage_inst_dmem_n16085), .ZN(MEM_stage_inst_dmem_n11267) );
NAND2_X1 MEM_stage_inst_dmem_U13686 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n16102), .ZN(MEM_stage_inst_dmem_n16085) );
NAND2_X1 MEM_stage_inst_dmem_U13685 ( .A1(MEM_stage_inst_dmem_ram_1992), .A2(MEM_stage_inst_dmem_n16101), .ZN(MEM_stage_inst_dmem_n16086) );
NAND2_X1 MEM_stage_inst_dmem_U13684 ( .A1(MEM_stage_inst_dmem_n16084), .A2(MEM_stage_inst_dmem_n16083), .ZN(MEM_stage_inst_dmem_n11268) );
NAND2_X1 MEM_stage_inst_dmem_U13683 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n16102), .ZN(MEM_stage_inst_dmem_n16083) );
NAND2_X1 MEM_stage_inst_dmem_U13682 ( .A1(MEM_stage_inst_dmem_ram_1993), .A2(MEM_stage_inst_dmem_n16101), .ZN(MEM_stage_inst_dmem_n16084) );
NAND2_X1 MEM_stage_inst_dmem_U13681 ( .A1(MEM_stage_inst_dmem_n16082), .A2(MEM_stage_inst_dmem_n16081), .ZN(MEM_stage_inst_dmem_n11269) );
NAND2_X1 MEM_stage_inst_dmem_U13680 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n16102), .ZN(MEM_stage_inst_dmem_n16081) );
NAND2_X1 MEM_stage_inst_dmem_U13679 ( .A1(MEM_stage_inst_dmem_ram_1994), .A2(MEM_stage_inst_dmem_n16101), .ZN(MEM_stage_inst_dmem_n16082) );
NAND2_X1 MEM_stage_inst_dmem_U13678 ( .A1(MEM_stage_inst_dmem_n16080), .A2(MEM_stage_inst_dmem_n16079), .ZN(MEM_stage_inst_dmem_n11270) );
NAND2_X1 MEM_stage_inst_dmem_U13677 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n16102), .ZN(MEM_stage_inst_dmem_n16079) );
NAND2_X1 MEM_stage_inst_dmem_U13676 ( .A1(MEM_stage_inst_dmem_ram_1995), .A2(MEM_stage_inst_dmem_n16101), .ZN(MEM_stage_inst_dmem_n16080) );
NAND2_X1 MEM_stage_inst_dmem_U13675 ( .A1(MEM_stage_inst_dmem_n16078), .A2(MEM_stage_inst_dmem_n16077), .ZN(MEM_stage_inst_dmem_n11271) );
NAND2_X1 MEM_stage_inst_dmem_U13674 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n16102), .ZN(MEM_stage_inst_dmem_n16077) );
NAND2_X1 MEM_stage_inst_dmem_U13673 ( .A1(MEM_stage_inst_dmem_ram_1996), .A2(MEM_stage_inst_dmem_n16101), .ZN(MEM_stage_inst_dmem_n16078) );
NAND2_X1 MEM_stage_inst_dmem_U13672 ( .A1(MEM_stage_inst_dmem_n16076), .A2(MEM_stage_inst_dmem_n16075), .ZN(MEM_stage_inst_dmem_n11272) );
NAND2_X1 MEM_stage_inst_dmem_U13671 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n16102), .ZN(MEM_stage_inst_dmem_n16075) );
NAND2_X1 MEM_stage_inst_dmem_U13670 ( .A1(MEM_stage_inst_dmem_ram_1997), .A2(MEM_stage_inst_dmem_n16101), .ZN(MEM_stage_inst_dmem_n16076) );
NAND2_X1 MEM_stage_inst_dmem_U13669 ( .A1(MEM_stage_inst_dmem_n16074), .A2(MEM_stage_inst_dmem_n16073), .ZN(MEM_stage_inst_dmem_n11273) );
NAND2_X1 MEM_stage_inst_dmem_U13668 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n16102), .ZN(MEM_stage_inst_dmem_n16073) );
NAND2_X1 MEM_stage_inst_dmem_U13667 ( .A1(MEM_stage_inst_dmem_ram_1998), .A2(MEM_stage_inst_dmem_n16101), .ZN(MEM_stage_inst_dmem_n16074) );
NAND2_X1 MEM_stage_inst_dmem_U13666 ( .A1(MEM_stage_inst_dmem_n16072), .A2(MEM_stage_inst_dmem_n16071), .ZN(MEM_stage_inst_dmem_n11274) );
NAND2_X1 MEM_stage_inst_dmem_U13665 ( .A1(MEM_stage_inst_dmem_n15110), .A2(MEM_stage_inst_dmem_n16102), .ZN(MEM_stage_inst_dmem_n16071) );
INV_X1 MEM_stage_inst_dmem_U13664 ( .A(MEM_stage_inst_dmem_n16101), .ZN(MEM_stage_inst_dmem_n16102) );
NAND2_X1 MEM_stage_inst_dmem_U13663 ( .A1(MEM_stage_inst_dmem_ram_1999), .A2(MEM_stage_inst_dmem_n16101), .ZN(MEM_stage_inst_dmem_n16072) );
NAND2_X1 MEM_stage_inst_dmem_U13662 ( .A1(MEM_stage_inst_dmem_n21039), .A2(MEM_stage_inst_dmem_n16484), .ZN(MEM_stage_inst_dmem_n16101) );
NAND2_X1 MEM_stage_inst_dmem_U13661 ( .A1(MEM_stage_inst_dmem_n16070), .A2(MEM_stage_inst_dmem_n16069), .ZN(MEM_stage_inst_dmem_n11275) );
NAND2_X1 MEM_stage_inst_dmem_U13660 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n16068), .ZN(MEM_stage_inst_dmem_n16069) );
NAND2_X1 MEM_stage_inst_dmem_U13659 ( .A1(MEM_stage_inst_dmem_ram_2000), .A2(MEM_stage_inst_dmem_n16067), .ZN(MEM_stage_inst_dmem_n16070) );
NAND2_X1 MEM_stage_inst_dmem_U13658 ( .A1(MEM_stage_inst_dmem_n16066), .A2(MEM_stage_inst_dmem_n16065), .ZN(MEM_stage_inst_dmem_n11276) );
NAND2_X1 MEM_stage_inst_dmem_U13657 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n16068), .ZN(MEM_stage_inst_dmem_n16065) );
NAND2_X1 MEM_stage_inst_dmem_U13656 ( .A1(MEM_stage_inst_dmem_ram_2001), .A2(MEM_stage_inst_dmem_n16067), .ZN(MEM_stage_inst_dmem_n16066) );
NAND2_X1 MEM_stage_inst_dmem_U13655 ( .A1(MEM_stage_inst_dmem_n16064), .A2(MEM_stage_inst_dmem_n16063), .ZN(MEM_stage_inst_dmem_n11277) );
NAND2_X1 MEM_stage_inst_dmem_U13654 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n16068), .ZN(MEM_stage_inst_dmem_n16063) );
NAND2_X1 MEM_stage_inst_dmem_U13653 ( .A1(MEM_stage_inst_dmem_ram_2002), .A2(MEM_stage_inst_dmem_n16067), .ZN(MEM_stage_inst_dmem_n16064) );
NAND2_X1 MEM_stage_inst_dmem_U13652 ( .A1(MEM_stage_inst_dmem_n16062), .A2(MEM_stage_inst_dmem_n16061), .ZN(MEM_stage_inst_dmem_n11278) );
NAND2_X1 MEM_stage_inst_dmem_U13651 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n16068), .ZN(MEM_stage_inst_dmem_n16061) );
NAND2_X1 MEM_stage_inst_dmem_U13650 ( .A1(MEM_stage_inst_dmem_ram_2003), .A2(MEM_stage_inst_dmem_n16067), .ZN(MEM_stage_inst_dmem_n16062) );
NAND2_X1 MEM_stage_inst_dmem_U13649 ( .A1(MEM_stage_inst_dmem_n16060), .A2(MEM_stage_inst_dmem_n16059), .ZN(MEM_stage_inst_dmem_n11279) );
NAND2_X1 MEM_stage_inst_dmem_U13648 ( .A1(MEM_stage_inst_dmem_n16368), .A2(MEM_stage_inst_dmem_n16068), .ZN(MEM_stage_inst_dmem_n16059) );
NAND2_X1 MEM_stage_inst_dmem_U13647 ( .A1(MEM_stage_inst_dmem_ram_2004), .A2(MEM_stage_inst_dmem_n16067), .ZN(MEM_stage_inst_dmem_n16060) );
NAND2_X1 MEM_stage_inst_dmem_U13646 ( .A1(MEM_stage_inst_dmem_n16058), .A2(MEM_stage_inst_dmem_n16057), .ZN(MEM_stage_inst_dmem_n11280) );
NAND2_X1 MEM_stage_inst_dmem_U13645 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n16068), .ZN(MEM_stage_inst_dmem_n16057) );
NAND2_X1 MEM_stage_inst_dmem_U13644 ( .A1(MEM_stage_inst_dmem_ram_2005), .A2(MEM_stage_inst_dmem_n16067), .ZN(MEM_stage_inst_dmem_n16058) );
NAND2_X1 MEM_stage_inst_dmem_U13643 ( .A1(MEM_stage_inst_dmem_n16056), .A2(MEM_stage_inst_dmem_n16055), .ZN(MEM_stage_inst_dmem_n11281) );
NAND2_X1 MEM_stage_inst_dmem_U13642 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n16068), .ZN(MEM_stage_inst_dmem_n16055) );
NAND2_X1 MEM_stage_inst_dmem_U13641 ( .A1(MEM_stage_inst_dmem_ram_2006), .A2(MEM_stage_inst_dmem_n16067), .ZN(MEM_stage_inst_dmem_n16056) );
NAND2_X1 MEM_stage_inst_dmem_U13640 ( .A1(MEM_stage_inst_dmem_n16054), .A2(MEM_stage_inst_dmem_n16053), .ZN(MEM_stage_inst_dmem_n11282) );
NAND2_X1 MEM_stage_inst_dmem_U13639 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n16068), .ZN(MEM_stage_inst_dmem_n16053) );
NAND2_X1 MEM_stage_inst_dmem_U13638 ( .A1(MEM_stage_inst_dmem_ram_2007), .A2(MEM_stage_inst_dmem_n16067), .ZN(MEM_stage_inst_dmem_n16054) );
NAND2_X1 MEM_stage_inst_dmem_U13637 ( .A1(MEM_stage_inst_dmem_n16052), .A2(MEM_stage_inst_dmem_n16051), .ZN(MEM_stage_inst_dmem_n11283) );
NAND2_X1 MEM_stage_inst_dmem_U13636 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n16068), .ZN(MEM_stage_inst_dmem_n16051) );
NAND2_X1 MEM_stage_inst_dmem_U13635 ( .A1(MEM_stage_inst_dmem_ram_2008), .A2(MEM_stage_inst_dmem_n16067), .ZN(MEM_stage_inst_dmem_n16052) );
NAND2_X1 MEM_stage_inst_dmem_U13634 ( .A1(MEM_stage_inst_dmem_n16050), .A2(MEM_stage_inst_dmem_n16049), .ZN(MEM_stage_inst_dmem_n11284) );
NAND2_X1 MEM_stage_inst_dmem_U13633 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n16068), .ZN(MEM_stage_inst_dmem_n16049) );
NAND2_X1 MEM_stage_inst_dmem_U13632 ( .A1(MEM_stage_inst_dmem_ram_2009), .A2(MEM_stage_inst_dmem_n16067), .ZN(MEM_stage_inst_dmem_n16050) );
NAND2_X1 MEM_stage_inst_dmem_U13631 ( .A1(MEM_stage_inst_dmem_n16048), .A2(MEM_stage_inst_dmem_n16047), .ZN(MEM_stage_inst_dmem_n11285) );
NAND2_X1 MEM_stage_inst_dmem_U13630 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n16068), .ZN(MEM_stage_inst_dmem_n16047) );
NAND2_X1 MEM_stage_inst_dmem_U13629 ( .A1(MEM_stage_inst_dmem_ram_2010), .A2(MEM_stage_inst_dmem_n16067), .ZN(MEM_stage_inst_dmem_n16048) );
NAND2_X1 MEM_stage_inst_dmem_U13628 ( .A1(MEM_stage_inst_dmem_n16046), .A2(MEM_stage_inst_dmem_n16045), .ZN(MEM_stage_inst_dmem_n11286) );
NAND2_X1 MEM_stage_inst_dmem_U13627 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n16068), .ZN(MEM_stage_inst_dmem_n16045) );
NAND2_X1 MEM_stage_inst_dmem_U13626 ( .A1(MEM_stage_inst_dmem_ram_2011), .A2(MEM_stage_inst_dmem_n16067), .ZN(MEM_stage_inst_dmem_n16046) );
NAND2_X1 MEM_stage_inst_dmem_U13625 ( .A1(MEM_stage_inst_dmem_n16044), .A2(MEM_stage_inst_dmem_n16043), .ZN(MEM_stage_inst_dmem_n11287) );
NAND2_X1 MEM_stage_inst_dmem_U13624 ( .A1(MEM_stage_inst_dmem_n14702), .A2(MEM_stage_inst_dmem_n16068), .ZN(MEM_stage_inst_dmem_n16043) );
NAND2_X1 MEM_stage_inst_dmem_U13623 ( .A1(MEM_stage_inst_dmem_ram_2012), .A2(MEM_stage_inst_dmem_n16067), .ZN(MEM_stage_inst_dmem_n16044) );
NAND2_X1 MEM_stage_inst_dmem_U13622 ( .A1(MEM_stage_inst_dmem_n16042), .A2(MEM_stage_inst_dmem_n16041), .ZN(MEM_stage_inst_dmem_n11288) );
NAND2_X1 MEM_stage_inst_dmem_U13621 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n16068), .ZN(MEM_stage_inst_dmem_n16041) );
NAND2_X1 MEM_stage_inst_dmem_U13620 ( .A1(MEM_stage_inst_dmem_ram_2013), .A2(MEM_stage_inst_dmem_n16067), .ZN(MEM_stage_inst_dmem_n16042) );
NAND2_X1 MEM_stage_inst_dmem_U13619 ( .A1(MEM_stage_inst_dmem_n16040), .A2(MEM_stage_inst_dmem_n16039), .ZN(MEM_stage_inst_dmem_n11289) );
NAND2_X1 MEM_stage_inst_dmem_U13618 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n16068), .ZN(MEM_stage_inst_dmem_n16039) );
NAND2_X1 MEM_stage_inst_dmem_U13617 ( .A1(MEM_stage_inst_dmem_ram_2014), .A2(MEM_stage_inst_dmem_n16067), .ZN(MEM_stage_inst_dmem_n16040) );
NAND2_X1 MEM_stage_inst_dmem_U13616 ( .A1(MEM_stage_inst_dmem_n16038), .A2(MEM_stage_inst_dmem_n16037), .ZN(MEM_stage_inst_dmem_n11290) );
NAND2_X1 MEM_stage_inst_dmem_U13615 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n16068), .ZN(MEM_stage_inst_dmem_n16037) );
INV_X1 MEM_stage_inst_dmem_U13614 ( .A(MEM_stage_inst_dmem_n16067), .ZN(MEM_stage_inst_dmem_n16068) );
NAND2_X1 MEM_stage_inst_dmem_U13613 ( .A1(MEM_stage_inst_dmem_ram_2015), .A2(MEM_stage_inst_dmem_n16067), .ZN(MEM_stage_inst_dmem_n16038) );
NAND2_X1 MEM_stage_inst_dmem_U13612 ( .A1(MEM_stage_inst_dmem_n21004), .A2(MEM_stage_inst_dmem_n16484), .ZN(MEM_stage_inst_dmem_n16067) );
NAND2_X1 MEM_stage_inst_dmem_U13611 ( .A1(MEM_stage_inst_dmem_n16036), .A2(MEM_stage_inst_dmem_n16035), .ZN(MEM_stage_inst_dmem_n11291) );
NAND2_X1 MEM_stage_inst_dmem_U13610 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n16034), .ZN(MEM_stage_inst_dmem_n16035) );
NAND2_X1 MEM_stage_inst_dmem_U13609 ( .A1(MEM_stage_inst_dmem_ram_2016), .A2(MEM_stage_inst_dmem_n16033), .ZN(MEM_stage_inst_dmem_n16036) );
NAND2_X1 MEM_stage_inst_dmem_U13608 ( .A1(MEM_stage_inst_dmem_n16032), .A2(MEM_stage_inst_dmem_n16031), .ZN(MEM_stage_inst_dmem_n11292) );
NAND2_X1 MEM_stage_inst_dmem_U13607 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n16034), .ZN(MEM_stage_inst_dmem_n16031) );
NAND2_X1 MEM_stage_inst_dmem_U13606 ( .A1(MEM_stage_inst_dmem_ram_2017), .A2(MEM_stage_inst_dmem_n16033), .ZN(MEM_stage_inst_dmem_n16032) );
NAND2_X1 MEM_stage_inst_dmem_U13605 ( .A1(MEM_stage_inst_dmem_n16030), .A2(MEM_stage_inst_dmem_n16029), .ZN(MEM_stage_inst_dmem_n11293) );
NAND2_X1 MEM_stage_inst_dmem_U13604 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n16034), .ZN(MEM_stage_inst_dmem_n16029) );
NAND2_X1 MEM_stage_inst_dmem_U13603 ( .A1(MEM_stage_inst_dmem_ram_2018), .A2(MEM_stage_inst_dmem_n16033), .ZN(MEM_stage_inst_dmem_n16030) );
NAND2_X1 MEM_stage_inst_dmem_U13602 ( .A1(MEM_stage_inst_dmem_n16028), .A2(MEM_stage_inst_dmem_n16027), .ZN(MEM_stage_inst_dmem_n11294) );
NAND2_X1 MEM_stage_inst_dmem_U13601 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n16034), .ZN(MEM_stage_inst_dmem_n16027) );
NAND2_X1 MEM_stage_inst_dmem_U13600 ( .A1(MEM_stage_inst_dmem_ram_2019), .A2(MEM_stage_inst_dmem_n16033), .ZN(MEM_stage_inst_dmem_n16028) );
NAND2_X1 MEM_stage_inst_dmem_U13599 ( .A1(MEM_stage_inst_dmem_n16026), .A2(MEM_stage_inst_dmem_n16025), .ZN(MEM_stage_inst_dmem_n11295) );
NAND2_X1 MEM_stage_inst_dmem_U13598 ( .A1(MEM_stage_inst_dmem_n16368), .A2(MEM_stage_inst_dmem_n16034), .ZN(MEM_stage_inst_dmem_n16025) );
NAND2_X1 MEM_stage_inst_dmem_U13597 ( .A1(MEM_stage_inst_dmem_ram_2020), .A2(MEM_stage_inst_dmem_n16033), .ZN(MEM_stage_inst_dmem_n16026) );
NAND2_X1 MEM_stage_inst_dmem_U13596 ( .A1(MEM_stage_inst_dmem_n16024), .A2(MEM_stage_inst_dmem_n16023), .ZN(MEM_stage_inst_dmem_n11296) );
NAND2_X1 MEM_stage_inst_dmem_U13595 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n16034), .ZN(MEM_stage_inst_dmem_n16023) );
NAND2_X1 MEM_stage_inst_dmem_U13594 ( .A1(MEM_stage_inst_dmem_ram_2021), .A2(MEM_stage_inst_dmem_n16033), .ZN(MEM_stage_inst_dmem_n16024) );
NAND2_X1 MEM_stage_inst_dmem_U13593 ( .A1(MEM_stage_inst_dmem_n16022), .A2(MEM_stage_inst_dmem_n16021), .ZN(MEM_stage_inst_dmem_n11297) );
NAND2_X1 MEM_stage_inst_dmem_U13592 ( .A1(MEM_stage_inst_dmem_n14717), .A2(MEM_stage_inst_dmem_n16034), .ZN(MEM_stage_inst_dmem_n16021) );
NAND2_X1 MEM_stage_inst_dmem_U13591 ( .A1(MEM_stage_inst_dmem_ram_2022), .A2(MEM_stage_inst_dmem_n16033), .ZN(MEM_stage_inst_dmem_n16022) );
NAND2_X1 MEM_stage_inst_dmem_U13590 ( .A1(MEM_stage_inst_dmem_n16020), .A2(MEM_stage_inst_dmem_n16019), .ZN(MEM_stage_inst_dmem_n11298) );
NAND2_X1 MEM_stage_inst_dmem_U13589 ( .A1(MEM_stage_inst_dmem_n112), .A2(MEM_stage_inst_dmem_n16034), .ZN(MEM_stage_inst_dmem_n16019) );
NAND2_X1 MEM_stage_inst_dmem_U13588 ( .A1(MEM_stage_inst_dmem_ram_2023), .A2(MEM_stage_inst_dmem_n16033), .ZN(MEM_stage_inst_dmem_n16020) );
NAND2_X1 MEM_stage_inst_dmem_U13587 ( .A1(MEM_stage_inst_dmem_n16018), .A2(MEM_stage_inst_dmem_n16017), .ZN(MEM_stage_inst_dmem_n11299) );
NAND2_X1 MEM_stage_inst_dmem_U13586 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n16034), .ZN(MEM_stage_inst_dmem_n16017) );
NAND2_X1 MEM_stage_inst_dmem_U13585 ( .A1(MEM_stage_inst_dmem_ram_2024), .A2(MEM_stage_inst_dmem_n16033), .ZN(MEM_stage_inst_dmem_n16018) );
NAND2_X1 MEM_stage_inst_dmem_U13584 ( .A1(MEM_stage_inst_dmem_n16016), .A2(MEM_stage_inst_dmem_n16015), .ZN(MEM_stage_inst_dmem_n11300) );
NAND2_X1 MEM_stage_inst_dmem_U13583 ( .A1(MEM_stage_inst_dmem_n19251), .A2(MEM_stage_inst_dmem_n16034), .ZN(MEM_stage_inst_dmem_n16015) );
NAND2_X1 MEM_stage_inst_dmem_U13582 ( .A1(MEM_stage_inst_dmem_ram_2025), .A2(MEM_stage_inst_dmem_n16033), .ZN(MEM_stage_inst_dmem_n16016) );
NAND2_X1 MEM_stage_inst_dmem_U13581 ( .A1(MEM_stage_inst_dmem_n16014), .A2(MEM_stage_inst_dmem_n16013), .ZN(MEM_stage_inst_dmem_n11301) );
NAND2_X1 MEM_stage_inst_dmem_U13580 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n16034), .ZN(MEM_stage_inst_dmem_n16013) );
NAND2_X1 MEM_stage_inst_dmem_U13579 ( .A1(MEM_stage_inst_dmem_ram_2026), .A2(MEM_stage_inst_dmem_n16033), .ZN(MEM_stage_inst_dmem_n16014) );
NAND2_X1 MEM_stage_inst_dmem_U13578 ( .A1(MEM_stage_inst_dmem_n16012), .A2(MEM_stage_inst_dmem_n16011), .ZN(MEM_stage_inst_dmem_n11302) );
NAND2_X1 MEM_stage_inst_dmem_U13577 ( .A1(MEM_stage_inst_dmem_n18004), .A2(MEM_stage_inst_dmem_n16034), .ZN(MEM_stage_inst_dmem_n16011) );
NAND2_X1 MEM_stage_inst_dmem_U13576 ( .A1(MEM_stage_inst_dmem_ram_2027), .A2(MEM_stage_inst_dmem_n16033), .ZN(MEM_stage_inst_dmem_n16012) );
NAND2_X1 MEM_stage_inst_dmem_U13575 ( .A1(MEM_stage_inst_dmem_n16010), .A2(MEM_stage_inst_dmem_n16009), .ZN(MEM_stage_inst_dmem_n11303) );
NAND2_X1 MEM_stage_inst_dmem_U13574 ( .A1(MEM_stage_inst_dmem_n18001), .A2(MEM_stage_inst_dmem_n16034), .ZN(MEM_stage_inst_dmem_n16009) );
NAND2_X1 MEM_stage_inst_dmem_U13573 ( .A1(MEM_stage_inst_dmem_ram_2028), .A2(MEM_stage_inst_dmem_n16033), .ZN(MEM_stage_inst_dmem_n16010) );
NAND2_X1 MEM_stage_inst_dmem_U13572 ( .A1(MEM_stage_inst_dmem_n16008), .A2(MEM_stage_inst_dmem_n16007), .ZN(MEM_stage_inst_dmem_n11304) );
NAND2_X1 MEM_stage_inst_dmem_U13571 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n16034), .ZN(MEM_stage_inst_dmem_n16007) );
NAND2_X1 MEM_stage_inst_dmem_U13570 ( .A1(MEM_stage_inst_dmem_ram_2029), .A2(MEM_stage_inst_dmem_n16033), .ZN(MEM_stage_inst_dmem_n16008) );
NAND2_X1 MEM_stage_inst_dmem_U13569 ( .A1(MEM_stage_inst_dmem_n16006), .A2(MEM_stage_inst_dmem_n16005), .ZN(MEM_stage_inst_dmem_n11305) );
NAND2_X1 MEM_stage_inst_dmem_U13568 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n16034), .ZN(MEM_stage_inst_dmem_n16005) );
NAND2_X1 MEM_stage_inst_dmem_U13567 ( .A1(MEM_stage_inst_dmem_ram_2030), .A2(MEM_stage_inst_dmem_n16033), .ZN(MEM_stage_inst_dmem_n16006) );
NAND2_X1 MEM_stage_inst_dmem_U13566 ( .A1(MEM_stage_inst_dmem_n16004), .A2(MEM_stage_inst_dmem_n16003), .ZN(MEM_stage_inst_dmem_n11306) );
NAND2_X1 MEM_stage_inst_dmem_U13565 ( .A1(MEM_stage_inst_dmem_n16343), .A2(MEM_stage_inst_dmem_n16034), .ZN(MEM_stage_inst_dmem_n16003) );
INV_X1 MEM_stage_inst_dmem_U13564 ( .A(MEM_stage_inst_dmem_n16033), .ZN(MEM_stage_inst_dmem_n16034) );
NAND2_X1 MEM_stage_inst_dmem_U13563 ( .A1(MEM_stage_inst_dmem_ram_2031), .A2(MEM_stage_inst_dmem_n16033), .ZN(MEM_stage_inst_dmem_n16004) );
NAND2_X1 MEM_stage_inst_dmem_U13562 ( .A1(MEM_stage_inst_dmem_n20969), .A2(MEM_stage_inst_dmem_n16484), .ZN(MEM_stage_inst_dmem_n16033) );
NAND2_X1 MEM_stage_inst_dmem_U13561 ( .A1(MEM_stage_inst_dmem_n16002), .A2(MEM_stage_inst_dmem_n16001), .ZN(MEM_stage_inst_dmem_n11307) );
NAND2_X1 MEM_stage_inst_dmem_U13560 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n16000), .ZN(MEM_stage_inst_dmem_n16001) );
NAND2_X1 MEM_stage_inst_dmem_U13559 ( .A1(MEM_stage_inst_dmem_ram_2032), .A2(MEM_stage_inst_dmem_n15999), .ZN(MEM_stage_inst_dmem_n16002) );
NAND2_X1 MEM_stage_inst_dmem_U13558 ( .A1(MEM_stage_inst_dmem_n15998), .A2(MEM_stage_inst_dmem_n15997), .ZN(MEM_stage_inst_dmem_n11308) );
NAND2_X1 MEM_stage_inst_dmem_U13557 ( .A1(MEM_stage_inst_dmem_n20547), .A2(MEM_stage_inst_dmem_n16000), .ZN(MEM_stage_inst_dmem_n15997) );
NAND2_X1 MEM_stage_inst_dmem_U13556 ( .A1(MEM_stage_inst_dmem_ram_2033), .A2(MEM_stage_inst_dmem_n15999), .ZN(MEM_stage_inst_dmem_n15998) );
NAND2_X1 MEM_stage_inst_dmem_U13555 ( .A1(MEM_stage_inst_dmem_n15996), .A2(MEM_stage_inst_dmem_n15995), .ZN(MEM_stage_inst_dmem_n11309) );
NAND2_X1 MEM_stage_inst_dmem_U13554 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n16000), .ZN(MEM_stage_inst_dmem_n15995) );
NAND2_X1 MEM_stage_inst_dmem_U13553 ( .A1(MEM_stage_inst_dmem_ram_2034), .A2(MEM_stage_inst_dmem_n15999), .ZN(MEM_stage_inst_dmem_n15996) );
NAND2_X1 MEM_stage_inst_dmem_U13552 ( .A1(MEM_stage_inst_dmem_n15994), .A2(MEM_stage_inst_dmem_n15993), .ZN(MEM_stage_inst_dmem_n11310) );
NAND2_X1 MEM_stage_inst_dmem_U13551 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n16000), .ZN(MEM_stage_inst_dmem_n15993) );
NAND2_X1 MEM_stage_inst_dmem_U13550 ( .A1(MEM_stage_inst_dmem_ram_2035), .A2(MEM_stage_inst_dmem_n15999), .ZN(MEM_stage_inst_dmem_n15994) );
NAND2_X1 MEM_stage_inst_dmem_U13549 ( .A1(MEM_stage_inst_dmem_n15992), .A2(MEM_stage_inst_dmem_n15991), .ZN(MEM_stage_inst_dmem_n11311) );
NAND2_X1 MEM_stage_inst_dmem_U13548 ( .A1(MEM_stage_inst_dmem_n16368), .A2(MEM_stage_inst_dmem_n16000), .ZN(MEM_stage_inst_dmem_n15991) );
NAND2_X1 MEM_stage_inst_dmem_U13547 ( .A1(MEM_stage_inst_dmem_ram_2036), .A2(MEM_stage_inst_dmem_n15999), .ZN(MEM_stage_inst_dmem_n15992) );
NAND2_X1 MEM_stage_inst_dmem_U13546 ( .A1(MEM_stage_inst_dmem_n15990), .A2(MEM_stage_inst_dmem_n15989), .ZN(MEM_stage_inst_dmem_n11312) );
NAND2_X1 MEM_stage_inst_dmem_U13545 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n16000), .ZN(MEM_stage_inst_dmem_n15989) );
NAND2_X1 MEM_stage_inst_dmem_U13544 ( .A1(MEM_stage_inst_dmem_ram_2037), .A2(MEM_stage_inst_dmem_n15999), .ZN(MEM_stage_inst_dmem_n15990) );
NAND2_X1 MEM_stage_inst_dmem_U13543 ( .A1(MEM_stage_inst_dmem_n15988), .A2(MEM_stage_inst_dmem_n15987), .ZN(MEM_stage_inst_dmem_n11313) );
NAND2_X1 MEM_stage_inst_dmem_U13542 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n16000), .ZN(MEM_stage_inst_dmem_n15987) );
NAND2_X1 MEM_stage_inst_dmem_U13541 ( .A1(MEM_stage_inst_dmem_ram_2038), .A2(MEM_stage_inst_dmem_n15999), .ZN(MEM_stage_inst_dmem_n15988) );
NAND2_X1 MEM_stage_inst_dmem_U13540 ( .A1(MEM_stage_inst_dmem_n15986), .A2(MEM_stage_inst_dmem_n15985), .ZN(MEM_stage_inst_dmem_n11314) );
NAND2_X1 MEM_stage_inst_dmem_U13539 ( .A1(MEM_stage_inst_dmem_n16361), .A2(MEM_stage_inst_dmem_n16000), .ZN(MEM_stage_inst_dmem_n15985) );
NAND2_X1 MEM_stage_inst_dmem_U13538 ( .A1(MEM_stage_inst_dmem_ram_2039), .A2(MEM_stage_inst_dmem_n15999), .ZN(MEM_stage_inst_dmem_n15986) );
NAND2_X1 MEM_stage_inst_dmem_U13537 ( .A1(MEM_stage_inst_dmem_n15984), .A2(MEM_stage_inst_dmem_n15983), .ZN(MEM_stage_inst_dmem_n11315) );
NAND2_X1 MEM_stage_inst_dmem_U13536 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n16000), .ZN(MEM_stage_inst_dmem_n15983) );
NAND2_X1 MEM_stage_inst_dmem_U13535 ( .A1(MEM_stage_inst_dmem_ram_2040), .A2(MEM_stage_inst_dmem_n15999), .ZN(MEM_stage_inst_dmem_n15984) );
NAND2_X1 MEM_stage_inst_dmem_U13534 ( .A1(MEM_stage_inst_dmem_n15982), .A2(MEM_stage_inst_dmem_n15981), .ZN(MEM_stage_inst_dmem_n11316) );
NAND2_X1 MEM_stage_inst_dmem_U13533 ( .A1(MEM_stage_inst_dmem_n20524), .A2(MEM_stage_inst_dmem_n16000), .ZN(MEM_stage_inst_dmem_n15981) );
NAND2_X1 MEM_stage_inst_dmem_U13532 ( .A1(MEM_stage_inst_dmem_ram_2041), .A2(MEM_stage_inst_dmem_n15999), .ZN(MEM_stage_inst_dmem_n15982) );
NAND2_X1 MEM_stage_inst_dmem_U13531 ( .A1(MEM_stage_inst_dmem_n15980), .A2(MEM_stage_inst_dmem_n15979), .ZN(MEM_stage_inst_dmem_n11317) );
NAND2_X1 MEM_stage_inst_dmem_U13530 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n16000), .ZN(MEM_stage_inst_dmem_n15979) );
NAND2_X1 MEM_stage_inst_dmem_U13529 ( .A1(MEM_stage_inst_dmem_ram_2042), .A2(MEM_stage_inst_dmem_n15999), .ZN(MEM_stage_inst_dmem_n15980) );
NAND2_X1 MEM_stage_inst_dmem_U13528 ( .A1(MEM_stage_inst_dmem_n15978), .A2(MEM_stage_inst_dmem_n15977), .ZN(MEM_stage_inst_dmem_n11318) );
NAND2_X1 MEM_stage_inst_dmem_U13527 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n16000), .ZN(MEM_stage_inst_dmem_n15977) );
NAND2_X1 MEM_stage_inst_dmem_U13526 ( .A1(MEM_stage_inst_dmem_ram_2043), .A2(MEM_stage_inst_dmem_n15999), .ZN(MEM_stage_inst_dmem_n15978) );
NAND2_X1 MEM_stage_inst_dmem_U13525 ( .A1(MEM_stage_inst_dmem_n15976), .A2(MEM_stage_inst_dmem_n15975), .ZN(MEM_stage_inst_dmem_n11319) );
NAND2_X1 MEM_stage_inst_dmem_U13524 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n16000), .ZN(MEM_stage_inst_dmem_n15975) );
NAND2_X1 MEM_stage_inst_dmem_U13523 ( .A1(MEM_stage_inst_dmem_ram_2044), .A2(MEM_stage_inst_dmem_n15999), .ZN(MEM_stage_inst_dmem_n15976) );
NAND2_X1 MEM_stage_inst_dmem_U13522 ( .A1(MEM_stage_inst_dmem_n15974), .A2(MEM_stage_inst_dmem_n15973), .ZN(MEM_stage_inst_dmem_n11320) );
NAND2_X1 MEM_stage_inst_dmem_U13521 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n16000), .ZN(MEM_stage_inst_dmem_n15973) );
NAND2_X1 MEM_stage_inst_dmem_U13520 ( .A1(MEM_stage_inst_dmem_ram_2045), .A2(MEM_stage_inst_dmem_n15999), .ZN(MEM_stage_inst_dmem_n15974) );
NAND2_X1 MEM_stage_inst_dmem_U13519 ( .A1(MEM_stage_inst_dmem_n15972), .A2(MEM_stage_inst_dmem_n15971), .ZN(MEM_stage_inst_dmem_n11321) );
NAND2_X1 MEM_stage_inst_dmem_U13518 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n16000), .ZN(MEM_stage_inst_dmem_n15971) );
NAND2_X1 MEM_stage_inst_dmem_U13517 ( .A1(MEM_stage_inst_dmem_ram_2046), .A2(MEM_stage_inst_dmem_n15999), .ZN(MEM_stage_inst_dmem_n15972) );
NAND2_X1 MEM_stage_inst_dmem_U13516 ( .A1(MEM_stage_inst_dmem_n15970), .A2(MEM_stage_inst_dmem_n15969), .ZN(MEM_stage_inst_dmem_n11322) );
NAND2_X1 MEM_stage_inst_dmem_U13515 ( .A1(MEM_stage_inst_dmem_n14693), .A2(MEM_stage_inst_dmem_n16000), .ZN(MEM_stage_inst_dmem_n15969) );
INV_X1 MEM_stage_inst_dmem_U13514 ( .A(MEM_stage_inst_dmem_n15999), .ZN(MEM_stage_inst_dmem_n16000) );
BUF_X1 MEM_stage_inst_dmem_U13513 ( .A(MEM_stage_inst_dmem_n20506), .Z(MEM_stage_inst_dmem_n16343) );
NAND2_X1 MEM_stage_inst_dmem_U13512 ( .A1(MEM_stage_inst_dmem_ram_2047), .A2(MEM_stage_inst_dmem_n15999), .ZN(MEM_stage_inst_dmem_n15970) );
NAND2_X1 MEM_stage_inst_dmem_U13511 ( .A1(MEM_stage_inst_dmem_n20934), .A2(MEM_stage_inst_dmem_n16484), .ZN(MEM_stage_inst_dmem_n15999) );
NOR2_X2 MEM_stage_inst_dmem_U13510 ( .A1(MEM_stage_inst_dmem_n15968), .A2(MEM_stage_inst_dmem_n20933), .ZN(MEM_stage_inst_dmem_n16484) );
NAND2_X1 MEM_stage_inst_dmem_U13509 ( .A1(MEM_stage_inst_dmem_n15967), .A2(MEM_stage_inst_dmem_n15966), .ZN(MEM_stage_inst_dmem_n20933) );
NAND2_X1 MEM_stage_inst_dmem_U13508 ( .A1(MEM_stage_inst_dmem_n15965), .A2(MEM_stage_inst_dmem_n15964), .ZN(MEM_stage_inst_dmem_n11323) );
NAND2_X1 MEM_stage_inst_dmem_U13507 ( .A1(MEM_stage_inst_dmem_n19275), .A2(MEM_stage_inst_dmem_n15963), .ZN(MEM_stage_inst_dmem_n15964) );
NAND2_X1 MEM_stage_inst_dmem_U13506 ( .A1(MEM_stage_inst_dmem_ram_1024), .A2(MEM_stage_inst_dmem_n15962), .ZN(MEM_stage_inst_dmem_n15965) );
NAND2_X1 MEM_stage_inst_dmem_U13505 ( .A1(MEM_stage_inst_dmem_n15961), .A2(MEM_stage_inst_dmem_n15960), .ZN(MEM_stage_inst_dmem_n11324) );
NAND2_X1 MEM_stage_inst_dmem_U13504 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n15963), .ZN(MEM_stage_inst_dmem_n15960) );
NAND2_X1 MEM_stage_inst_dmem_U13503 ( .A1(MEM_stage_inst_dmem_ram_1025), .A2(MEM_stage_inst_dmem_n15962), .ZN(MEM_stage_inst_dmem_n15961) );
NAND2_X1 MEM_stage_inst_dmem_U13502 ( .A1(MEM_stage_inst_dmem_n15959), .A2(MEM_stage_inst_dmem_n15958), .ZN(MEM_stage_inst_dmem_n11325) );
NAND2_X1 MEM_stage_inst_dmem_U13501 ( .A1(MEM_stage_inst_dmem_n16789), .A2(MEM_stage_inst_dmem_n15963), .ZN(MEM_stage_inst_dmem_n15958) );
NAND2_X1 MEM_stage_inst_dmem_U13500 ( .A1(MEM_stage_inst_dmem_ram_1026), .A2(MEM_stage_inst_dmem_n15962), .ZN(MEM_stage_inst_dmem_n15959) );
NAND2_X1 MEM_stage_inst_dmem_U13499 ( .A1(MEM_stage_inst_dmem_n15957), .A2(MEM_stage_inst_dmem_n15956), .ZN(MEM_stage_inst_dmem_n11326) );
NAND2_X1 MEM_stage_inst_dmem_U13498 ( .A1(MEM_stage_inst_dmem_n13064), .A2(MEM_stage_inst_dmem_n15963), .ZN(MEM_stage_inst_dmem_n15956) );
NAND2_X1 MEM_stage_inst_dmem_U13497 ( .A1(MEM_stage_inst_dmem_ram_1027), .A2(MEM_stage_inst_dmem_n15962), .ZN(MEM_stage_inst_dmem_n15957) );
NAND2_X1 MEM_stage_inst_dmem_U13496 ( .A1(MEM_stage_inst_dmem_n15955), .A2(MEM_stage_inst_dmem_n15954), .ZN(MEM_stage_inst_dmem_n11327) );
NAND2_X1 MEM_stage_inst_dmem_U13495 ( .A1(MEM_stage_inst_dmem_n16784), .A2(MEM_stage_inst_dmem_n15963), .ZN(MEM_stage_inst_dmem_n15954) );
NAND2_X1 MEM_stage_inst_dmem_U13494 ( .A1(MEM_stage_inst_dmem_ram_1028), .A2(MEM_stage_inst_dmem_n15962), .ZN(MEM_stage_inst_dmem_n15955) );
NAND2_X1 MEM_stage_inst_dmem_U13493 ( .A1(MEM_stage_inst_dmem_n15953), .A2(MEM_stage_inst_dmem_n15952), .ZN(MEM_stage_inst_dmem_n11328) );
NAND2_X1 MEM_stage_inst_dmem_U13492 ( .A1(MEM_stage_inst_dmem_n13059), .A2(MEM_stage_inst_dmem_n15963), .ZN(MEM_stage_inst_dmem_n15952) );
NAND2_X1 MEM_stage_inst_dmem_U13491 ( .A1(MEM_stage_inst_dmem_ram_1029), .A2(MEM_stage_inst_dmem_n15962), .ZN(MEM_stage_inst_dmem_n15953) );
NAND2_X1 MEM_stage_inst_dmem_U13490 ( .A1(MEM_stage_inst_dmem_n15951), .A2(MEM_stage_inst_dmem_n15950), .ZN(MEM_stage_inst_dmem_n11329) );
NAND2_X1 MEM_stage_inst_dmem_U13489 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n15963), .ZN(MEM_stage_inst_dmem_n15950) );
NAND2_X1 MEM_stage_inst_dmem_U13488 ( .A1(MEM_stage_inst_dmem_ram_1030), .A2(MEM_stage_inst_dmem_n15962), .ZN(MEM_stage_inst_dmem_n15951) );
NAND2_X1 MEM_stage_inst_dmem_U13487 ( .A1(MEM_stage_inst_dmem_n15949), .A2(MEM_stage_inst_dmem_n15948), .ZN(MEM_stage_inst_dmem_n11330) );
NAND2_X1 MEM_stage_inst_dmem_U13486 ( .A1(MEM_stage_inst_dmem_n16777), .A2(MEM_stage_inst_dmem_n15963), .ZN(MEM_stage_inst_dmem_n15948) );
NAND2_X1 MEM_stage_inst_dmem_U13485 ( .A1(MEM_stage_inst_dmem_ram_1031), .A2(MEM_stage_inst_dmem_n15962), .ZN(MEM_stage_inst_dmem_n15949) );
NAND2_X1 MEM_stage_inst_dmem_U13484 ( .A1(MEM_stage_inst_dmem_n15947), .A2(MEM_stage_inst_dmem_n15946), .ZN(MEM_stage_inst_dmem_n11331) );
NAND2_X1 MEM_stage_inst_dmem_U13483 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n15963), .ZN(MEM_stage_inst_dmem_n15946) );
NAND2_X1 MEM_stage_inst_dmem_U13482 ( .A1(MEM_stage_inst_dmem_ram_1032), .A2(MEM_stage_inst_dmem_n15962), .ZN(MEM_stage_inst_dmem_n15947) );
NAND2_X1 MEM_stage_inst_dmem_U13481 ( .A1(MEM_stage_inst_dmem_n15945), .A2(MEM_stage_inst_dmem_n15944), .ZN(MEM_stage_inst_dmem_n11332) );
NAND2_X1 MEM_stage_inst_dmem_U13480 ( .A1(MEM_stage_inst_dmem_n16772), .A2(MEM_stage_inst_dmem_n15963), .ZN(MEM_stage_inst_dmem_n15944) );
NAND2_X1 MEM_stage_inst_dmem_U13479 ( .A1(MEM_stage_inst_dmem_ram_1033), .A2(MEM_stage_inst_dmem_n15962), .ZN(MEM_stage_inst_dmem_n15945) );
NAND2_X1 MEM_stage_inst_dmem_U13478 ( .A1(MEM_stage_inst_dmem_n15943), .A2(MEM_stage_inst_dmem_n15942), .ZN(MEM_stage_inst_dmem_n11333) );
NAND2_X1 MEM_stage_inst_dmem_U13477 ( .A1(MEM_stage_inst_dmem_n16769), .A2(MEM_stage_inst_dmem_n15963), .ZN(MEM_stage_inst_dmem_n15942) );
NAND2_X1 MEM_stage_inst_dmem_U13476 ( .A1(MEM_stage_inst_dmem_ram_1034), .A2(MEM_stage_inst_dmem_n15962), .ZN(MEM_stage_inst_dmem_n15943) );
NAND2_X1 MEM_stage_inst_dmem_U13475 ( .A1(MEM_stage_inst_dmem_n15941), .A2(MEM_stage_inst_dmem_n15940), .ZN(MEM_stage_inst_dmem_n11334) );
NAND2_X1 MEM_stage_inst_dmem_U13474 ( .A1(MEM_stage_inst_dmem_n20904), .A2(MEM_stage_inst_dmem_n15963), .ZN(MEM_stage_inst_dmem_n15940) );
NAND2_X1 MEM_stage_inst_dmem_U13473 ( .A1(MEM_stage_inst_dmem_ram_1035), .A2(MEM_stage_inst_dmem_n15962), .ZN(MEM_stage_inst_dmem_n15941) );
NAND2_X1 MEM_stage_inst_dmem_U13472 ( .A1(MEM_stage_inst_dmem_n15939), .A2(MEM_stage_inst_dmem_n15938), .ZN(MEM_stage_inst_dmem_n11335) );
NAND2_X1 MEM_stage_inst_dmem_U13471 ( .A1(MEM_stage_inst_dmem_n21474), .A2(MEM_stage_inst_dmem_n15963), .ZN(MEM_stage_inst_dmem_n15938) );
NAND2_X1 MEM_stage_inst_dmem_U13470 ( .A1(MEM_stage_inst_dmem_ram_1036), .A2(MEM_stage_inst_dmem_n15962), .ZN(MEM_stage_inst_dmem_n15939) );
NAND2_X1 MEM_stage_inst_dmem_U13469 ( .A1(MEM_stage_inst_dmem_n15937), .A2(MEM_stage_inst_dmem_n15936), .ZN(MEM_stage_inst_dmem_n11336) );
NAND2_X1 MEM_stage_inst_dmem_U13468 ( .A1(MEM_stage_inst_dmem_n19242), .A2(MEM_stage_inst_dmem_n15963), .ZN(MEM_stage_inst_dmem_n15936) );
NAND2_X1 MEM_stage_inst_dmem_U13467 ( .A1(MEM_stage_inst_dmem_ram_1037), .A2(MEM_stage_inst_dmem_n15962), .ZN(MEM_stage_inst_dmem_n15937) );
NAND2_X1 MEM_stage_inst_dmem_U13466 ( .A1(MEM_stage_inst_dmem_n15935), .A2(MEM_stage_inst_dmem_n15934), .ZN(MEM_stage_inst_dmem_n11337) );
NAND2_X1 MEM_stage_inst_dmem_U13465 ( .A1(MEM_stage_inst_dmem_n115), .A2(MEM_stage_inst_dmem_n15963), .ZN(MEM_stage_inst_dmem_n15934) );
NAND2_X1 MEM_stage_inst_dmem_U13464 ( .A1(MEM_stage_inst_dmem_ram_1038), .A2(MEM_stage_inst_dmem_n15962), .ZN(MEM_stage_inst_dmem_n15935) );
NAND2_X1 MEM_stage_inst_dmem_U13463 ( .A1(MEM_stage_inst_dmem_n15933), .A2(MEM_stage_inst_dmem_n15932), .ZN(MEM_stage_inst_dmem_n11338) );
NAND2_X1 MEM_stage_inst_dmem_U13462 ( .A1(MEM_stage_inst_dmem_n16758), .A2(MEM_stage_inst_dmem_n15963), .ZN(MEM_stage_inst_dmem_n15932) );
INV_X1 MEM_stage_inst_dmem_U13461 ( .A(MEM_stage_inst_dmem_n15962), .ZN(MEM_stage_inst_dmem_n15963) );
NAND2_X1 MEM_stage_inst_dmem_U13460 ( .A1(MEM_stage_inst_dmem_ram_1039), .A2(MEM_stage_inst_dmem_n15962), .ZN(MEM_stage_inst_dmem_n15933) );
NAND2_X1 MEM_stage_inst_dmem_U13459 ( .A1(MEM_stage_inst_dmem_n21465), .A2(MEM_stage_inst_dmem_n15931), .ZN(MEM_stage_inst_dmem_n15962) );
NAND2_X1 MEM_stage_inst_dmem_U13458 ( .A1(MEM_stage_inst_dmem_n15930), .A2(MEM_stage_inst_dmem_n15929), .ZN(MEM_stage_inst_dmem_n11339) );
NAND2_X1 MEM_stage_inst_dmem_U13457 ( .A1(EX_pipeline_reg_out_5), .A2(MEM_stage_inst_dmem_n15928), .ZN(MEM_stage_inst_dmem_n15929) );
NAND2_X1 MEM_stage_inst_dmem_U13456 ( .A1(MEM_stage_inst_dmem_ram_1040), .A2(MEM_stage_inst_dmem_n15927), .ZN(MEM_stage_inst_dmem_n15930) );
NAND2_X1 MEM_stage_inst_dmem_U13455 ( .A1(MEM_stage_inst_dmem_n15926), .A2(MEM_stage_inst_dmem_n15925), .ZN(MEM_stage_inst_dmem_n11340) );
NAND2_X1 MEM_stage_inst_dmem_U13454 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n15928), .ZN(MEM_stage_inst_dmem_n15925) );
NAND2_X1 MEM_stage_inst_dmem_U13453 ( .A1(MEM_stage_inst_dmem_ram_1041), .A2(MEM_stage_inst_dmem_n15927), .ZN(MEM_stage_inst_dmem_n15926) );
NAND2_X1 MEM_stage_inst_dmem_U13452 ( .A1(MEM_stage_inst_dmem_n15924), .A2(MEM_stage_inst_dmem_n15923), .ZN(MEM_stage_inst_dmem_n11341) );
NAND2_X1 MEM_stage_inst_dmem_U13451 ( .A1(MEM_stage_inst_dmem_n16789), .A2(MEM_stage_inst_dmem_n15928), .ZN(MEM_stage_inst_dmem_n15923) );
NAND2_X1 MEM_stage_inst_dmem_U13450 ( .A1(MEM_stage_inst_dmem_ram_1042), .A2(MEM_stage_inst_dmem_n15927), .ZN(MEM_stage_inst_dmem_n15924) );
NAND2_X1 MEM_stage_inst_dmem_U13449 ( .A1(MEM_stage_inst_dmem_n15922), .A2(MEM_stage_inst_dmem_n15921), .ZN(MEM_stage_inst_dmem_n11342) );
NAND2_X1 MEM_stage_inst_dmem_U13448 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n15928), .ZN(MEM_stage_inst_dmem_n15921) );
NAND2_X1 MEM_stage_inst_dmem_U13447 ( .A1(MEM_stage_inst_dmem_ram_1043), .A2(MEM_stage_inst_dmem_n15927), .ZN(MEM_stage_inst_dmem_n15922) );
NAND2_X1 MEM_stage_inst_dmem_U13446 ( .A1(MEM_stage_inst_dmem_n15920), .A2(MEM_stage_inst_dmem_n15919), .ZN(MEM_stage_inst_dmem_n11343) );
NAND2_X1 MEM_stage_inst_dmem_U13445 ( .A1(MEM_stage_inst_dmem_n16784), .A2(MEM_stage_inst_dmem_n15928), .ZN(MEM_stage_inst_dmem_n15919) );
NAND2_X1 MEM_stage_inst_dmem_U13444 ( .A1(MEM_stage_inst_dmem_ram_1044), .A2(MEM_stage_inst_dmem_n15927), .ZN(MEM_stage_inst_dmem_n15920) );
NAND2_X1 MEM_stage_inst_dmem_U13443 ( .A1(MEM_stage_inst_dmem_n15918), .A2(MEM_stage_inst_dmem_n15917), .ZN(MEM_stage_inst_dmem_n11344) );
NAND2_X1 MEM_stage_inst_dmem_U13442 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n15928), .ZN(MEM_stage_inst_dmem_n15917) );
NAND2_X1 MEM_stage_inst_dmem_U13441 ( .A1(MEM_stage_inst_dmem_ram_1045), .A2(MEM_stage_inst_dmem_n15927), .ZN(MEM_stage_inst_dmem_n15918) );
NAND2_X1 MEM_stage_inst_dmem_U13440 ( .A1(MEM_stage_inst_dmem_n15916), .A2(MEM_stage_inst_dmem_n15915), .ZN(MEM_stage_inst_dmem_n11345) );
NAND2_X1 MEM_stage_inst_dmem_U13439 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n15928), .ZN(MEM_stage_inst_dmem_n15915) );
NAND2_X1 MEM_stage_inst_dmem_U13438 ( .A1(MEM_stage_inst_dmem_ram_1046), .A2(MEM_stage_inst_dmem_n15927), .ZN(MEM_stage_inst_dmem_n15916) );
NAND2_X1 MEM_stage_inst_dmem_U13437 ( .A1(MEM_stage_inst_dmem_n15914), .A2(MEM_stage_inst_dmem_n15913), .ZN(MEM_stage_inst_dmem_n11346) );
NAND2_X1 MEM_stage_inst_dmem_U13436 ( .A1(MEM_stage_inst_dmem_n16777), .A2(MEM_stage_inst_dmem_n15928), .ZN(MEM_stage_inst_dmem_n15913) );
NAND2_X1 MEM_stage_inst_dmem_U13435 ( .A1(MEM_stage_inst_dmem_ram_1047), .A2(MEM_stage_inst_dmem_n15927), .ZN(MEM_stage_inst_dmem_n15914) );
NAND2_X1 MEM_stage_inst_dmem_U13434 ( .A1(MEM_stage_inst_dmem_n15912), .A2(MEM_stage_inst_dmem_n15911), .ZN(MEM_stage_inst_dmem_n11347) );
NAND2_X1 MEM_stage_inst_dmem_U13433 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n15928), .ZN(MEM_stage_inst_dmem_n15911) );
NAND2_X1 MEM_stage_inst_dmem_U13432 ( .A1(MEM_stage_inst_dmem_ram_1048), .A2(MEM_stage_inst_dmem_n15927), .ZN(MEM_stage_inst_dmem_n15912) );
NAND2_X1 MEM_stage_inst_dmem_U13431 ( .A1(MEM_stage_inst_dmem_n15910), .A2(MEM_stage_inst_dmem_n15909), .ZN(MEM_stage_inst_dmem_n11348) );
NAND2_X1 MEM_stage_inst_dmem_U13430 ( .A1(MEM_stage_inst_dmem_n16772), .A2(MEM_stage_inst_dmem_n15928), .ZN(MEM_stage_inst_dmem_n15909) );
NAND2_X1 MEM_stage_inst_dmem_U13429 ( .A1(MEM_stage_inst_dmem_ram_1049), .A2(MEM_stage_inst_dmem_n15927), .ZN(MEM_stage_inst_dmem_n15910) );
NAND2_X1 MEM_stage_inst_dmem_U13428 ( .A1(MEM_stage_inst_dmem_n15908), .A2(MEM_stage_inst_dmem_n15907), .ZN(MEM_stage_inst_dmem_n11349) );
NAND2_X1 MEM_stage_inst_dmem_U13427 ( .A1(MEM_stage_inst_dmem_n16769), .A2(MEM_stage_inst_dmem_n15928), .ZN(MEM_stage_inst_dmem_n15907) );
NAND2_X1 MEM_stage_inst_dmem_U13426 ( .A1(MEM_stage_inst_dmem_ram_1050), .A2(MEM_stage_inst_dmem_n15927), .ZN(MEM_stage_inst_dmem_n15908) );
NAND2_X1 MEM_stage_inst_dmem_U13425 ( .A1(MEM_stage_inst_dmem_n15906), .A2(MEM_stage_inst_dmem_n15905), .ZN(MEM_stage_inst_dmem_n11350) );
NAND2_X1 MEM_stage_inst_dmem_U13424 ( .A1(MEM_stage_inst_dmem_n20518), .A2(MEM_stage_inst_dmem_n15928), .ZN(MEM_stage_inst_dmem_n15905) );
NAND2_X1 MEM_stage_inst_dmem_U13423 ( .A1(MEM_stage_inst_dmem_ram_1051), .A2(MEM_stage_inst_dmem_n15927), .ZN(MEM_stage_inst_dmem_n15906) );
NAND2_X1 MEM_stage_inst_dmem_U13422 ( .A1(MEM_stage_inst_dmem_n15904), .A2(MEM_stage_inst_dmem_n15903), .ZN(MEM_stage_inst_dmem_n11351) );
NAND2_X1 MEM_stage_inst_dmem_U13421 ( .A1(MEM_stage_inst_dmem_n20515), .A2(MEM_stage_inst_dmem_n15928), .ZN(MEM_stage_inst_dmem_n15903) );
NAND2_X1 MEM_stage_inst_dmem_U13420 ( .A1(MEM_stage_inst_dmem_ram_1052), .A2(MEM_stage_inst_dmem_n15927), .ZN(MEM_stage_inst_dmem_n15904) );
NAND2_X1 MEM_stage_inst_dmem_U13419 ( .A1(MEM_stage_inst_dmem_n15902), .A2(MEM_stage_inst_dmem_n15901), .ZN(MEM_stage_inst_dmem_n11352) );
NAND2_X1 MEM_stage_inst_dmem_U13418 ( .A1(EX_pipeline_reg_out_18), .A2(MEM_stage_inst_dmem_n15928), .ZN(MEM_stage_inst_dmem_n15901) );
NAND2_X1 MEM_stage_inst_dmem_U13417 ( .A1(MEM_stage_inst_dmem_ram_1053), .A2(MEM_stage_inst_dmem_n15927), .ZN(MEM_stage_inst_dmem_n15902) );
NAND2_X1 MEM_stage_inst_dmem_U13416 ( .A1(MEM_stage_inst_dmem_n15900), .A2(MEM_stage_inst_dmem_n15899), .ZN(MEM_stage_inst_dmem_n11353) );
NAND2_X1 MEM_stage_inst_dmem_U13415 ( .A1(EX_pipeline_reg_out_19), .A2(MEM_stage_inst_dmem_n15928), .ZN(MEM_stage_inst_dmem_n15899) );
NAND2_X1 MEM_stage_inst_dmem_U13414 ( .A1(MEM_stage_inst_dmem_ram_1054), .A2(MEM_stage_inst_dmem_n15927), .ZN(MEM_stage_inst_dmem_n15900) );
NAND2_X1 MEM_stage_inst_dmem_U13413 ( .A1(MEM_stage_inst_dmem_n15898), .A2(MEM_stage_inst_dmem_n15897), .ZN(MEM_stage_inst_dmem_n11354) );
NAND2_X1 MEM_stage_inst_dmem_U13412 ( .A1(MEM_stage_inst_dmem_n16758), .A2(MEM_stage_inst_dmem_n15928), .ZN(MEM_stage_inst_dmem_n15897) );
INV_X1 MEM_stage_inst_dmem_U13411 ( .A(MEM_stage_inst_dmem_n15927), .ZN(MEM_stage_inst_dmem_n15928) );
NAND2_X1 MEM_stage_inst_dmem_U13410 ( .A1(MEM_stage_inst_dmem_ram_1055), .A2(MEM_stage_inst_dmem_n15927), .ZN(MEM_stage_inst_dmem_n15898) );
NAND2_X1 MEM_stage_inst_dmem_U13409 ( .A1(MEM_stage_inst_dmem_n21429), .A2(MEM_stage_inst_dmem_n15931), .ZN(MEM_stage_inst_dmem_n15927) );
NAND2_X1 MEM_stage_inst_dmem_U13408 ( .A1(MEM_stage_inst_dmem_n15896), .A2(MEM_stage_inst_dmem_n15895), .ZN(MEM_stage_inst_dmem_n11355) );
NAND2_X1 MEM_stage_inst_dmem_U13407 ( .A1(MEM_stage_inst_dmem_n14732), .A2(MEM_stage_inst_dmem_n15894), .ZN(MEM_stage_inst_dmem_n15895) );
NAND2_X1 MEM_stage_inst_dmem_U13406 ( .A1(MEM_stage_inst_dmem_ram_1056), .A2(MEM_stage_inst_dmem_n15893), .ZN(MEM_stage_inst_dmem_n15896) );
NAND2_X1 MEM_stage_inst_dmem_U13405 ( .A1(MEM_stage_inst_dmem_n15892), .A2(MEM_stage_inst_dmem_n15891), .ZN(MEM_stage_inst_dmem_n11356) );
NAND2_X1 MEM_stage_inst_dmem_U13404 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n15894), .ZN(MEM_stage_inst_dmem_n15891) );
NAND2_X1 MEM_stage_inst_dmem_U13403 ( .A1(MEM_stage_inst_dmem_ram_1057), .A2(MEM_stage_inst_dmem_n15893), .ZN(MEM_stage_inst_dmem_n15892) );
NAND2_X1 MEM_stage_inst_dmem_U13402 ( .A1(MEM_stage_inst_dmem_n15890), .A2(MEM_stage_inst_dmem_n15889), .ZN(MEM_stage_inst_dmem_n11357) );
NAND2_X1 MEM_stage_inst_dmem_U13401 ( .A1(MEM_stage_inst_dmem_n16789), .A2(MEM_stage_inst_dmem_n15894), .ZN(MEM_stage_inst_dmem_n15889) );
NAND2_X1 MEM_stage_inst_dmem_U13400 ( .A1(MEM_stage_inst_dmem_ram_1058), .A2(MEM_stage_inst_dmem_n15893), .ZN(MEM_stage_inst_dmem_n15890) );
NAND2_X1 MEM_stage_inst_dmem_U13399 ( .A1(MEM_stage_inst_dmem_n15888), .A2(MEM_stage_inst_dmem_n15887), .ZN(MEM_stage_inst_dmem_n11358) );
NAND2_X1 MEM_stage_inst_dmem_U13398 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n15894), .ZN(MEM_stage_inst_dmem_n15887) );
NAND2_X1 MEM_stage_inst_dmem_U13397 ( .A1(MEM_stage_inst_dmem_ram_1059), .A2(MEM_stage_inst_dmem_n15893), .ZN(MEM_stage_inst_dmem_n15888) );
NAND2_X1 MEM_stage_inst_dmem_U13396 ( .A1(MEM_stage_inst_dmem_n15886), .A2(MEM_stage_inst_dmem_n15885), .ZN(MEM_stage_inst_dmem_n11359) );
NAND2_X1 MEM_stage_inst_dmem_U13395 ( .A1(MEM_stage_inst_dmem_n16784), .A2(MEM_stage_inst_dmem_n15894), .ZN(MEM_stage_inst_dmem_n15885) );
NAND2_X1 MEM_stage_inst_dmem_U13394 ( .A1(MEM_stage_inst_dmem_ram_1060), .A2(MEM_stage_inst_dmem_n15893), .ZN(MEM_stage_inst_dmem_n15886) );
NAND2_X1 MEM_stage_inst_dmem_U13393 ( .A1(MEM_stage_inst_dmem_n15884), .A2(MEM_stage_inst_dmem_n15883), .ZN(MEM_stage_inst_dmem_n11360) );
NAND2_X1 MEM_stage_inst_dmem_U13392 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n15894), .ZN(MEM_stage_inst_dmem_n15883) );
NAND2_X1 MEM_stage_inst_dmem_U13391 ( .A1(MEM_stage_inst_dmem_ram_1061), .A2(MEM_stage_inst_dmem_n15893), .ZN(MEM_stage_inst_dmem_n15884) );
NAND2_X1 MEM_stage_inst_dmem_U13390 ( .A1(MEM_stage_inst_dmem_n15882), .A2(MEM_stage_inst_dmem_n15881), .ZN(MEM_stage_inst_dmem_n11361) );
NAND2_X1 MEM_stage_inst_dmem_U13389 ( .A1(MEM_stage_inst_dmem_n13056), .A2(MEM_stage_inst_dmem_n15894), .ZN(MEM_stage_inst_dmem_n15881) );
NAND2_X1 MEM_stage_inst_dmem_U13388 ( .A1(MEM_stage_inst_dmem_ram_1062), .A2(MEM_stage_inst_dmem_n15893), .ZN(MEM_stage_inst_dmem_n15882) );
NAND2_X1 MEM_stage_inst_dmem_U13387 ( .A1(MEM_stage_inst_dmem_n15880), .A2(MEM_stage_inst_dmem_n15879), .ZN(MEM_stage_inst_dmem_n11362) );
NAND2_X1 MEM_stage_inst_dmem_U13386 ( .A1(MEM_stage_inst_dmem_n16777), .A2(MEM_stage_inst_dmem_n15894), .ZN(MEM_stage_inst_dmem_n15879) );
NAND2_X1 MEM_stage_inst_dmem_U13385 ( .A1(MEM_stage_inst_dmem_ram_1063), .A2(MEM_stage_inst_dmem_n15893), .ZN(MEM_stage_inst_dmem_n15880) );
NAND2_X1 MEM_stage_inst_dmem_U13384 ( .A1(MEM_stage_inst_dmem_n15878), .A2(MEM_stage_inst_dmem_n15877), .ZN(MEM_stage_inst_dmem_n11363) );
NAND2_X1 MEM_stage_inst_dmem_U13383 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n15894), .ZN(MEM_stage_inst_dmem_n15877) );
NAND2_X1 MEM_stage_inst_dmem_U13382 ( .A1(MEM_stage_inst_dmem_ram_1064), .A2(MEM_stage_inst_dmem_n15893), .ZN(MEM_stage_inst_dmem_n15878) );
NAND2_X1 MEM_stage_inst_dmem_U13381 ( .A1(MEM_stage_inst_dmem_n15876), .A2(MEM_stage_inst_dmem_n15875), .ZN(MEM_stage_inst_dmem_n11364) );
NAND2_X1 MEM_stage_inst_dmem_U13380 ( .A1(MEM_stage_inst_dmem_n16772), .A2(MEM_stage_inst_dmem_n15894), .ZN(MEM_stage_inst_dmem_n15875) );
NAND2_X1 MEM_stage_inst_dmem_U13379 ( .A1(MEM_stage_inst_dmem_ram_1065), .A2(MEM_stage_inst_dmem_n15893), .ZN(MEM_stage_inst_dmem_n15876) );
NAND2_X1 MEM_stage_inst_dmem_U13378 ( .A1(MEM_stage_inst_dmem_n15874), .A2(MEM_stage_inst_dmem_n15873), .ZN(MEM_stage_inst_dmem_n11365) );
NAND2_X1 MEM_stage_inst_dmem_U13377 ( .A1(MEM_stage_inst_dmem_n16769), .A2(MEM_stage_inst_dmem_n15894), .ZN(MEM_stage_inst_dmem_n15873) );
NAND2_X1 MEM_stage_inst_dmem_U13376 ( .A1(MEM_stage_inst_dmem_ram_1066), .A2(MEM_stage_inst_dmem_n15893), .ZN(MEM_stage_inst_dmem_n15874) );
NAND2_X1 MEM_stage_inst_dmem_U13375 ( .A1(MEM_stage_inst_dmem_n15872), .A2(MEM_stage_inst_dmem_n15871), .ZN(MEM_stage_inst_dmem_n11366) );
NAND2_X1 MEM_stage_inst_dmem_U13374 ( .A1(MEM_stage_inst_dmem_n13044), .A2(MEM_stage_inst_dmem_n15894), .ZN(MEM_stage_inst_dmem_n15871) );
NAND2_X1 MEM_stage_inst_dmem_U13373 ( .A1(MEM_stage_inst_dmem_ram_1067), .A2(MEM_stage_inst_dmem_n15893), .ZN(MEM_stage_inst_dmem_n15872) );
NAND2_X1 MEM_stage_inst_dmem_U13372 ( .A1(MEM_stage_inst_dmem_n15870), .A2(MEM_stage_inst_dmem_n15869), .ZN(MEM_stage_inst_dmem_n11367) );
NAND2_X1 MEM_stage_inst_dmem_U13371 ( .A1(MEM_stage_inst_dmem_n13041), .A2(MEM_stage_inst_dmem_n15894), .ZN(MEM_stage_inst_dmem_n15869) );
NAND2_X1 MEM_stage_inst_dmem_U13370 ( .A1(MEM_stage_inst_dmem_ram_1068), .A2(MEM_stage_inst_dmem_n15893), .ZN(MEM_stage_inst_dmem_n15870) );
NAND2_X1 MEM_stage_inst_dmem_U13369 ( .A1(MEM_stage_inst_dmem_n15868), .A2(MEM_stage_inst_dmem_n15867), .ZN(MEM_stage_inst_dmem_n11368) );
NAND2_X1 MEM_stage_inst_dmem_U13368 ( .A1(MEM_stage_inst_dmem_n116), .A2(MEM_stage_inst_dmem_n15894), .ZN(MEM_stage_inst_dmem_n15867) );
NAND2_X1 MEM_stage_inst_dmem_U13367 ( .A1(MEM_stage_inst_dmem_ram_1069), .A2(MEM_stage_inst_dmem_n15893), .ZN(MEM_stage_inst_dmem_n15868) );
NAND2_X1 MEM_stage_inst_dmem_U13366 ( .A1(MEM_stage_inst_dmem_n15866), .A2(MEM_stage_inst_dmem_n15865), .ZN(MEM_stage_inst_dmem_n11369) );
NAND2_X1 MEM_stage_inst_dmem_U13365 ( .A1(MEM_stage_inst_dmem_n14696), .A2(MEM_stage_inst_dmem_n15894), .ZN(MEM_stage_inst_dmem_n15865) );
NAND2_X1 MEM_stage_inst_dmem_U13364 ( .A1(MEM_stage_inst_dmem_ram_1070), .A2(MEM_stage_inst_dmem_n15893), .ZN(MEM_stage_inst_dmem_n15866) );
NAND2_X1 MEM_stage_inst_dmem_U13363 ( .A1(MEM_stage_inst_dmem_n15864), .A2(MEM_stage_inst_dmem_n15863), .ZN(MEM_stage_inst_dmem_n11370) );
NAND2_X1 MEM_stage_inst_dmem_U13362 ( .A1(MEM_stage_inst_dmem_n16758), .A2(MEM_stage_inst_dmem_n15894), .ZN(MEM_stage_inst_dmem_n15863) );
NAND2_X1 MEM_stage_inst_dmem_U13361 ( .A1(MEM_stage_inst_dmem_ram_1071), .A2(MEM_stage_inst_dmem_n15893), .ZN(MEM_stage_inst_dmem_n15864) );
NAND2_X1 MEM_stage_inst_dmem_U13360 ( .A1(MEM_stage_inst_dmem_n21394), .A2(MEM_stage_inst_dmem_n15931), .ZN(MEM_stage_inst_dmem_n15893) );
NAND2_X1 MEM_stage_inst_dmem_U13359 ( .A1(MEM_stage_inst_dmem_n15862), .A2(MEM_stage_inst_dmem_n15861), .ZN(MEM_stage_inst_dmem_n11371) );
NAND2_X1 MEM_stage_inst_dmem_U13358 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n15860), .ZN(MEM_stage_inst_dmem_n15861) );
NAND2_X1 MEM_stage_inst_dmem_U13357 ( .A1(MEM_stage_inst_dmem_ram_1072), .A2(MEM_stage_inst_dmem_n15859), .ZN(MEM_stage_inst_dmem_n15862) );
NAND2_X1 MEM_stage_inst_dmem_U13356 ( .A1(MEM_stage_inst_dmem_n15858), .A2(MEM_stage_inst_dmem_n15857), .ZN(MEM_stage_inst_dmem_n11372) );
NAND2_X1 MEM_stage_inst_dmem_U13355 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n15860), .ZN(MEM_stage_inst_dmem_n15857) );
NAND2_X1 MEM_stage_inst_dmem_U13354 ( .A1(MEM_stage_inst_dmem_ram_1073), .A2(MEM_stage_inst_dmem_n15859), .ZN(MEM_stage_inst_dmem_n15858) );
NAND2_X1 MEM_stage_inst_dmem_U13353 ( .A1(MEM_stage_inst_dmem_n15856), .A2(MEM_stage_inst_dmem_n15855), .ZN(MEM_stage_inst_dmem_n11373) );
NAND2_X1 MEM_stage_inst_dmem_U13352 ( .A1(MEM_stage_inst_dmem_n16789), .A2(MEM_stage_inst_dmem_n15860), .ZN(MEM_stage_inst_dmem_n15855) );
NAND2_X1 MEM_stage_inst_dmem_U13351 ( .A1(MEM_stage_inst_dmem_ram_1074), .A2(MEM_stage_inst_dmem_n15859), .ZN(MEM_stage_inst_dmem_n15856) );
NAND2_X1 MEM_stage_inst_dmem_U13350 ( .A1(MEM_stage_inst_dmem_n15854), .A2(MEM_stage_inst_dmem_n15853), .ZN(MEM_stage_inst_dmem_n11374) );
NAND2_X1 MEM_stage_inst_dmem_U13349 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n15860), .ZN(MEM_stage_inst_dmem_n15853) );
NAND2_X1 MEM_stage_inst_dmem_U13348 ( .A1(MEM_stage_inst_dmem_ram_1075), .A2(MEM_stage_inst_dmem_n15859), .ZN(MEM_stage_inst_dmem_n15854) );
NAND2_X1 MEM_stage_inst_dmem_U13347 ( .A1(MEM_stage_inst_dmem_n15852), .A2(MEM_stage_inst_dmem_n15851), .ZN(MEM_stage_inst_dmem_n11375) );
NAND2_X1 MEM_stage_inst_dmem_U13346 ( .A1(MEM_stage_inst_dmem_n16784), .A2(MEM_stage_inst_dmem_n15860), .ZN(MEM_stage_inst_dmem_n15851) );
NAND2_X1 MEM_stage_inst_dmem_U13345 ( .A1(MEM_stage_inst_dmem_ram_1076), .A2(MEM_stage_inst_dmem_n15859), .ZN(MEM_stage_inst_dmem_n15852) );
NAND2_X1 MEM_stage_inst_dmem_U13344 ( .A1(MEM_stage_inst_dmem_n15850), .A2(MEM_stage_inst_dmem_n15849), .ZN(MEM_stage_inst_dmem_n11376) );
NAND2_X1 MEM_stage_inst_dmem_U13343 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n15860), .ZN(MEM_stage_inst_dmem_n15849) );
NAND2_X1 MEM_stage_inst_dmem_U13342 ( .A1(MEM_stage_inst_dmem_ram_1077), .A2(MEM_stage_inst_dmem_n15859), .ZN(MEM_stage_inst_dmem_n15850) );
NAND2_X1 MEM_stage_inst_dmem_U13341 ( .A1(MEM_stage_inst_dmem_n15848), .A2(MEM_stage_inst_dmem_n15847), .ZN(MEM_stage_inst_dmem_n11377) );
NAND2_X1 MEM_stage_inst_dmem_U13340 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n15860), .ZN(MEM_stage_inst_dmem_n15847) );
NAND2_X1 MEM_stage_inst_dmem_U13339 ( .A1(MEM_stage_inst_dmem_ram_1078), .A2(MEM_stage_inst_dmem_n15859), .ZN(MEM_stage_inst_dmem_n15848) );
NAND2_X1 MEM_stage_inst_dmem_U13338 ( .A1(MEM_stage_inst_dmem_n15846), .A2(MEM_stage_inst_dmem_n15845), .ZN(MEM_stage_inst_dmem_n11378) );
NAND2_X1 MEM_stage_inst_dmem_U13337 ( .A1(MEM_stage_inst_dmem_n16777), .A2(MEM_stage_inst_dmem_n15860), .ZN(MEM_stage_inst_dmem_n15845) );
NAND2_X1 MEM_stage_inst_dmem_U13336 ( .A1(MEM_stage_inst_dmem_ram_1079), .A2(MEM_stage_inst_dmem_n15859), .ZN(MEM_stage_inst_dmem_n15846) );
NAND2_X1 MEM_stage_inst_dmem_U13335 ( .A1(MEM_stage_inst_dmem_n15844), .A2(MEM_stage_inst_dmem_n15843), .ZN(MEM_stage_inst_dmem_n11379) );
NAND2_X1 MEM_stage_inst_dmem_U13334 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n15860), .ZN(MEM_stage_inst_dmem_n15843) );
NAND2_X1 MEM_stage_inst_dmem_U13333 ( .A1(MEM_stage_inst_dmem_ram_1080), .A2(MEM_stage_inst_dmem_n15859), .ZN(MEM_stage_inst_dmem_n15844) );
NAND2_X1 MEM_stage_inst_dmem_U13332 ( .A1(MEM_stage_inst_dmem_n15842), .A2(MEM_stage_inst_dmem_n15841), .ZN(MEM_stage_inst_dmem_n11380) );
NAND2_X1 MEM_stage_inst_dmem_U13331 ( .A1(MEM_stage_inst_dmem_n16772), .A2(MEM_stage_inst_dmem_n15860), .ZN(MEM_stage_inst_dmem_n15841) );
NAND2_X1 MEM_stage_inst_dmem_U13330 ( .A1(MEM_stage_inst_dmem_ram_1081), .A2(MEM_stage_inst_dmem_n15859), .ZN(MEM_stage_inst_dmem_n15842) );
NAND2_X1 MEM_stage_inst_dmem_U13329 ( .A1(MEM_stage_inst_dmem_n15840), .A2(MEM_stage_inst_dmem_n15839), .ZN(MEM_stage_inst_dmem_n11381) );
NAND2_X1 MEM_stage_inst_dmem_U13328 ( .A1(MEM_stage_inst_dmem_n16769), .A2(MEM_stage_inst_dmem_n15860), .ZN(MEM_stage_inst_dmem_n15839) );
NAND2_X1 MEM_stage_inst_dmem_U13327 ( .A1(MEM_stage_inst_dmem_ram_1082), .A2(MEM_stage_inst_dmem_n15859), .ZN(MEM_stage_inst_dmem_n15840) );
NAND2_X1 MEM_stage_inst_dmem_U13326 ( .A1(MEM_stage_inst_dmem_n15838), .A2(MEM_stage_inst_dmem_n15837), .ZN(MEM_stage_inst_dmem_n11382) );
NAND2_X1 MEM_stage_inst_dmem_U13325 ( .A1(MEM_stage_inst_dmem_n20904), .A2(MEM_stage_inst_dmem_n15860), .ZN(MEM_stage_inst_dmem_n15837) );
NAND2_X1 MEM_stage_inst_dmem_U13324 ( .A1(MEM_stage_inst_dmem_ram_1083), .A2(MEM_stage_inst_dmem_n15859), .ZN(MEM_stage_inst_dmem_n15838) );
NAND2_X1 MEM_stage_inst_dmem_U13323 ( .A1(MEM_stage_inst_dmem_n15836), .A2(MEM_stage_inst_dmem_n15835), .ZN(MEM_stage_inst_dmem_n11383) );
NAND2_X1 MEM_stage_inst_dmem_U13322 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n15860), .ZN(MEM_stage_inst_dmem_n15835) );
NAND2_X1 MEM_stage_inst_dmem_U13321 ( .A1(MEM_stage_inst_dmem_ram_1084), .A2(MEM_stage_inst_dmem_n15859), .ZN(MEM_stage_inst_dmem_n15836) );
NAND2_X1 MEM_stage_inst_dmem_U13320 ( .A1(MEM_stage_inst_dmem_n15834), .A2(MEM_stage_inst_dmem_n15833), .ZN(MEM_stage_inst_dmem_n11384) );
NAND2_X1 MEM_stage_inst_dmem_U13319 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n15860), .ZN(MEM_stage_inst_dmem_n15833) );
NAND2_X1 MEM_stage_inst_dmem_U13318 ( .A1(MEM_stage_inst_dmem_ram_1085), .A2(MEM_stage_inst_dmem_n15859), .ZN(MEM_stage_inst_dmem_n15834) );
NAND2_X1 MEM_stage_inst_dmem_U13317 ( .A1(MEM_stage_inst_dmem_n15832), .A2(MEM_stage_inst_dmem_n15831), .ZN(MEM_stage_inst_dmem_n11385) );
NAND2_X1 MEM_stage_inst_dmem_U13316 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n15860), .ZN(MEM_stage_inst_dmem_n15831) );
NAND2_X1 MEM_stage_inst_dmem_U13315 ( .A1(MEM_stage_inst_dmem_ram_1086), .A2(MEM_stage_inst_dmem_n15859), .ZN(MEM_stage_inst_dmem_n15832) );
NAND2_X1 MEM_stage_inst_dmem_U13314 ( .A1(MEM_stage_inst_dmem_n15830), .A2(MEM_stage_inst_dmem_n15829), .ZN(MEM_stage_inst_dmem_n11386) );
NAND2_X1 MEM_stage_inst_dmem_U13313 ( .A1(MEM_stage_inst_dmem_n16758), .A2(MEM_stage_inst_dmem_n15860), .ZN(MEM_stage_inst_dmem_n15829) );
INV_X1 MEM_stage_inst_dmem_U13312 ( .A(MEM_stage_inst_dmem_n15859), .ZN(MEM_stage_inst_dmem_n15860) );
NAND2_X1 MEM_stage_inst_dmem_U13311 ( .A1(MEM_stage_inst_dmem_ram_1087), .A2(MEM_stage_inst_dmem_n15859), .ZN(MEM_stage_inst_dmem_n15830) );
NAND2_X1 MEM_stage_inst_dmem_U13310 ( .A1(MEM_stage_inst_dmem_n21359), .A2(MEM_stage_inst_dmem_n15931), .ZN(MEM_stage_inst_dmem_n15859) );
NAND2_X1 MEM_stage_inst_dmem_U13309 ( .A1(MEM_stage_inst_dmem_n15828), .A2(MEM_stage_inst_dmem_n15827), .ZN(MEM_stage_inst_dmem_n11387) );
NAND2_X1 MEM_stage_inst_dmem_U13308 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n15826), .ZN(MEM_stage_inst_dmem_n15827) );
NAND2_X1 MEM_stage_inst_dmem_U13307 ( .A1(MEM_stage_inst_dmem_ram_1088), .A2(MEM_stage_inst_dmem_n15825), .ZN(MEM_stage_inst_dmem_n15828) );
NAND2_X1 MEM_stage_inst_dmem_U13306 ( .A1(MEM_stage_inst_dmem_n15824), .A2(MEM_stage_inst_dmem_n15823), .ZN(MEM_stage_inst_dmem_n11388) );
NAND2_X1 MEM_stage_inst_dmem_U13305 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n15826), .ZN(MEM_stage_inst_dmem_n15823) );
NAND2_X1 MEM_stage_inst_dmem_U13304 ( .A1(MEM_stage_inst_dmem_ram_1089), .A2(MEM_stage_inst_dmem_n15825), .ZN(MEM_stage_inst_dmem_n15824) );
NAND2_X1 MEM_stage_inst_dmem_U13303 ( .A1(MEM_stage_inst_dmem_n15822), .A2(MEM_stage_inst_dmem_n15821), .ZN(MEM_stage_inst_dmem_n11389) );
NAND2_X1 MEM_stage_inst_dmem_U13302 ( .A1(MEM_stage_inst_dmem_n16789), .A2(MEM_stage_inst_dmem_n15826), .ZN(MEM_stage_inst_dmem_n15821) );
NAND2_X1 MEM_stage_inst_dmem_U13301 ( .A1(MEM_stage_inst_dmem_ram_1090), .A2(MEM_stage_inst_dmem_n15825), .ZN(MEM_stage_inst_dmem_n15822) );
NAND2_X1 MEM_stage_inst_dmem_U13300 ( .A1(MEM_stage_inst_dmem_n15820), .A2(MEM_stage_inst_dmem_n15819), .ZN(MEM_stage_inst_dmem_n11390) );
NAND2_X1 MEM_stage_inst_dmem_U13299 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n15826), .ZN(MEM_stage_inst_dmem_n15819) );
NAND2_X1 MEM_stage_inst_dmem_U13298 ( .A1(MEM_stage_inst_dmem_ram_1091), .A2(MEM_stage_inst_dmem_n15825), .ZN(MEM_stage_inst_dmem_n15820) );
NAND2_X1 MEM_stage_inst_dmem_U13297 ( .A1(MEM_stage_inst_dmem_n15818), .A2(MEM_stage_inst_dmem_n15817), .ZN(MEM_stage_inst_dmem_n11391) );
NAND2_X1 MEM_stage_inst_dmem_U13296 ( .A1(MEM_stage_inst_dmem_n16784), .A2(MEM_stage_inst_dmem_n15826), .ZN(MEM_stage_inst_dmem_n15817) );
NAND2_X1 MEM_stage_inst_dmem_U13295 ( .A1(MEM_stage_inst_dmem_ram_1092), .A2(MEM_stage_inst_dmem_n15825), .ZN(MEM_stage_inst_dmem_n15818) );
NAND2_X1 MEM_stage_inst_dmem_U13294 ( .A1(MEM_stage_inst_dmem_n15816), .A2(MEM_stage_inst_dmem_n15815), .ZN(MEM_stage_inst_dmem_n11392) );
NAND2_X1 MEM_stage_inst_dmem_U13293 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n15826), .ZN(MEM_stage_inst_dmem_n15815) );
NAND2_X1 MEM_stage_inst_dmem_U13292 ( .A1(MEM_stage_inst_dmem_ram_1093), .A2(MEM_stage_inst_dmem_n15825), .ZN(MEM_stage_inst_dmem_n15816) );
NAND2_X1 MEM_stage_inst_dmem_U13291 ( .A1(MEM_stage_inst_dmem_n15814), .A2(MEM_stage_inst_dmem_n15813), .ZN(MEM_stage_inst_dmem_n11393) );
NAND2_X1 MEM_stage_inst_dmem_U13290 ( .A1(MEM_stage_inst_dmem_n13056), .A2(MEM_stage_inst_dmem_n15826), .ZN(MEM_stage_inst_dmem_n15813) );
NAND2_X1 MEM_stage_inst_dmem_U13289 ( .A1(MEM_stage_inst_dmem_ram_1094), .A2(MEM_stage_inst_dmem_n15825), .ZN(MEM_stage_inst_dmem_n15814) );
NAND2_X1 MEM_stage_inst_dmem_U13288 ( .A1(MEM_stage_inst_dmem_n15812), .A2(MEM_stage_inst_dmem_n15811), .ZN(MEM_stage_inst_dmem_n11394) );
NAND2_X1 MEM_stage_inst_dmem_U13287 ( .A1(MEM_stage_inst_dmem_n16777), .A2(MEM_stage_inst_dmem_n15826), .ZN(MEM_stage_inst_dmem_n15811) );
NAND2_X1 MEM_stage_inst_dmem_U13286 ( .A1(MEM_stage_inst_dmem_ram_1095), .A2(MEM_stage_inst_dmem_n15825), .ZN(MEM_stage_inst_dmem_n15812) );
NAND2_X1 MEM_stage_inst_dmem_U13285 ( .A1(MEM_stage_inst_dmem_n15810), .A2(MEM_stage_inst_dmem_n15809), .ZN(MEM_stage_inst_dmem_n11395) );
NAND2_X1 MEM_stage_inst_dmem_U13284 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n15826), .ZN(MEM_stage_inst_dmem_n15809) );
NAND2_X1 MEM_stage_inst_dmem_U13283 ( .A1(MEM_stage_inst_dmem_ram_1096), .A2(MEM_stage_inst_dmem_n15825), .ZN(MEM_stage_inst_dmem_n15810) );
NAND2_X1 MEM_stage_inst_dmem_U13282 ( .A1(MEM_stage_inst_dmem_n15808), .A2(MEM_stage_inst_dmem_n15807), .ZN(MEM_stage_inst_dmem_n11396) );
NAND2_X1 MEM_stage_inst_dmem_U13281 ( .A1(MEM_stage_inst_dmem_n16772), .A2(MEM_stage_inst_dmem_n15826), .ZN(MEM_stage_inst_dmem_n15807) );
NAND2_X1 MEM_stage_inst_dmem_U13280 ( .A1(MEM_stage_inst_dmem_ram_1097), .A2(MEM_stage_inst_dmem_n15825), .ZN(MEM_stage_inst_dmem_n15808) );
NAND2_X1 MEM_stage_inst_dmem_U13279 ( .A1(MEM_stage_inst_dmem_n15806), .A2(MEM_stage_inst_dmem_n15805), .ZN(MEM_stage_inst_dmem_n11397) );
NAND2_X1 MEM_stage_inst_dmem_U13278 ( .A1(MEM_stage_inst_dmem_n16769), .A2(MEM_stage_inst_dmem_n15826), .ZN(MEM_stage_inst_dmem_n15805) );
NAND2_X1 MEM_stage_inst_dmem_U13277 ( .A1(MEM_stage_inst_dmem_ram_1098), .A2(MEM_stage_inst_dmem_n15825), .ZN(MEM_stage_inst_dmem_n15806) );
NAND2_X1 MEM_stage_inst_dmem_U13276 ( .A1(MEM_stage_inst_dmem_n15804), .A2(MEM_stage_inst_dmem_n15803), .ZN(MEM_stage_inst_dmem_n11398) );
NAND2_X1 MEM_stage_inst_dmem_U13275 ( .A1(MEM_stage_inst_dmem_n14705), .A2(MEM_stage_inst_dmem_n15826), .ZN(MEM_stage_inst_dmem_n15803) );
NAND2_X1 MEM_stage_inst_dmem_U13274 ( .A1(MEM_stage_inst_dmem_ram_1099), .A2(MEM_stage_inst_dmem_n15825), .ZN(MEM_stage_inst_dmem_n15804) );
NAND2_X1 MEM_stage_inst_dmem_U13273 ( .A1(MEM_stage_inst_dmem_n15802), .A2(MEM_stage_inst_dmem_n15801), .ZN(MEM_stage_inst_dmem_n11399) );
NAND2_X1 MEM_stage_inst_dmem_U13272 ( .A1(MEM_stage_inst_dmem_n14702), .A2(MEM_stage_inst_dmem_n15826), .ZN(MEM_stage_inst_dmem_n15801) );
NAND2_X1 MEM_stage_inst_dmem_U13271 ( .A1(MEM_stage_inst_dmem_ram_1100), .A2(MEM_stage_inst_dmem_n15825), .ZN(MEM_stage_inst_dmem_n15802) );
NAND2_X1 MEM_stage_inst_dmem_U13270 ( .A1(MEM_stage_inst_dmem_n15800), .A2(MEM_stage_inst_dmem_n15799), .ZN(MEM_stage_inst_dmem_n11400) );
NAND2_X1 MEM_stage_inst_dmem_U13269 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n15826), .ZN(MEM_stage_inst_dmem_n15799) );
NAND2_X1 MEM_stage_inst_dmem_U13268 ( .A1(MEM_stage_inst_dmem_ram_1101), .A2(MEM_stage_inst_dmem_n15825), .ZN(MEM_stage_inst_dmem_n15800) );
NAND2_X1 MEM_stage_inst_dmem_U13267 ( .A1(MEM_stage_inst_dmem_n15798), .A2(MEM_stage_inst_dmem_n15797), .ZN(MEM_stage_inst_dmem_n11401) );
NAND2_X1 MEM_stage_inst_dmem_U13266 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n15826), .ZN(MEM_stage_inst_dmem_n15797) );
NAND2_X1 MEM_stage_inst_dmem_U13265 ( .A1(MEM_stage_inst_dmem_ram_1102), .A2(MEM_stage_inst_dmem_n15825), .ZN(MEM_stage_inst_dmem_n15798) );
NAND2_X1 MEM_stage_inst_dmem_U13264 ( .A1(MEM_stage_inst_dmem_n15796), .A2(MEM_stage_inst_dmem_n15795), .ZN(MEM_stage_inst_dmem_n11402) );
NAND2_X1 MEM_stage_inst_dmem_U13263 ( .A1(MEM_stage_inst_dmem_n16758), .A2(MEM_stage_inst_dmem_n15826), .ZN(MEM_stage_inst_dmem_n15795) );
INV_X1 MEM_stage_inst_dmem_U13262 ( .A(MEM_stage_inst_dmem_n15825), .ZN(MEM_stage_inst_dmem_n15826) );
NAND2_X1 MEM_stage_inst_dmem_U13261 ( .A1(MEM_stage_inst_dmem_ram_1103), .A2(MEM_stage_inst_dmem_n15825), .ZN(MEM_stage_inst_dmem_n15796) );
NAND2_X1 MEM_stage_inst_dmem_U13260 ( .A1(MEM_stage_inst_dmem_n21319), .A2(MEM_stage_inst_dmem_n15931), .ZN(MEM_stage_inst_dmem_n15825) );
NAND2_X1 MEM_stage_inst_dmem_U13259 ( .A1(MEM_stage_inst_dmem_n15794), .A2(MEM_stage_inst_dmem_n15793), .ZN(MEM_stage_inst_dmem_n11403) );
NAND2_X1 MEM_stage_inst_dmem_U13258 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n15792), .ZN(MEM_stage_inst_dmem_n15793) );
NAND2_X1 MEM_stage_inst_dmem_U13257 ( .A1(MEM_stage_inst_dmem_ram_1104), .A2(MEM_stage_inst_dmem_n15791), .ZN(MEM_stage_inst_dmem_n15794) );
NAND2_X1 MEM_stage_inst_dmem_U13256 ( .A1(MEM_stage_inst_dmem_n15790), .A2(MEM_stage_inst_dmem_n15789), .ZN(MEM_stage_inst_dmem_n11404) );
NAND2_X1 MEM_stage_inst_dmem_U13255 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n15792), .ZN(MEM_stage_inst_dmem_n15789) );
NAND2_X1 MEM_stage_inst_dmem_U13254 ( .A1(MEM_stage_inst_dmem_ram_1105), .A2(MEM_stage_inst_dmem_n15791), .ZN(MEM_stage_inst_dmem_n15790) );
NAND2_X1 MEM_stage_inst_dmem_U13253 ( .A1(MEM_stage_inst_dmem_n15788), .A2(MEM_stage_inst_dmem_n15787), .ZN(MEM_stage_inst_dmem_n11405) );
NAND2_X1 MEM_stage_inst_dmem_U13252 ( .A1(MEM_stage_inst_dmem_n20544), .A2(MEM_stage_inst_dmem_n15792), .ZN(MEM_stage_inst_dmem_n15787) );
NAND2_X1 MEM_stage_inst_dmem_U13251 ( .A1(MEM_stage_inst_dmem_ram_1106), .A2(MEM_stage_inst_dmem_n15791), .ZN(MEM_stage_inst_dmem_n15788) );
NAND2_X1 MEM_stage_inst_dmem_U13250 ( .A1(MEM_stage_inst_dmem_n15786), .A2(MEM_stage_inst_dmem_n15785), .ZN(MEM_stage_inst_dmem_n11406) );
NAND2_X1 MEM_stage_inst_dmem_U13249 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n15792), .ZN(MEM_stage_inst_dmem_n15785) );
NAND2_X1 MEM_stage_inst_dmem_U13248 ( .A1(MEM_stage_inst_dmem_ram_1107), .A2(MEM_stage_inst_dmem_n15791), .ZN(MEM_stage_inst_dmem_n15786) );
NAND2_X1 MEM_stage_inst_dmem_U13247 ( .A1(MEM_stage_inst_dmem_n15784), .A2(MEM_stage_inst_dmem_n15783), .ZN(MEM_stage_inst_dmem_n11407) );
NAND2_X1 MEM_stage_inst_dmem_U13246 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n15792), .ZN(MEM_stage_inst_dmem_n15783) );
NAND2_X1 MEM_stage_inst_dmem_U13245 ( .A1(MEM_stage_inst_dmem_ram_1108), .A2(MEM_stage_inst_dmem_n15791), .ZN(MEM_stage_inst_dmem_n15784) );
NAND2_X1 MEM_stage_inst_dmem_U13244 ( .A1(MEM_stage_inst_dmem_n15782), .A2(MEM_stage_inst_dmem_n15781), .ZN(MEM_stage_inst_dmem_n11408) );
NAND2_X1 MEM_stage_inst_dmem_U13243 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n15792), .ZN(MEM_stage_inst_dmem_n15781) );
NAND2_X1 MEM_stage_inst_dmem_U13242 ( .A1(MEM_stage_inst_dmem_ram_1109), .A2(MEM_stage_inst_dmem_n15791), .ZN(MEM_stage_inst_dmem_n15782) );
NAND2_X1 MEM_stage_inst_dmem_U13241 ( .A1(MEM_stage_inst_dmem_n15780), .A2(MEM_stage_inst_dmem_n15779), .ZN(MEM_stage_inst_dmem_n11409) );
NAND2_X1 MEM_stage_inst_dmem_U13240 ( .A1(EX_pipeline_reg_out_11), .A2(MEM_stage_inst_dmem_n15792), .ZN(MEM_stage_inst_dmem_n15779) );
NAND2_X1 MEM_stage_inst_dmem_U13239 ( .A1(MEM_stage_inst_dmem_ram_1110), .A2(MEM_stage_inst_dmem_n15791), .ZN(MEM_stage_inst_dmem_n15780) );
NAND2_X1 MEM_stage_inst_dmem_U13238 ( .A1(MEM_stage_inst_dmem_n15778), .A2(MEM_stage_inst_dmem_n15777), .ZN(MEM_stage_inst_dmem_n11410) );
NAND2_X1 MEM_stage_inst_dmem_U13237 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n15792), .ZN(MEM_stage_inst_dmem_n15777) );
NAND2_X1 MEM_stage_inst_dmem_U13236 ( .A1(MEM_stage_inst_dmem_ram_1111), .A2(MEM_stage_inst_dmem_n15791), .ZN(MEM_stage_inst_dmem_n15778) );
NAND2_X1 MEM_stage_inst_dmem_U13235 ( .A1(MEM_stage_inst_dmem_n15776), .A2(MEM_stage_inst_dmem_n15775), .ZN(MEM_stage_inst_dmem_n11411) );
NAND2_X1 MEM_stage_inst_dmem_U13234 ( .A1(MEM_stage_inst_dmem_n20527), .A2(MEM_stage_inst_dmem_n15792), .ZN(MEM_stage_inst_dmem_n15775) );
NAND2_X1 MEM_stage_inst_dmem_U13233 ( .A1(MEM_stage_inst_dmem_ram_1112), .A2(MEM_stage_inst_dmem_n15791), .ZN(MEM_stage_inst_dmem_n15776) );
NAND2_X1 MEM_stage_inst_dmem_U13232 ( .A1(MEM_stage_inst_dmem_n15774), .A2(MEM_stage_inst_dmem_n15773), .ZN(MEM_stage_inst_dmem_n11412) );
NAND2_X1 MEM_stage_inst_dmem_U13231 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n15792), .ZN(MEM_stage_inst_dmem_n15773) );
NAND2_X1 MEM_stage_inst_dmem_U13230 ( .A1(MEM_stage_inst_dmem_ram_1113), .A2(MEM_stage_inst_dmem_n15791), .ZN(MEM_stage_inst_dmem_n15774) );
NAND2_X1 MEM_stage_inst_dmem_U13229 ( .A1(MEM_stage_inst_dmem_n15772), .A2(MEM_stage_inst_dmem_n15771), .ZN(MEM_stage_inst_dmem_n11413) );
NAND2_X1 MEM_stage_inst_dmem_U13228 ( .A1(MEM_stage_inst_dmem_n20521), .A2(MEM_stage_inst_dmem_n15792), .ZN(MEM_stage_inst_dmem_n15771) );
NAND2_X1 MEM_stage_inst_dmem_U13227 ( .A1(MEM_stage_inst_dmem_ram_1114), .A2(MEM_stage_inst_dmem_n15791), .ZN(MEM_stage_inst_dmem_n15772) );
NAND2_X1 MEM_stage_inst_dmem_U13226 ( .A1(MEM_stage_inst_dmem_n15770), .A2(MEM_stage_inst_dmem_n15769), .ZN(MEM_stage_inst_dmem_n11414) );
NAND2_X1 MEM_stage_inst_dmem_U13225 ( .A1(MEM_stage_inst_dmem_n20518), .A2(MEM_stage_inst_dmem_n15792), .ZN(MEM_stage_inst_dmem_n15769) );
NAND2_X1 MEM_stage_inst_dmem_U13224 ( .A1(MEM_stage_inst_dmem_ram_1115), .A2(MEM_stage_inst_dmem_n15791), .ZN(MEM_stage_inst_dmem_n15770) );
NAND2_X1 MEM_stage_inst_dmem_U13223 ( .A1(MEM_stage_inst_dmem_n15768), .A2(MEM_stage_inst_dmem_n15767), .ZN(MEM_stage_inst_dmem_n11415) );
NAND2_X1 MEM_stage_inst_dmem_U13222 ( .A1(MEM_stage_inst_dmem_n20515), .A2(MEM_stage_inst_dmem_n15792), .ZN(MEM_stage_inst_dmem_n15767) );
NAND2_X1 MEM_stage_inst_dmem_U13221 ( .A1(MEM_stage_inst_dmem_ram_1116), .A2(MEM_stage_inst_dmem_n15791), .ZN(MEM_stage_inst_dmem_n15768) );
NAND2_X1 MEM_stage_inst_dmem_U13220 ( .A1(MEM_stage_inst_dmem_n15766), .A2(MEM_stage_inst_dmem_n15765), .ZN(MEM_stage_inst_dmem_n11416) );
NAND2_X1 MEM_stage_inst_dmem_U13219 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n15792), .ZN(MEM_stage_inst_dmem_n15765) );
NAND2_X1 MEM_stage_inst_dmem_U13218 ( .A1(MEM_stage_inst_dmem_ram_1117), .A2(MEM_stage_inst_dmem_n15791), .ZN(MEM_stage_inst_dmem_n15766) );
NAND2_X1 MEM_stage_inst_dmem_U13217 ( .A1(MEM_stage_inst_dmem_n15764), .A2(MEM_stage_inst_dmem_n15763), .ZN(MEM_stage_inst_dmem_n11417) );
NAND2_X1 MEM_stage_inst_dmem_U13216 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n15792), .ZN(MEM_stage_inst_dmem_n15763) );
NAND2_X1 MEM_stage_inst_dmem_U13215 ( .A1(MEM_stage_inst_dmem_ram_1118), .A2(MEM_stage_inst_dmem_n15791), .ZN(MEM_stage_inst_dmem_n15764) );
NAND2_X1 MEM_stage_inst_dmem_U13214 ( .A1(MEM_stage_inst_dmem_n15762), .A2(MEM_stage_inst_dmem_n15761), .ZN(MEM_stage_inst_dmem_n11418) );
NAND2_X1 MEM_stage_inst_dmem_U13213 ( .A1(MEM_stage_inst_dmem_n15110), .A2(MEM_stage_inst_dmem_n15792), .ZN(MEM_stage_inst_dmem_n15761) );
INV_X1 MEM_stage_inst_dmem_U13212 ( .A(MEM_stage_inst_dmem_n15791), .ZN(MEM_stage_inst_dmem_n15792) );
NAND2_X1 MEM_stage_inst_dmem_U13211 ( .A1(MEM_stage_inst_dmem_ram_1119), .A2(MEM_stage_inst_dmem_n15791), .ZN(MEM_stage_inst_dmem_n15762) );
NAND2_X1 MEM_stage_inst_dmem_U13210 ( .A1(MEM_stage_inst_dmem_n21284), .A2(MEM_stage_inst_dmem_n15931), .ZN(MEM_stage_inst_dmem_n15791) );
NAND2_X1 MEM_stage_inst_dmem_U13209 ( .A1(MEM_stage_inst_dmem_n15760), .A2(MEM_stage_inst_dmem_n15759), .ZN(MEM_stage_inst_dmem_n11419) );
NAND2_X1 MEM_stage_inst_dmem_U13208 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n15758), .ZN(MEM_stage_inst_dmem_n15759) );
NAND2_X1 MEM_stage_inst_dmem_U13207 ( .A1(MEM_stage_inst_dmem_ram_1120), .A2(MEM_stage_inst_dmem_n15757), .ZN(MEM_stage_inst_dmem_n15760) );
NAND2_X1 MEM_stage_inst_dmem_U13206 ( .A1(MEM_stage_inst_dmem_n15756), .A2(MEM_stage_inst_dmem_n15755), .ZN(MEM_stage_inst_dmem_n11420) );
NAND2_X1 MEM_stage_inst_dmem_U13205 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n15758), .ZN(MEM_stage_inst_dmem_n15755) );
NAND2_X1 MEM_stage_inst_dmem_U13204 ( .A1(MEM_stage_inst_dmem_ram_1121), .A2(MEM_stage_inst_dmem_n15757), .ZN(MEM_stage_inst_dmem_n15756) );
NAND2_X1 MEM_stage_inst_dmem_U13203 ( .A1(MEM_stage_inst_dmem_n15754), .A2(MEM_stage_inst_dmem_n15753), .ZN(MEM_stage_inst_dmem_n11421) );
NAND2_X1 MEM_stage_inst_dmem_U13202 ( .A1(MEM_stage_inst_dmem_n16789), .A2(MEM_stage_inst_dmem_n15758), .ZN(MEM_stage_inst_dmem_n15753) );
NAND2_X1 MEM_stage_inst_dmem_U13201 ( .A1(MEM_stage_inst_dmem_ram_1122), .A2(MEM_stage_inst_dmem_n15757), .ZN(MEM_stage_inst_dmem_n15754) );
NAND2_X1 MEM_stage_inst_dmem_U13200 ( .A1(MEM_stage_inst_dmem_n15752), .A2(MEM_stage_inst_dmem_n15751), .ZN(MEM_stage_inst_dmem_n11422) );
NAND2_X1 MEM_stage_inst_dmem_U13199 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n15758), .ZN(MEM_stage_inst_dmem_n15751) );
NAND2_X1 MEM_stage_inst_dmem_U13198 ( .A1(MEM_stage_inst_dmem_ram_1123), .A2(MEM_stage_inst_dmem_n15757), .ZN(MEM_stage_inst_dmem_n15752) );
NAND2_X1 MEM_stage_inst_dmem_U13197 ( .A1(MEM_stage_inst_dmem_n15750), .A2(MEM_stage_inst_dmem_n15749), .ZN(MEM_stage_inst_dmem_n11423) );
NAND2_X1 MEM_stage_inst_dmem_U13196 ( .A1(MEM_stage_inst_dmem_n16784), .A2(MEM_stage_inst_dmem_n15758), .ZN(MEM_stage_inst_dmem_n15749) );
NAND2_X1 MEM_stage_inst_dmem_U13195 ( .A1(MEM_stage_inst_dmem_ram_1124), .A2(MEM_stage_inst_dmem_n15757), .ZN(MEM_stage_inst_dmem_n15750) );
NAND2_X1 MEM_stage_inst_dmem_U13194 ( .A1(MEM_stage_inst_dmem_n15748), .A2(MEM_stage_inst_dmem_n15747), .ZN(MEM_stage_inst_dmem_n11424) );
NAND2_X1 MEM_stage_inst_dmem_U13193 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n15758), .ZN(MEM_stage_inst_dmem_n15747) );
NAND2_X1 MEM_stage_inst_dmem_U13192 ( .A1(MEM_stage_inst_dmem_ram_1125), .A2(MEM_stage_inst_dmem_n15757), .ZN(MEM_stage_inst_dmem_n15748) );
NAND2_X1 MEM_stage_inst_dmem_U13191 ( .A1(MEM_stage_inst_dmem_n15746), .A2(MEM_stage_inst_dmem_n15745), .ZN(MEM_stage_inst_dmem_n11425) );
NAND2_X1 MEM_stage_inst_dmem_U13190 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n15758), .ZN(MEM_stage_inst_dmem_n15745) );
NAND2_X1 MEM_stage_inst_dmem_U13189 ( .A1(MEM_stage_inst_dmem_ram_1126), .A2(MEM_stage_inst_dmem_n15757), .ZN(MEM_stage_inst_dmem_n15746) );
NAND2_X1 MEM_stage_inst_dmem_U13188 ( .A1(MEM_stage_inst_dmem_n15744), .A2(MEM_stage_inst_dmem_n15743), .ZN(MEM_stage_inst_dmem_n11426) );
NAND2_X1 MEM_stage_inst_dmem_U13187 ( .A1(MEM_stage_inst_dmem_n16777), .A2(MEM_stage_inst_dmem_n15758), .ZN(MEM_stage_inst_dmem_n15743) );
NAND2_X1 MEM_stage_inst_dmem_U13186 ( .A1(MEM_stage_inst_dmem_ram_1127), .A2(MEM_stage_inst_dmem_n15757), .ZN(MEM_stage_inst_dmem_n15744) );
NAND2_X1 MEM_stage_inst_dmem_U13185 ( .A1(MEM_stage_inst_dmem_n15742), .A2(MEM_stage_inst_dmem_n15741), .ZN(MEM_stage_inst_dmem_n11427) );
NAND2_X1 MEM_stage_inst_dmem_U13184 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n15758), .ZN(MEM_stage_inst_dmem_n15741) );
NAND2_X1 MEM_stage_inst_dmem_U13183 ( .A1(MEM_stage_inst_dmem_ram_1128), .A2(MEM_stage_inst_dmem_n15757), .ZN(MEM_stage_inst_dmem_n15742) );
NAND2_X1 MEM_stage_inst_dmem_U13182 ( .A1(MEM_stage_inst_dmem_n15740), .A2(MEM_stage_inst_dmem_n15739), .ZN(MEM_stage_inst_dmem_n11428) );
NAND2_X1 MEM_stage_inst_dmem_U13181 ( .A1(MEM_stage_inst_dmem_n16772), .A2(MEM_stage_inst_dmem_n15758), .ZN(MEM_stage_inst_dmem_n15739) );
NAND2_X1 MEM_stage_inst_dmem_U13180 ( .A1(MEM_stage_inst_dmem_ram_1129), .A2(MEM_stage_inst_dmem_n15757), .ZN(MEM_stage_inst_dmem_n15740) );
NAND2_X1 MEM_stage_inst_dmem_U13179 ( .A1(MEM_stage_inst_dmem_n15738), .A2(MEM_stage_inst_dmem_n15737), .ZN(MEM_stage_inst_dmem_n11429) );
NAND2_X1 MEM_stage_inst_dmem_U13178 ( .A1(MEM_stage_inst_dmem_n16769), .A2(MEM_stage_inst_dmem_n15758), .ZN(MEM_stage_inst_dmem_n15737) );
NAND2_X1 MEM_stage_inst_dmem_U13177 ( .A1(MEM_stage_inst_dmem_ram_1130), .A2(MEM_stage_inst_dmem_n15757), .ZN(MEM_stage_inst_dmem_n15738) );
NAND2_X1 MEM_stage_inst_dmem_U13176 ( .A1(MEM_stage_inst_dmem_n15736), .A2(MEM_stage_inst_dmem_n15735), .ZN(MEM_stage_inst_dmem_n11430) );
NAND2_X1 MEM_stage_inst_dmem_U13175 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n15758), .ZN(MEM_stage_inst_dmem_n15735) );
NAND2_X1 MEM_stage_inst_dmem_U13174 ( .A1(MEM_stage_inst_dmem_ram_1131), .A2(MEM_stage_inst_dmem_n15757), .ZN(MEM_stage_inst_dmem_n15736) );
NAND2_X1 MEM_stage_inst_dmem_U13173 ( .A1(MEM_stage_inst_dmem_n15734), .A2(MEM_stage_inst_dmem_n15733), .ZN(MEM_stage_inst_dmem_n11431) );
NAND2_X1 MEM_stage_inst_dmem_U13172 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n15758), .ZN(MEM_stage_inst_dmem_n15733) );
NAND2_X1 MEM_stage_inst_dmem_U13171 ( .A1(MEM_stage_inst_dmem_ram_1132), .A2(MEM_stage_inst_dmem_n15757), .ZN(MEM_stage_inst_dmem_n15734) );
NAND2_X1 MEM_stage_inst_dmem_U13170 ( .A1(MEM_stage_inst_dmem_n15732), .A2(MEM_stage_inst_dmem_n15731), .ZN(MEM_stage_inst_dmem_n11432) );
NAND2_X1 MEM_stage_inst_dmem_U13169 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n15758), .ZN(MEM_stage_inst_dmem_n15731) );
NAND2_X1 MEM_stage_inst_dmem_U13168 ( .A1(MEM_stage_inst_dmem_ram_1133), .A2(MEM_stage_inst_dmem_n15757), .ZN(MEM_stage_inst_dmem_n15732) );
NAND2_X1 MEM_stage_inst_dmem_U13167 ( .A1(MEM_stage_inst_dmem_n15730), .A2(MEM_stage_inst_dmem_n15729), .ZN(MEM_stage_inst_dmem_n11433) );
NAND2_X1 MEM_stage_inst_dmem_U13166 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n15758), .ZN(MEM_stage_inst_dmem_n15729) );
NAND2_X1 MEM_stage_inst_dmem_U13165 ( .A1(MEM_stage_inst_dmem_ram_1134), .A2(MEM_stage_inst_dmem_n15757), .ZN(MEM_stage_inst_dmem_n15730) );
NAND2_X1 MEM_stage_inst_dmem_U13164 ( .A1(MEM_stage_inst_dmem_n15728), .A2(MEM_stage_inst_dmem_n15727), .ZN(MEM_stage_inst_dmem_n11434) );
NAND2_X1 MEM_stage_inst_dmem_U13163 ( .A1(MEM_stage_inst_dmem_n16758), .A2(MEM_stage_inst_dmem_n15758), .ZN(MEM_stage_inst_dmem_n15727) );
INV_X1 MEM_stage_inst_dmem_U13162 ( .A(MEM_stage_inst_dmem_n15757), .ZN(MEM_stage_inst_dmem_n15758) );
NAND2_X1 MEM_stage_inst_dmem_U13161 ( .A1(MEM_stage_inst_dmem_ram_1135), .A2(MEM_stage_inst_dmem_n15757), .ZN(MEM_stage_inst_dmem_n15728) );
NAND2_X1 MEM_stage_inst_dmem_U13160 ( .A1(MEM_stage_inst_dmem_n21249), .A2(MEM_stage_inst_dmem_n15931), .ZN(MEM_stage_inst_dmem_n15757) );
NAND2_X1 MEM_stage_inst_dmem_U13159 ( .A1(MEM_stage_inst_dmem_n15726), .A2(MEM_stage_inst_dmem_n15725), .ZN(MEM_stage_inst_dmem_n11435) );
NAND2_X1 MEM_stage_inst_dmem_U13158 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n15724), .ZN(MEM_stage_inst_dmem_n15725) );
NAND2_X1 MEM_stage_inst_dmem_U13157 ( .A1(MEM_stage_inst_dmem_ram_1136), .A2(MEM_stage_inst_dmem_n15723), .ZN(MEM_stage_inst_dmem_n15726) );
NAND2_X1 MEM_stage_inst_dmem_U13156 ( .A1(MEM_stage_inst_dmem_n15722), .A2(MEM_stage_inst_dmem_n15721), .ZN(MEM_stage_inst_dmem_n11436) );
NAND2_X1 MEM_stage_inst_dmem_U13155 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n15724), .ZN(MEM_stage_inst_dmem_n15721) );
NAND2_X1 MEM_stage_inst_dmem_U13154 ( .A1(MEM_stage_inst_dmem_ram_1137), .A2(MEM_stage_inst_dmem_n15723), .ZN(MEM_stage_inst_dmem_n15722) );
NAND2_X1 MEM_stage_inst_dmem_U13153 ( .A1(MEM_stage_inst_dmem_n15720), .A2(MEM_stage_inst_dmem_n15719), .ZN(MEM_stage_inst_dmem_n11437) );
NAND2_X1 MEM_stage_inst_dmem_U13152 ( .A1(EX_pipeline_reg_out_7), .A2(MEM_stage_inst_dmem_n15724), .ZN(MEM_stage_inst_dmem_n15719) );
NAND2_X1 MEM_stage_inst_dmem_U13151 ( .A1(MEM_stage_inst_dmem_ram_1138), .A2(MEM_stage_inst_dmem_n15723), .ZN(MEM_stage_inst_dmem_n15720) );
NAND2_X1 MEM_stage_inst_dmem_U13150 ( .A1(MEM_stage_inst_dmem_n15718), .A2(MEM_stage_inst_dmem_n15717), .ZN(MEM_stage_inst_dmem_n11438) );
NAND2_X1 MEM_stage_inst_dmem_U13149 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n15724), .ZN(MEM_stage_inst_dmem_n15717) );
NAND2_X1 MEM_stage_inst_dmem_U13148 ( .A1(MEM_stage_inst_dmem_ram_1139), .A2(MEM_stage_inst_dmem_n15723), .ZN(MEM_stage_inst_dmem_n15718) );
NAND2_X1 MEM_stage_inst_dmem_U13147 ( .A1(MEM_stage_inst_dmem_n15716), .A2(MEM_stage_inst_dmem_n15715), .ZN(MEM_stage_inst_dmem_n11439) );
NAND2_X1 MEM_stage_inst_dmem_U13146 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n15724), .ZN(MEM_stage_inst_dmem_n15715) );
NAND2_X1 MEM_stage_inst_dmem_U13145 ( .A1(MEM_stage_inst_dmem_ram_1140), .A2(MEM_stage_inst_dmem_n15723), .ZN(MEM_stage_inst_dmem_n15716) );
NAND2_X1 MEM_stage_inst_dmem_U13144 ( .A1(MEM_stage_inst_dmem_n15714), .A2(MEM_stage_inst_dmem_n15713), .ZN(MEM_stage_inst_dmem_n11440) );
NAND2_X1 MEM_stage_inst_dmem_U13143 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n15724), .ZN(MEM_stage_inst_dmem_n15713) );
NAND2_X1 MEM_stage_inst_dmem_U13142 ( .A1(MEM_stage_inst_dmem_ram_1141), .A2(MEM_stage_inst_dmem_n15723), .ZN(MEM_stage_inst_dmem_n15714) );
NAND2_X1 MEM_stage_inst_dmem_U13141 ( .A1(MEM_stage_inst_dmem_n15712), .A2(MEM_stage_inst_dmem_n15711), .ZN(MEM_stage_inst_dmem_n11441) );
NAND2_X1 MEM_stage_inst_dmem_U13140 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n15724), .ZN(MEM_stage_inst_dmem_n15711) );
NAND2_X1 MEM_stage_inst_dmem_U13139 ( .A1(MEM_stage_inst_dmem_ram_1142), .A2(MEM_stage_inst_dmem_n15723), .ZN(MEM_stage_inst_dmem_n15712) );
NAND2_X1 MEM_stage_inst_dmem_U13138 ( .A1(MEM_stage_inst_dmem_n15710), .A2(MEM_stage_inst_dmem_n15709), .ZN(MEM_stage_inst_dmem_n11442) );
NAND2_X1 MEM_stage_inst_dmem_U13137 ( .A1(MEM_stage_inst_dmem_n13886), .A2(MEM_stage_inst_dmem_n15724), .ZN(MEM_stage_inst_dmem_n15709) );
NAND2_X1 MEM_stage_inst_dmem_U13136 ( .A1(MEM_stage_inst_dmem_ram_1143), .A2(MEM_stage_inst_dmem_n15723), .ZN(MEM_stage_inst_dmem_n15710) );
NAND2_X1 MEM_stage_inst_dmem_U13135 ( .A1(MEM_stage_inst_dmem_n15708), .A2(MEM_stage_inst_dmem_n15707), .ZN(MEM_stage_inst_dmem_n11443) );
NAND2_X1 MEM_stage_inst_dmem_U13134 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n15724), .ZN(MEM_stage_inst_dmem_n15707) );
NAND2_X1 MEM_stage_inst_dmem_U13133 ( .A1(MEM_stage_inst_dmem_ram_1144), .A2(MEM_stage_inst_dmem_n15723), .ZN(MEM_stage_inst_dmem_n15708) );
NAND2_X1 MEM_stage_inst_dmem_U13132 ( .A1(MEM_stage_inst_dmem_n15706), .A2(MEM_stage_inst_dmem_n15705), .ZN(MEM_stage_inst_dmem_n11444) );
NAND2_X1 MEM_stage_inst_dmem_U13131 ( .A1(MEM_stage_inst_dmem_n19251), .A2(MEM_stage_inst_dmem_n15724), .ZN(MEM_stage_inst_dmem_n15705) );
NAND2_X1 MEM_stage_inst_dmem_U13130 ( .A1(MEM_stage_inst_dmem_ram_1145), .A2(MEM_stage_inst_dmem_n15723), .ZN(MEM_stage_inst_dmem_n15706) );
NAND2_X1 MEM_stage_inst_dmem_U13129 ( .A1(MEM_stage_inst_dmem_n15704), .A2(MEM_stage_inst_dmem_n15703), .ZN(MEM_stage_inst_dmem_n11445) );
NAND2_X1 MEM_stage_inst_dmem_U13128 ( .A1(EX_pipeline_reg_out_15), .A2(MEM_stage_inst_dmem_n15724), .ZN(MEM_stage_inst_dmem_n15703) );
NAND2_X1 MEM_stage_inst_dmem_U13127 ( .A1(MEM_stage_inst_dmem_ram_1146), .A2(MEM_stage_inst_dmem_n15723), .ZN(MEM_stage_inst_dmem_n15704) );
NAND2_X1 MEM_stage_inst_dmem_U13126 ( .A1(MEM_stage_inst_dmem_n15702), .A2(MEM_stage_inst_dmem_n15701), .ZN(MEM_stage_inst_dmem_n11446) );
NAND2_X1 MEM_stage_inst_dmem_U13125 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n15724), .ZN(MEM_stage_inst_dmem_n15701) );
NAND2_X1 MEM_stage_inst_dmem_U13124 ( .A1(MEM_stage_inst_dmem_ram_1147), .A2(MEM_stage_inst_dmem_n15723), .ZN(MEM_stage_inst_dmem_n15702) );
NAND2_X1 MEM_stage_inst_dmem_U13123 ( .A1(MEM_stage_inst_dmem_n15700), .A2(MEM_stage_inst_dmem_n15699), .ZN(MEM_stage_inst_dmem_n11447) );
NAND2_X1 MEM_stage_inst_dmem_U13122 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n15724), .ZN(MEM_stage_inst_dmem_n15699) );
NAND2_X1 MEM_stage_inst_dmem_U13121 ( .A1(MEM_stage_inst_dmem_ram_1148), .A2(MEM_stage_inst_dmem_n15723), .ZN(MEM_stage_inst_dmem_n15700) );
NAND2_X1 MEM_stage_inst_dmem_U13120 ( .A1(MEM_stage_inst_dmem_n15698), .A2(MEM_stage_inst_dmem_n15697), .ZN(MEM_stage_inst_dmem_n11448) );
NAND2_X1 MEM_stage_inst_dmem_U13119 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n15724), .ZN(MEM_stage_inst_dmem_n15697) );
NAND2_X1 MEM_stage_inst_dmem_U13118 ( .A1(MEM_stage_inst_dmem_ram_1149), .A2(MEM_stage_inst_dmem_n15723), .ZN(MEM_stage_inst_dmem_n15698) );
NAND2_X1 MEM_stage_inst_dmem_U13117 ( .A1(MEM_stage_inst_dmem_n15696), .A2(MEM_stage_inst_dmem_n15695), .ZN(MEM_stage_inst_dmem_n11449) );
NAND2_X1 MEM_stage_inst_dmem_U13116 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n15724), .ZN(MEM_stage_inst_dmem_n15695) );
NAND2_X1 MEM_stage_inst_dmem_U13115 ( .A1(MEM_stage_inst_dmem_ram_1150), .A2(MEM_stage_inst_dmem_n15723), .ZN(MEM_stage_inst_dmem_n15696) );
NAND2_X1 MEM_stage_inst_dmem_U13114 ( .A1(MEM_stage_inst_dmem_n15694), .A2(MEM_stage_inst_dmem_n15693), .ZN(MEM_stage_inst_dmem_n11450) );
NAND2_X1 MEM_stage_inst_dmem_U13113 ( .A1(MEM_stage_inst_dmem_n14693), .A2(MEM_stage_inst_dmem_n15724), .ZN(MEM_stage_inst_dmem_n15693) );
INV_X1 MEM_stage_inst_dmem_U13112 ( .A(MEM_stage_inst_dmem_n15723), .ZN(MEM_stage_inst_dmem_n15724) );
NAND2_X1 MEM_stage_inst_dmem_U13111 ( .A1(MEM_stage_inst_dmem_ram_1151), .A2(MEM_stage_inst_dmem_n15723), .ZN(MEM_stage_inst_dmem_n15694) );
NAND2_X1 MEM_stage_inst_dmem_U13110 ( .A1(MEM_stage_inst_dmem_n21214), .A2(MEM_stage_inst_dmem_n15931), .ZN(MEM_stage_inst_dmem_n15723) );
NAND2_X1 MEM_stage_inst_dmem_U13109 ( .A1(MEM_stage_inst_dmem_n15692), .A2(MEM_stage_inst_dmem_n15691), .ZN(MEM_stage_inst_dmem_n11451) );
NAND2_X1 MEM_stage_inst_dmem_U13108 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n15690), .ZN(MEM_stage_inst_dmem_n15691) );
NAND2_X1 MEM_stage_inst_dmem_U13107 ( .A1(MEM_stage_inst_dmem_ram_1152), .A2(MEM_stage_inst_dmem_n15689), .ZN(MEM_stage_inst_dmem_n15692) );
NAND2_X1 MEM_stage_inst_dmem_U13106 ( .A1(MEM_stage_inst_dmem_n15688), .A2(MEM_stage_inst_dmem_n15687), .ZN(MEM_stage_inst_dmem_n11452) );
NAND2_X1 MEM_stage_inst_dmem_U13105 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n15690), .ZN(MEM_stage_inst_dmem_n15687) );
NAND2_X1 MEM_stage_inst_dmem_U13104 ( .A1(MEM_stage_inst_dmem_ram_1153), .A2(MEM_stage_inst_dmem_n15689), .ZN(MEM_stage_inst_dmem_n15688) );
NAND2_X1 MEM_stage_inst_dmem_U13103 ( .A1(MEM_stage_inst_dmem_n15686), .A2(MEM_stage_inst_dmem_n15685), .ZN(MEM_stage_inst_dmem_n11453) );
NAND2_X1 MEM_stage_inst_dmem_U13102 ( .A1(MEM_stage_inst_dmem_n16789), .A2(MEM_stage_inst_dmem_n15690), .ZN(MEM_stage_inst_dmem_n15685) );
NAND2_X1 MEM_stage_inst_dmem_U13101 ( .A1(MEM_stage_inst_dmem_ram_1154), .A2(MEM_stage_inst_dmem_n15689), .ZN(MEM_stage_inst_dmem_n15686) );
NAND2_X1 MEM_stage_inst_dmem_U13100 ( .A1(MEM_stage_inst_dmem_n15684), .A2(MEM_stage_inst_dmem_n15683), .ZN(MEM_stage_inst_dmem_n11454) );
NAND2_X1 MEM_stage_inst_dmem_U13099 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n15690), .ZN(MEM_stage_inst_dmem_n15683) );
NAND2_X1 MEM_stage_inst_dmem_U13098 ( .A1(MEM_stage_inst_dmem_ram_1155), .A2(MEM_stage_inst_dmem_n15689), .ZN(MEM_stage_inst_dmem_n15684) );
NAND2_X1 MEM_stage_inst_dmem_U13097 ( .A1(MEM_stage_inst_dmem_n15682), .A2(MEM_stage_inst_dmem_n15681), .ZN(MEM_stage_inst_dmem_n11455) );
NAND2_X1 MEM_stage_inst_dmem_U13096 ( .A1(MEM_stage_inst_dmem_n16784), .A2(MEM_stage_inst_dmem_n15690), .ZN(MEM_stage_inst_dmem_n15681) );
NAND2_X1 MEM_stage_inst_dmem_U13095 ( .A1(MEM_stage_inst_dmem_ram_1156), .A2(MEM_stage_inst_dmem_n15689), .ZN(MEM_stage_inst_dmem_n15682) );
NAND2_X1 MEM_stage_inst_dmem_U13094 ( .A1(MEM_stage_inst_dmem_n15680), .A2(MEM_stage_inst_dmem_n15679), .ZN(MEM_stage_inst_dmem_n11456) );
NAND2_X1 MEM_stage_inst_dmem_U13093 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n15690), .ZN(MEM_stage_inst_dmem_n15679) );
NAND2_X1 MEM_stage_inst_dmem_U13092 ( .A1(MEM_stage_inst_dmem_ram_1157), .A2(MEM_stage_inst_dmem_n15689), .ZN(MEM_stage_inst_dmem_n15680) );
NAND2_X1 MEM_stage_inst_dmem_U13091 ( .A1(MEM_stage_inst_dmem_n15678), .A2(MEM_stage_inst_dmem_n15677), .ZN(MEM_stage_inst_dmem_n11457) );
NAND2_X1 MEM_stage_inst_dmem_U13090 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n15690), .ZN(MEM_stage_inst_dmem_n15677) );
NAND2_X1 MEM_stage_inst_dmem_U13089 ( .A1(MEM_stage_inst_dmem_ram_1158), .A2(MEM_stage_inst_dmem_n15689), .ZN(MEM_stage_inst_dmem_n15678) );
NAND2_X1 MEM_stage_inst_dmem_U13088 ( .A1(MEM_stage_inst_dmem_n15676), .A2(MEM_stage_inst_dmem_n15675), .ZN(MEM_stage_inst_dmem_n11458) );
NAND2_X1 MEM_stage_inst_dmem_U13087 ( .A1(MEM_stage_inst_dmem_n16777), .A2(MEM_stage_inst_dmem_n15690), .ZN(MEM_stage_inst_dmem_n15675) );
NAND2_X1 MEM_stage_inst_dmem_U13086 ( .A1(MEM_stage_inst_dmem_ram_1159), .A2(MEM_stage_inst_dmem_n15689), .ZN(MEM_stage_inst_dmem_n15676) );
NAND2_X1 MEM_stage_inst_dmem_U13085 ( .A1(MEM_stage_inst_dmem_n15674), .A2(MEM_stage_inst_dmem_n15673), .ZN(MEM_stage_inst_dmem_n11459) );
NAND2_X1 MEM_stage_inst_dmem_U13084 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n15690), .ZN(MEM_stage_inst_dmem_n15673) );
NAND2_X1 MEM_stage_inst_dmem_U13083 ( .A1(MEM_stage_inst_dmem_ram_1160), .A2(MEM_stage_inst_dmem_n15689), .ZN(MEM_stage_inst_dmem_n15674) );
NAND2_X1 MEM_stage_inst_dmem_U13082 ( .A1(MEM_stage_inst_dmem_n15672), .A2(MEM_stage_inst_dmem_n15671), .ZN(MEM_stage_inst_dmem_n11460) );
NAND2_X1 MEM_stage_inst_dmem_U13081 ( .A1(MEM_stage_inst_dmem_n16772), .A2(MEM_stage_inst_dmem_n15690), .ZN(MEM_stage_inst_dmem_n15671) );
NAND2_X1 MEM_stage_inst_dmem_U13080 ( .A1(MEM_stage_inst_dmem_ram_1161), .A2(MEM_stage_inst_dmem_n15689), .ZN(MEM_stage_inst_dmem_n15672) );
NAND2_X1 MEM_stage_inst_dmem_U13079 ( .A1(MEM_stage_inst_dmem_n15670), .A2(MEM_stage_inst_dmem_n15669), .ZN(MEM_stage_inst_dmem_n11461) );
NAND2_X1 MEM_stage_inst_dmem_U13078 ( .A1(MEM_stage_inst_dmem_n16769), .A2(MEM_stage_inst_dmem_n15690), .ZN(MEM_stage_inst_dmem_n15669) );
NAND2_X1 MEM_stage_inst_dmem_U13077 ( .A1(MEM_stage_inst_dmem_ram_1162), .A2(MEM_stage_inst_dmem_n15689), .ZN(MEM_stage_inst_dmem_n15670) );
NAND2_X1 MEM_stage_inst_dmem_U13076 ( .A1(MEM_stage_inst_dmem_n15668), .A2(MEM_stage_inst_dmem_n15667), .ZN(MEM_stage_inst_dmem_n11462) );
NAND2_X1 MEM_stage_inst_dmem_U13075 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n15690), .ZN(MEM_stage_inst_dmem_n15667) );
NAND2_X1 MEM_stage_inst_dmem_U13074 ( .A1(MEM_stage_inst_dmem_ram_1163), .A2(MEM_stage_inst_dmem_n15689), .ZN(MEM_stage_inst_dmem_n15668) );
NAND2_X1 MEM_stage_inst_dmem_U13073 ( .A1(MEM_stage_inst_dmem_n15666), .A2(MEM_stage_inst_dmem_n15665), .ZN(MEM_stage_inst_dmem_n11463) );
NAND2_X1 MEM_stage_inst_dmem_U13072 ( .A1(MEM_stage_inst_dmem_n21474), .A2(MEM_stage_inst_dmem_n15690), .ZN(MEM_stage_inst_dmem_n15665) );
NAND2_X1 MEM_stage_inst_dmem_U13071 ( .A1(MEM_stage_inst_dmem_ram_1164), .A2(MEM_stage_inst_dmem_n15689), .ZN(MEM_stage_inst_dmem_n15666) );
NAND2_X1 MEM_stage_inst_dmem_U13070 ( .A1(MEM_stage_inst_dmem_n15664), .A2(MEM_stage_inst_dmem_n15663), .ZN(MEM_stage_inst_dmem_n11464) );
NAND2_X1 MEM_stage_inst_dmem_U13069 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n15690), .ZN(MEM_stage_inst_dmem_n15663) );
NAND2_X1 MEM_stage_inst_dmem_U13068 ( .A1(MEM_stage_inst_dmem_ram_1165), .A2(MEM_stage_inst_dmem_n15689), .ZN(MEM_stage_inst_dmem_n15664) );
NAND2_X1 MEM_stage_inst_dmem_U13067 ( .A1(MEM_stage_inst_dmem_n15662), .A2(MEM_stage_inst_dmem_n15661), .ZN(MEM_stage_inst_dmem_n11465) );
NAND2_X1 MEM_stage_inst_dmem_U13066 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n15690), .ZN(MEM_stage_inst_dmem_n15661) );
NAND2_X1 MEM_stage_inst_dmem_U13065 ( .A1(MEM_stage_inst_dmem_ram_1166), .A2(MEM_stage_inst_dmem_n15689), .ZN(MEM_stage_inst_dmem_n15662) );
NAND2_X1 MEM_stage_inst_dmem_U13064 ( .A1(MEM_stage_inst_dmem_n15660), .A2(MEM_stage_inst_dmem_n15659), .ZN(MEM_stage_inst_dmem_n11466) );
NAND2_X1 MEM_stage_inst_dmem_U13063 ( .A1(MEM_stage_inst_dmem_n16758), .A2(MEM_stage_inst_dmem_n15690), .ZN(MEM_stage_inst_dmem_n15659) );
INV_X1 MEM_stage_inst_dmem_U13062 ( .A(MEM_stage_inst_dmem_n15689), .ZN(MEM_stage_inst_dmem_n15690) );
NAND2_X1 MEM_stage_inst_dmem_U13061 ( .A1(MEM_stage_inst_dmem_ram_1167), .A2(MEM_stage_inst_dmem_n15689), .ZN(MEM_stage_inst_dmem_n15660) );
NAND2_X1 MEM_stage_inst_dmem_U13060 ( .A1(MEM_stage_inst_dmem_n21179), .A2(MEM_stage_inst_dmem_n15931), .ZN(MEM_stage_inst_dmem_n15689) );
NAND2_X1 MEM_stage_inst_dmem_U13059 ( .A1(MEM_stage_inst_dmem_n15658), .A2(MEM_stage_inst_dmem_n15657), .ZN(MEM_stage_inst_dmem_n11467) );
NAND2_X1 MEM_stage_inst_dmem_U13058 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n15656), .ZN(MEM_stage_inst_dmem_n15657) );
NAND2_X1 MEM_stage_inst_dmem_U13057 ( .A1(MEM_stage_inst_dmem_ram_1168), .A2(MEM_stage_inst_dmem_n15655), .ZN(MEM_stage_inst_dmem_n15658) );
NAND2_X1 MEM_stage_inst_dmem_U13056 ( .A1(MEM_stage_inst_dmem_n15654), .A2(MEM_stage_inst_dmem_n15653), .ZN(MEM_stage_inst_dmem_n11468) );
NAND2_X1 MEM_stage_inst_dmem_U13055 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n15656), .ZN(MEM_stage_inst_dmem_n15653) );
NAND2_X1 MEM_stage_inst_dmem_U13054 ( .A1(MEM_stage_inst_dmem_ram_1169), .A2(MEM_stage_inst_dmem_n15655), .ZN(MEM_stage_inst_dmem_n15654) );
NAND2_X1 MEM_stage_inst_dmem_U13053 ( .A1(MEM_stage_inst_dmem_n15652), .A2(MEM_stage_inst_dmem_n15651), .ZN(MEM_stage_inst_dmem_n11469) );
NAND2_X1 MEM_stage_inst_dmem_U13052 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n15656), .ZN(MEM_stage_inst_dmem_n15651) );
NAND2_X1 MEM_stage_inst_dmem_U13051 ( .A1(MEM_stage_inst_dmem_ram_1170), .A2(MEM_stage_inst_dmem_n15655), .ZN(MEM_stage_inst_dmem_n15652) );
NAND2_X1 MEM_stage_inst_dmem_U13050 ( .A1(MEM_stage_inst_dmem_n15650), .A2(MEM_stage_inst_dmem_n15649), .ZN(MEM_stage_inst_dmem_n11470) );
NAND2_X1 MEM_stage_inst_dmem_U13049 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n15656), .ZN(MEM_stage_inst_dmem_n15649) );
NAND2_X1 MEM_stage_inst_dmem_U13048 ( .A1(MEM_stage_inst_dmem_ram_1171), .A2(MEM_stage_inst_dmem_n15655), .ZN(MEM_stage_inst_dmem_n15650) );
NAND2_X1 MEM_stage_inst_dmem_U13047 ( .A1(MEM_stage_inst_dmem_n15648), .A2(MEM_stage_inst_dmem_n15647), .ZN(MEM_stage_inst_dmem_n11471) );
NAND2_X1 MEM_stage_inst_dmem_U13046 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n15656), .ZN(MEM_stage_inst_dmem_n15647) );
NAND2_X1 MEM_stage_inst_dmem_U13045 ( .A1(MEM_stage_inst_dmem_ram_1172), .A2(MEM_stage_inst_dmem_n15655), .ZN(MEM_stage_inst_dmem_n15648) );
NAND2_X1 MEM_stage_inst_dmem_U13044 ( .A1(MEM_stage_inst_dmem_n15646), .A2(MEM_stage_inst_dmem_n15645), .ZN(MEM_stage_inst_dmem_n11472) );
NAND2_X1 MEM_stage_inst_dmem_U13043 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n15656), .ZN(MEM_stage_inst_dmem_n15645) );
NAND2_X1 MEM_stage_inst_dmem_U13042 ( .A1(MEM_stage_inst_dmem_ram_1173), .A2(MEM_stage_inst_dmem_n15655), .ZN(MEM_stage_inst_dmem_n15646) );
NAND2_X1 MEM_stage_inst_dmem_U13041 ( .A1(MEM_stage_inst_dmem_n15644), .A2(MEM_stage_inst_dmem_n15643), .ZN(MEM_stage_inst_dmem_n11473) );
NAND2_X1 MEM_stage_inst_dmem_U13040 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n15656), .ZN(MEM_stage_inst_dmem_n15643) );
NAND2_X1 MEM_stage_inst_dmem_U13039 ( .A1(MEM_stage_inst_dmem_ram_1174), .A2(MEM_stage_inst_dmem_n15655), .ZN(MEM_stage_inst_dmem_n15644) );
NAND2_X1 MEM_stage_inst_dmem_U13038 ( .A1(MEM_stage_inst_dmem_n15642), .A2(MEM_stage_inst_dmem_n15641), .ZN(MEM_stage_inst_dmem_n11474) );
NAND2_X1 MEM_stage_inst_dmem_U13037 ( .A1(EX_pipeline_reg_out_12), .A2(MEM_stage_inst_dmem_n15656), .ZN(MEM_stage_inst_dmem_n15641) );
NAND2_X1 MEM_stage_inst_dmem_U13036 ( .A1(MEM_stage_inst_dmem_ram_1175), .A2(MEM_stage_inst_dmem_n15655), .ZN(MEM_stage_inst_dmem_n15642) );
NAND2_X1 MEM_stage_inst_dmem_U13035 ( .A1(MEM_stage_inst_dmem_n15640), .A2(MEM_stage_inst_dmem_n15639), .ZN(MEM_stage_inst_dmem_n11475) );
NAND2_X1 MEM_stage_inst_dmem_U13034 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n15656), .ZN(MEM_stage_inst_dmem_n15639) );
NAND2_X1 MEM_stage_inst_dmem_U13033 ( .A1(MEM_stage_inst_dmem_ram_1176), .A2(MEM_stage_inst_dmem_n15655), .ZN(MEM_stage_inst_dmem_n15640) );
NAND2_X1 MEM_stage_inst_dmem_U13032 ( .A1(MEM_stage_inst_dmem_n15638), .A2(MEM_stage_inst_dmem_n15637), .ZN(MEM_stage_inst_dmem_n11476) );
NAND2_X1 MEM_stage_inst_dmem_U13031 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n15656), .ZN(MEM_stage_inst_dmem_n15637) );
NAND2_X1 MEM_stage_inst_dmem_U13030 ( .A1(MEM_stage_inst_dmem_ram_1177), .A2(MEM_stage_inst_dmem_n15655), .ZN(MEM_stage_inst_dmem_n15638) );
NAND2_X1 MEM_stage_inst_dmem_U13029 ( .A1(MEM_stage_inst_dmem_n15636), .A2(MEM_stage_inst_dmem_n15635), .ZN(MEM_stage_inst_dmem_n11477) );
NAND2_X1 MEM_stage_inst_dmem_U13028 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n15656), .ZN(MEM_stage_inst_dmem_n15635) );
NAND2_X1 MEM_stage_inst_dmem_U13027 ( .A1(MEM_stage_inst_dmem_ram_1178), .A2(MEM_stage_inst_dmem_n15655), .ZN(MEM_stage_inst_dmem_n15636) );
NAND2_X1 MEM_stage_inst_dmem_U13026 ( .A1(MEM_stage_inst_dmem_n15634), .A2(MEM_stage_inst_dmem_n15633), .ZN(MEM_stage_inst_dmem_n11478) );
NAND2_X1 MEM_stage_inst_dmem_U13025 ( .A1(MEM_stage_inst_dmem_n20518), .A2(MEM_stage_inst_dmem_n15656), .ZN(MEM_stage_inst_dmem_n15633) );
NAND2_X1 MEM_stage_inst_dmem_U13024 ( .A1(MEM_stage_inst_dmem_ram_1179), .A2(MEM_stage_inst_dmem_n15655), .ZN(MEM_stage_inst_dmem_n15634) );
NAND2_X1 MEM_stage_inst_dmem_U13023 ( .A1(MEM_stage_inst_dmem_n15632), .A2(MEM_stage_inst_dmem_n15631), .ZN(MEM_stage_inst_dmem_n11479) );
NAND2_X1 MEM_stage_inst_dmem_U13022 ( .A1(MEM_stage_inst_dmem_n20515), .A2(MEM_stage_inst_dmem_n15656), .ZN(MEM_stage_inst_dmem_n15631) );
NAND2_X1 MEM_stage_inst_dmem_U13021 ( .A1(MEM_stage_inst_dmem_ram_1180), .A2(MEM_stage_inst_dmem_n15655), .ZN(MEM_stage_inst_dmem_n15632) );
NAND2_X1 MEM_stage_inst_dmem_U13020 ( .A1(MEM_stage_inst_dmem_n15630), .A2(MEM_stage_inst_dmem_n15629), .ZN(MEM_stage_inst_dmem_n11480) );
NAND2_X1 MEM_stage_inst_dmem_U13019 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n15656), .ZN(MEM_stage_inst_dmem_n15629) );
NAND2_X1 MEM_stage_inst_dmem_U13018 ( .A1(MEM_stage_inst_dmem_ram_1181), .A2(MEM_stage_inst_dmem_n15655), .ZN(MEM_stage_inst_dmem_n15630) );
NAND2_X1 MEM_stage_inst_dmem_U13017 ( .A1(MEM_stage_inst_dmem_n15628), .A2(MEM_stage_inst_dmem_n15627), .ZN(MEM_stage_inst_dmem_n11481) );
NAND2_X1 MEM_stage_inst_dmem_U13016 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n15656), .ZN(MEM_stage_inst_dmem_n15627) );
NAND2_X1 MEM_stage_inst_dmem_U13015 ( .A1(MEM_stage_inst_dmem_ram_1182), .A2(MEM_stage_inst_dmem_n15655), .ZN(MEM_stage_inst_dmem_n15628) );
NAND2_X1 MEM_stage_inst_dmem_U13014 ( .A1(MEM_stage_inst_dmem_n15626), .A2(MEM_stage_inst_dmem_n15625), .ZN(MEM_stage_inst_dmem_n11482) );
NAND2_X1 MEM_stage_inst_dmem_U13013 ( .A1(MEM_stage_inst_dmem_n16343), .A2(MEM_stage_inst_dmem_n15656), .ZN(MEM_stage_inst_dmem_n15625) );
INV_X1 MEM_stage_inst_dmem_U13012 ( .A(MEM_stage_inst_dmem_n15655), .ZN(MEM_stage_inst_dmem_n15656) );
NAND2_X1 MEM_stage_inst_dmem_U13011 ( .A1(MEM_stage_inst_dmem_ram_1183), .A2(MEM_stage_inst_dmem_n15655), .ZN(MEM_stage_inst_dmem_n15626) );
NAND2_X1 MEM_stage_inst_dmem_U13010 ( .A1(MEM_stage_inst_dmem_n21144), .A2(MEM_stage_inst_dmem_n15931), .ZN(MEM_stage_inst_dmem_n15655) );
NAND2_X1 MEM_stage_inst_dmem_U13009 ( .A1(MEM_stage_inst_dmem_n15624), .A2(MEM_stage_inst_dmem_n15623), .ZN(MEM_stage_inst_dmem_n11483) );
NAND2_X1 MEM_stage_inst_dmem_U13008 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n15622), .ZN(MEM_stage_inst_dmem_n15623) );
NAND2_X1 MEM_stage_inst_dmem_U13007 ( .A1(MEM_stage_inst_dmem_ram_1184), .A2(MEM_stage_inst_dmem_n15621), .ZN(MEM_stage_inst_dmem_n15624) );
NAND2_X1 MEM_stage_inst_dmem_U13006 ( .A1(MEM_stage_inst_dmem_n15620), .A2(MEM_stage_inst_dmem_n15619), .ZN(MEM_stage_inst_dmem_n11484) );
NAND2_X1 MEM_stage_inst_dmem_U13005 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n15622), .ZN(MEM_stage_inst_dmem_n15619) );
NAND2_X1 MEM_stage_inst_dmem_U13004 ( .A1(MEM_stage_inst_dmem_ram_1185), .A2(MEM_stage_inst_dmem_n15621), .ZN(MEM_stage_inst_dmem_n15620) );
NAND2_X1 MEM_stage_inst_dmem_U13003 ( .A1(MEM_stage_inst_dmem_n15618), .A2(MEM_stage_inst_dmem_n15617), .ZN(MEM_stage_inst_dmem_n11485) );
NAND2_X1 MEM_stage_inst_dmem_U13002 ( .A1(MEM_stage_inst_dmem_n16789), .A2(MEM_stage_inst_dmem_n15622), .ZN(MEM_stage_inst_dmem_n15617) );
BUF_X1 MEM_stage_inst_dmem_U13001 ( .A(MEM_stage_inst_dmem_n113), .Z(MEM_stage_inst_dmem_n16789) );
NAND2_X1 MEM_stage_inst_dmem_U13000 ( .A1(MEM_stage_inst_dmem_ram_1186), .A2(MEM_stage_inst_dmem_n15621), .ZN(MEM_stage_inst_dmem_n15618) );
NAND2_X1 MEM_stage_inst_dmem_U12999 ( .A1(MEM_stage_inst_dmem_n15616), .A2(MEM_stage_inst_dmem_n15615), .ZN(MEM_stage_inst_dmem_n11486) );
NAND2_X1 MEM_stage_inst_dmem_U12998 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n15622), .ZN(MEM_stage_inst_dmem_n15615) );
NAND2_X1 MEM_stage_inst_dmem_U12997 ( .A1(MEM_stage_inst_dmem_ram_1187), .A2(MEM_stage_inst_dmem_n15621), .ZN(MEM_stage_inst_dmem_n15616) );
NAND2_X1 MEM_stage_inst_dmem_U12996 ( .A1(MEM_stage_inst_dmem_n15614), .A2(MEM_stage_inst_dmem_n15613), .ZN(MEM_stage_inst_dmem_n11487) );
NAND2_X1 MEM_stage_inst_dmem_U12995 ( .A1(MEM_stage_inst_dmem_n16784), .A2(MEM_stage_inst_dmem_n15622), .ZN(MEM_stage_inst_dmem_n15613) );
NAND2_X1 MEM_stage_inst_dmem_U12994 ( .A1(MEM_stage_inst_dmem_ram_1188), .A2(MEM_stage_inst_dmem_n15621), .ZN(MEM_stage_inst_dmem_n15614) );
NAND2_X1 MEM_stage_inst_dmem_U12993 ( .A1(MEM_stage_inst_dmem_n15612), .A2(MEM_stage_inst_dmem_n15611), .ZN(MEM_stage_inst_dmem_n11488) );
NAND2_X1 MEM_stage_inst_dmem_U12992 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n15622), .ZN(MEM_stage_inst_dmem_n15611) );
NAND2_X1 MEM_stage_inst_dmem_U12991 ( .A1(MEM_stage_inst_dmem_ram_1189), .A2(MEM_stage_inst_dmem_n15621), .ZN(MEM_stage_inst_dmem_n15612) );
NAND2_X1 MEM_stage_inst_dmem_U12990 ( .A1(MEM_stage_inst_dmem_n15610), .A2(MEM_stage_inst_dmem_n15609), .ZN(MEM_stage_inst_dmem_n11489) );
NAND2_X1 MEM_stage_inst_dmem_U12989 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n15622), .ZN(MEM_stage_inst_dmem_n15609) );
NAND2_X1 MEM_stage_inst_dmem_U12988 ( .A1(MEM_stage_inst_dmem_ram_1190), .A2(MEM_stage_inst_dmem_n15621), .ZN(MEM_stage_inst_dmem_n15610) );
NAND2_X1 MEM_stage_inst_dmem_U12987 ( .A1(MEM_stage_inst_dmem_n15608), .A2(MEM_stage_inst_dmem_n15607), .ZN(MEM_stage_inst_dmem_n11490) );
NAND2_X1 MEM_stage_inst_dmem_U12986 ( .A1(MEM_stage_inst_dmem_n16777), .A2(MEM_stage_inst_dmem_n15622), .ZN(MEM_stage_inst_dmem_n15607) );
BUF_X1 MEM_stage_inst_dmem_U12985 ( .A(MEM_stage_inst_dmem_n17), .Z(MEM_stage_inst_dmem_n16777) );
NAND2_X1 MEM_stage_inst_dmem_U12984 ( .A1(MEM_stage_inst_dmem_ram_1191), .A2(MEM_stage_inst_dmem_n15621), .ZN(MEM_stage_inst_dmem_n15608) );
NAND2_X1 MEM_stage_inst_dmem_U12983 ( .A1(MEM_stage_inst_dmem_n15606), .A2(MEM_stage_inst_dmem_n15605), .ZN(MEM_stage_inst_dmem_n11491) );
NAND2_X1 MEM_stage_inst_dmem_U12982 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n15622), .ZN(MEM_stage_inst_dmem_n15605) );
NAND2_X1 MEM_stage_inst_dmem_U12981 ( .A1(MEM_stage_inst_dmem_ram_1192), .A2(MEM_stage_inst_dmem_n15621), .ZN(MEM_stage_inst_dmem_n15606) );
NAND2_X1 MEM_stage_inst_dmem_U12980 ( .A1(MEM_stage_inst_dmem_n15604), .A2(MEM_stage_inst_dmem_n15603), .ZN(MEM_stage_inst_dmem_n11492) );
NAND2_X1 MEM_stage_inst_dmem_U12979 ( .A1(MEM_stage_inst_dmem_n16772), .A2(MEM_stage_inst_dmem_n15622), .ZN(MEM_stage_inst_dmem_n15603) );
BUF_X1 MEM_stage_inst_dmem_U12978 ( .A(MEM_stage_inst_dmem_n100), .Z(MEM_stage_inst_dmem_n16772) );
NAND2_X1 MEM_stage_inst_dmem_U12977 ( .A1(MEM_stage_inst_dmem_ram_1193), .A2(MEM_stage_inst_dmem_n15621), .ZN(MEM_stage_inst_dmem_n15604) );
NAND2_X1 MEM_stage_inst_dmem_U12976 ( .A1(MEM_stage_inst_dmem_n15602), .A2(MEM_stage_inst_dmem_n15601), .ZN(MEM_stage_inst_dmem_n11493) );
NAND2_X1 MEM_stage_inst_dmem_U12975 ( .A1(MEM_stage_inst_dmem_n16769), .A2(MEM_stage_inst_dmem_n15622), .ZN(MEM_stage_inst_dmem_n15601) );
BUF_X1 MEM_stage_inst_dmem_U12974 ( .A(MEM_stage_inst_dmem_n102), .Z(MEM_stage_inst_dmem_n16769) );
NAND2_X1 MEM_stage_inst_dmem_U12973 ( .A1(MEM_stage_inst_dmem_ram_1194), .A2(MEM_stage_inst_dmem_n15621), .ZN(MEM_stage_inst_dmem_n15602) );
NAND2_X1 MEM_stage_inst_dmem_U12972 ( .A1(MEM_stage_inst_dmem_n15600), .A2(MEM_stage_inst_dmem_n15599), .ZN(MEM_stage_inst_dmem_n11494) );
NAND2_X1 MEM_stage_inst_dmem_U12971 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n15622), .ZN(MEM_stage_inst_dmem_n15599) );
NAND2_X1 MEM_stage_inst_dmem_U12970 ( .A1(MEM_stage_inst_dmem_ram_1195), .A2(MEM_stage_inst_dmem_n15621), .ZN(MEM_stage_inst_dmem_n15600) );
NAND2_X1 MEM_stage_inst_dmem_U12969 ( .A1(MEM_stage_inst_dmem_n15598), .A2(MEM_stage_inst_dmem_n15597), .ZN(MEM_stage_inst_dmem_n11495) );
NAND2_X1 MEM_stage_inst_dmem_U12968 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n15622), .ZN(MEM_stage_inst_dmem_n15597) );
NAND2_X1 MEM_stage_inst_dmem_U12967 ( .A1(MEM_stage_inst_dmem_ram_1196), .A2(MEM_stage_inst_dmem_n15621), .ZN(MEM_stage_inst_dmem_n15598) );
NAND2_X1 MEM_stage_inst_dmem_U12966 ( .A1(MEM_stage_inst_dmem_n15596), .A2(MEM_stage_inst_dmem_n15595), .ZN(MEM_stage_inst_dmem_n11496) );
NAND2_X1 MEM_stage_inst_dmem_U12965 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n15622), .ZN(MEM_stage_inst_dmem_n15595) );
NAND2_X1 MEM_stage_inst_dmem_U12964 ( .A1(MEM_stage_inst_dmem_ram_1197), .A2(MEM_stage_inst_dmem_n15621), .ZN(MEM_stage_inst_dmem_n15596) );
NAND2_X1 MEM_stage_inst_dmem_U12963 ( .A1(MEM_stage_inst_dmem_n15594), .A2(MEM_stage_inst_dmem_n15593), .ZN(MEM_stage_inst_dmem_n11497) );
NAND2_X1 MEM_stage_inst_dmem_U12962 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n15622), .ZN(MEM_stage_inst_dmem_n15593) );
NAND2_X1 MEM_stage_inst_dmem_U12961 ( .A1(MEM_stage_inst_dmem_ram_1198), .A2(MEM_stage_inst_dmem_n15621), .ZN(MEM_stage_inst_dmem_n15594) );
NAND2_X1 MEM_stage_inst_dmem_U12960 ( .A1(MEM_stage_inst_dmem_n15592), .A2(MEM_stage_inst_dmem_n15591), .ZN(MEM_stage_inst_dmem_n11498) );
NAND2_X1 MEM_stage_inst_dmem_U12959 ( .A1(MEM_stage_inst_dmem_n16758), .A2(MEM_stage_inst_dmem_n15622), .ZN(MEM_stage_inst_dmem_n15591) );
INV_X1 MEM_stage_inst_dmem_U12958 ( .A(MEM_stage_inst_dmem_n15621), .ZN(MEM_stage_inst_dmem_n15622) );
NAND2_X1 MEM_stage_inst_dmem_U12957 ( .A1(MEM_stage_inst_dmem_ram_1199), .A2(MEM_stage_inst_dmem_n15621), .ZN(MEM_stage_inst_dmem_n15592) );
NAND2_X1 MEM_stage_inst_dmem_U12956 ( .A1(MEM_stage_inst_dmem_n21109), .A2(MEM_stage_inst_dmem_n15931), .ZN(MEM_stage_inst_dmem_n15621) );
NAND2_X1 MEM_stage_inst_dmem_U12955 ( .A1(MEM_stage_inst_dmem_n15590), .A2(MEM_stage_inst_dmem_n15589), .ZN(MEM_stage_inst_dmem_n11499) );
NAND2_X1 MEM_stage_inst_dmem_U12954 ( .A1(MEM_stage_inst_dmem_n20551), .A2(MEM_stage_inst_dmem_n15588), .ZN(MEM_stage_inst_dmem_n15589) );
NAND2_X1 MEM_stage_inst_dmem_U12953 ( .A1(MEM_stage_inst_dmem_ram_1200), .A2(MEM_stage_inst_dmem_n15587), .ZN(MEM_stage_inst_dmem_n15590) );
NAND2_X1 MEM_stage_inst_dmem_U12952 ( .A1(MEM_stage_inst_dmem_n15586), .A2(MEM_stage_inst_dmem_n15585), .ZN(MEM_stage_inst_dmem_n11500) );
NAND2_X1 MEM_stage_inst_dmem_U12951 ( .A1(MEM_stage_inst_dmem_n20547), .A2(MEM_stage_inst_dmem_n15588), .ZN(MEM_stage_inst_dmem_n15585) );
NAND2_X1 MEM_stage_inst_dmem_U12950 ( .A1(MEM_stage_inst_dmem_ram_1201), .A2(MEM_stage_inst_dmem_n15587), .ZN(MEM_stage_inst_dmem_n15586) );
NAND2_X1 MEM_stage_inst_dmem_U12949 ( .A1(MEM_stage_inst_dmem_n15584), .A2(MEM_stage_inst_dmem_n15583), .ZN(MEM_stage_inst_dmem_n11501) );
NAND2_X1 MEM_stage_inst_dmem_U12948 ( .A1(MEM_stage_inst_dmem_n20544), .A2(MEM_stage_inst_dmem_n15588), .ZN(MEM_stage_inst_dmem_n15583) );
NAND2_X1 MEM_stage_inst_dmem_U12947 ( .A1(MEM_stage_inst_dmem_ram_1202), .A2(MEM_stage_inst_dmem_n15587), .ZN(MEM_stage_inst_dmem_n15584) );
NAND2_X1 MEM_stage_inst_dmem_U12946 ( .A1(MEM_stage_inst_dmem_n15582), .A2(MEM_stage_inst_dmem_n15581), .ZN(MEM_stage_inst_dmem_n11502) );
NAND2_X1 MEM_stage_inst_dmem_U12945 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n15588), .ZN(MEM_stage_inst_dmem_n15581) );
NAND2_X1 MEM_stage_inst_dmem_U12944 ( .A1(MEM_stage_inst_dmem_ram_1203), .A2(MEM_stage_inst_dmem_n15587), .ZN(MEM_stage_inst_dmem_n15582) );
NAND2_X1 MEM_stage_inst_dmem_U12943 ( .A1(MEM_stage_inst_dmem_n15580), .A2(MEM_stage_inst_dmem_n15579), .ZN(MEM_stage_inst_dmem_n11503) );
NAND2_X1 MEM_stage_inst_dmem_U12942 ( .A1(MEM_stage_inst_dmem_n16368), .A2(MEM_stage_inst_dmem_n15588), .ZN(MEM_stage_inst_dmem_n15579) );
NAND2_X1 MEM_stage_inst_dmem_U12941 ( .A1(MEM_stage_inst_dmem_ram_1204), .A2(MEM_stage_inst_dmem_n15587), .ZN(MEM_stage_inst_dmem_n15580) );
NAND2_X1 MEM_stage_inst_dmem_U12940 ( .A1(MEM_stage_inst_dmem_n15578), .A2(MEM_stage_inst_dmem_n15577), .ZN(MEM_stage_inst_dmem_n11504) );
NAND2_X1 MEM_stage_inst_dmem_U12939 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n15588), .ZN(MEM_stage_inst_dmem_n15577) );
NAND2_X1 MEM_stage_inst_dmem_U12938 ( .A1(MEM_stage_inst_dmem_ram_1205), .A2(MEM_stage_inst_dmem_n15587), .ZN(MEM_stage_inst_dmem_n15578) );
NAND2_X1 MEM_stage_inst_dmem_U12937 ( .A1(MEM_stage_inst_dmem_n15576), .A2(MEM_stage_inst_dmem_n15575), .ZN(MEM_stage_inst_dmem_n11505) );
NAND2_X1 MEM_stage_inst_dmem_U12936 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n15588), .ZN(MEM_stage_inst_dmem_n15575) );
NAND2_X1 MEM_stage_inst_dmem_U12935 ( .A1(MEM_stage_inst_dmem_ram_1206), .A2(MEM_stage_inst_dmem_n15587), .ZN(MEM_stage_inst_dmem_n15576) );
NAND2_X1 MEM_stage_inst_dmem_U12934 ( .A1(MEM_stage_inst_dmem_n15574), .A2(MEM_stage_inst_dmem_n15573), .ZN(MEM_stage_inst_dmem_n11506) );
NAND2_X1 MEM_stage_inst_dmem_U12933 ( .A1(MEM_stage_inst_dmem_n20530), .A2(MEM_stage_inst_dmem_n15588), .ZN(MEM_stage_inst_dmem_n15573) );
NAND2_X1 MEM_stage_inst_dmem_U12932 ( .A1(MEM_stage_inst_dmem_ram_1207), .A2(MEM_stage_inst_dmem_n15587), .ZN(MEM_stage_inst_dmem_n15574) );
NAND2_X1 MEM_stage_inst_dmem_U12931 ( .A1(MEM_stage_inst_dmem_n15572), .A2(MEM_stage_inst_dmem_n15571), .ZN(MEM_stage_inst_dmem_n11507) );
NAND2_X1 MEM_stage_inst_dmem_U12930 ( .A1(MEM_stage_inst_dmem_n20527), .A2(MEM_stage_inst_dmem_n15588), .ZN(MEM_stage_inst_dmem_n15571) );
NAND2_X1 MEM_stage_inst_dmem_U12929 ( .A1(MEM_stage_inst_dmem_ram_1208), .A2(MEM_stage_inst_dmem_n15587), .ZN(MEM_stage_inst_dmem_n15572) );
NAND2_X1 MEM_stage_inst_dmem_U12928 ( .A1(MEM_stage_inst_dmem_n15570), .A2(MEM_stage_inst_dmem_n15569), .ZN(MEM_stage_inst_dmem_n11508) );
NAND2_X1 MEM_stage_inst_dmem_U12927 ( .A1(MEM_stage_inst_dmem_n20524), .A2(MEM_stage_inst_dmem_n15588), .ZN(MEM_stage_inst_dmem_n15569) );
NAND2_X1 MEM_stage_inst_dmem_U12926 ( .A1(MEM_stage_inst_dmem_ram_1209), .A2(MEM_stage_inst_dmem_n15587), .ZN(MEM_stage_inst_dmem_n15570) );
NAND2_X1 MEM_stage_inst_dmem_U12925 ( .A1(MEM_stage_inst_dmem_n15568), .A2(MEM_stage_inst_dmem_n15567), .ZN(MEM_stage_inst_dmem_n11509) );
NAND2_X1 MEM_stage_inst_dmem_U12924 ( .A1(MEM_stage_inst_dmem_n20521), .A2(MEM_stage_inst_dmem_n15588), .ZN(MEM_stage_inst_dmem_n15567) );
NAND2_X1 MEM_stage_inst_dmem_U12923 ( .A1(MEM_stage_inst_dmem_ram_1210), .A2(MEM_stage_inst_dmem_n15587), .ZN(MEM_stage_inst_dmem_n15568) );
NAND2_X1 MEM_stage_inst_dmem_U12922 ( .A1(MEM_stage_inst_dmem_n15566), .A2(MEM_stage_inst_dmem_n15565), .ZN(MEM_stage_inst_dmem_n11510) );
NAND2_X1 MEM_stage_inst_dmem_U12921 ( .A1(MEM_stage_inst_dmem_n20518), .A2(MEM_stage_inst_dmem_n15588), .ZN(MEM_stage_inst_dmem_n15565) );
NAND2_X1 MEM_stage_inst_dmem_U12920 ( .A1(MEM_stage_inst_dmem_ram_1211), .A2(MEM_stage_inst_dmem_n15587), .ZN(MEM_stage_inst_dmem_n15566) );
NAND2_X1 MEM_stage_inst_dmem_U12919 ( .A1(MEM_stage_inst_dmem_n15564), .A2(MEM_stage_inst_dmem_n15563), .ZN(MEM_stage_inst_dmem_n11511) );
NAND2_X1 MEM_stage_inst_dmem_U12918 ( .A1(MEM_stage_inst_dmem_n20515), .A2(MEM_stage_inst_dmem_n15588), .ZN(MEM_stage_inst_dmem_n15563) );
NAND2_X1 MEM_stage_inst_dmem_U12917 ( .A1(MEM_stage_inst_dmem_ram_1212), .A2(MEM_stage_inst_dmem_n15587), .ZN(MEM_stage_inst_dmem_n15564) );
NAND2_X1 MEM_stage_inst_dmem_U12916 ( .A1(MEM_stage_inst_dmem_n15562), .A2(MEM_stage_inst_dmem_n15561), .ZN(MEM_stage_inst_dmem_n11512) );
NAND2_X1 MEM_stage_inst_dmem_U12915 ( .A1(MEM_stage_inst_dmem_n20512), .A2(MEM_stage_inst_dmem_n15588), .ZN(MEM_stage_inst_dmem_n15561) );
NAND2_X1 MEM_stage_inst_dmem_U12914 ( .A1(MEM_stage_inst_dmem_ram_1213), .A2(MEM_stage_inst_dmem_n15587), .ZN(MEM_stage_inst_dmem_n15562) );
NAND2_X1 MEM_stage_inst_dmem_U12913 ( .A1(MEM_stage_inst_dmem_n15560), .A2(MEM_stage_inst_dmem_n15559), .ZN(MEM_stage_inst_dmem_n11513) );
NAND2_X1 MEM_stage_inst_dmem_U12912 ( .A1(MEM_stage_inst_dmem_n20509), .A2(MEM_stage_inst_dmem_n15588), .ZN(MEM_stage_inst_dmem_n15559) );
NAND2_X1 MEM_stage_inst_dmem_U12911 ( .A1(MEM_stage_inst_dmem_ram_1214), .A2(MEM_stage_inst_dmem_n15587), .ZN(MEM_stage_inst_dmem_n15560) );
NAND2_X1 MEM_stage_inst_dmem_U12910 ( .A1(MEM_stage_inst_dmem_n15558), .A2(MEM_stage_inst_dmem_n15557), .ZN(MEM_stage_inst_dmem_n11514) );
NAND2_X1 MEM_stage_inst_dmem_U12909 ( .A1(MEM_stage_inst_dmem_n20506), .A2(MEM_stage_inst_dmem_n15588), .ZN(MEM_stage_inst_dmem_n15557) );
NAND2_X1 MEM_stage_inst_dmem_U12908 ( .A1(MEM_stage_inst_dmem_ram_1215), .A2(MEM_stage_inst_dmem_n15587), .ZN(MEM_stage_inst_dmem_n15558) );
NAND2_X1 MEM_stage_inst_dmem_U12907 ( .A1(MEM_stage_inst_dmem_n21074), .A2(MEM_stage_inst_dmem_n15931), .ZN(MEM_stage_inst_dmem_n15587) );
NAND2_X1 MEM_stage_inst_dmem_U12906 ( .A1(MEM_stage_inst_dmem_n15556), .A2(MEM_stage_inst_dmem_n15555), .ZN(MEM_stage_inst_dmem_n11515) );
NAND2_X1 MEM_stage_inst_dmem_U12905 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n15554), .ZN(MEM_stage_inst_dmem_n15555) );
NAND2_X1 MEM_stage_inst_dmem_U12904 ( .A1(MEM_stage_inst_dmem_ram_1216), .A2(MEM_stage_inst_dmem_n15553), .ZN(MEM_stage_inst_dmem_n15556) );
NAND2_X1 MEM_stage_inst_dmem_U12903 ( .A1(MEM_stage_inst_dmem_n15552), .A2(MEM_stage_inst_dmem_n15551), .ZN(MEM_stage_inst_dmem_n11516) );
NAND2_X1 MEM_stage_inst_dmem_U12902 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n15554), .ZN(MEM_stage_inst_dmem_n15551) );
NAND2_X1 MEM_stage_inst_dmem_U12901 ( .A1(MEM_stage_inst_dmem_ram_1217), .A2(MEM_stage_inst_dmem_n15553), .ZN(MEM_stage_inst_dmem_n15552) );
NAND2_X1 MEM_stage_inst_dmem_U12900 ( .A1(MEM_stage_inst_dmem_n15550), .A2(MEM_stage_inst_dmem_n15549), .ZN(MEM_stage_inst_dmem_n11517) );
NAND2_X1 MEM_stage_inst_dmem_U12899 ( .A1(MEM_stage_inst_dmem_n18887), .A2(MEM_stage_inst_dmem_n15554), .ZN(MEM_stage_inst_dmem_n15549) );
NAND2_X1 MEM_stage_inst_dmem_U12898 ( .A1(MEM_stage_inst_dmem_ram_1218), .A2(MEM_stage_inst_dmem_n15553), .ZN(MEM_stage_inst_dmem_n15550) );
NAND2_X1 MEM_stage_inst_dmem_U12897 ( .A1(MEM_stage_inst_dmem_n15548), .A2(MEM_stage_inst_dmem_n15547), .ZN(MEM_stage_inst_dmem_n11518) );
NAND2_X1 MEM_stage_inst_dmem_U12896 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n15554), .ZN(MEM_stage_inst_dmem_n15547) );
NAND2_X1 MEM_stage_inst_dmem_U12895 ( .A1(MEM_stage_inst_dmem_ram_1219), .A2(MEM_stage_inst_dmem_n15553), .ZN(MEM_stage_inst_dmem_n15548) );
NAND2_X1 MEM_stage_inst_dmem_U12894 ( .A1(MEM_stage_inst_dmem_n15546), .A2(MEM_stage_inst_dmem_n15545), .ZN(MEM_stage_inst_dmem_n11519) );
NAND2_X1 MEM_stage_inst_dmem_U12893 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n15554), .ZN(MEM_stage_inst_dmem_n15545) );
NAND2_X1 MEM_stage_inst_dmem_U12892 ( .A1(MEM_stage_inst_dmem_ram_1220), .A2(MEM_stage_inst_dmem_n15553), .ZN(MEM_stage_inst_dmem_n15546) );
NAND2_X1 MEM_stage_inst_dmem_U12891 ( .A1(MEM_stage_inst_dmem_n15544), .A2(MEM_stage_inst_dmem_n15543), .ZN(MEM_stage_inst_dmem_n11520) );
NAND2_X1 MEM_stage_inst_dmem_U12890 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n15554), .ZN(MEM_stage_inst_dmem_n15543) );
NAND2_X1 MEM_stage_inst_dmem_U12889 ( .A1(MEM_stage_inst_dmem_ram_1221), .A2(MEM_stage_inst_dmem_n15553), .ZN(MEM_stage_inst_dmem_n15544) );
NAND2_X1 MEM_stage_inst_dmem_U12888 ( .A1(MEM_stage_inst_dmem_n15542), .A2(MEM_stage_inst_dmem_n15541), .ZN(MEM_stage_inst_dmem_n11521) );
NAND2_X1 MEM_stage_inst_dmem_U12887 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n15554), .ZN(MEM_stage_inst_dmem_n15541) );
NAND2_X1 MEM_stage_inst_dmem_U12886 ( .A1(MEM_stage_inst_dmem_ram_1222), .A2(MEM_stage_inst_dmem_n15553), .ZN(MEM_stage_inst_dmem_n15542) );
NAND2_X1 MEM_stage_inst_dmem_U12885 ( .A1(MEM_stage_inst_dmem_n15540), .A2(MEM_stage_inst_dmem_n15539), .ZN(MEM_stage_inst_dmem_n11522) );
NAND2_X1 MEM_stage_inst_dmem_U12884 ( .A1(MEM_stage_inst_dmem_n18875), .A2(MEM_stage_inst_dmem_n15554), .ZN(MEM_stage_inst_dmem_n15539) );
NAND2_X1 MEM_stage_inst_dmem_U12883 ( .A1(MEM_stage_inst_dmem_ram_1223), .A2(MEM_stage_inst_dmem_n15553), .ZN(MEM_stage_inst_dmem_n15540) );
NAND2_X1 MEM_stage_inst_dmem_U12882 ( .A1(MEM_stage_inst_dmem_n15538), .A2(MEM_stage_inst_dmem_n15537), .ZN(MEM_stage_inst_dmem_n11523) );
NAND2_X1 MEM_stage_inst_dmem_U12881 ( .A1(MEM_stage_inst_dmem_n111), .A2(MEM_stage_inst_dmem_n15554), .ZN(MEM_stage_inst_dmem_n15537) );
NAND2_X1 MEM_stage_inst_dmem_U12880 ( .A1(MEM_stage_inst_dmem_ram_1224), .A2(MEM_stage_inst_dmem_n15553), .ZN(MEM_stage_inst_dmem_n15538) );
NAND2_X1 MEM_stage_inst_dmem_U12879 ( .A1(MEM_stage_inst_dmem_n15536), .A2(MEM_stage_inst_dmem_n15535), .ZN(MEM_stage_inst_dmem_n11524) );
NAND2_X1 MEM_stage_inst_dmem_U12878 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n15554), .ZN(MEM_stage_inst_dmem_n15535) );
NAND2_X1 MEM_stage_inst_dmem_U12877 ( .A1(MEM_stage_inst_dmem_ram_1225), .A2(MEM_stage_inst_dmem_n15553), .ZN(MEM_stage_inst_dmem_n15536) );
NAND2_X1 MEM_stage_inst_dmem_U12876 ( .A1(MEM_stage_inst_dmem_n15534), .A2(MEM_stage_inst_dmem_n15533), .ZN(MEM_stage_inst_dmem_n11525) );
NAND2_X1 MEM_stage_inst_dmem_U12875 ( .A1(MEM_stage_inst_dmem_n18867), .A2(MEM_stage_inst_dmem_n15554), .ZN(MEM_stage_inst_dmem_n15533) );
NAND2_X1 MEM_stage_inst_dmem_U12874 ( .A1(MEM_stage_inst_dmem_ram_1226), .A2(MEM_stage_inst_dmem_n15553), .ZN(MEM_stage_inst_dmem_n15534) );
NAND2_X1 MEM_stage_inst_dmem_U12873 ( .A1(MEM_stage_inst_dmem_n15532), .A2(MEM_stage_inst_dmem_n15531), .ZN(MEM_stage_inst_dmem_n11526) );
NAND2_X1 MEM_stage_inst_dmem_U12872 ( .A1(MEM_stage_inst_dmem_n18864), .A2(MEM_stage_inst_dmem_n15554), .ZN(MEM_stage_inst_dmem_n15531) );
NAND2_X1 MEM_stage_inst_dmem_U12871 ( .A1(MEM_stage_inst_dmem_ram_1227), .A2(MEM_stage_inst_dmem_n15553), .ZN(MEM_stage_inst_dmem_n15532) );
NAND2_X1 MEM_stage_inst_dmem_U12870 ( .A1(MEM_stage_inst_dmem_n15530), .A2(MEM_stage_inst_dmem_n15529), .ZN(MEM_stage_inst_dmem_n11527) );
NAND2_X1 MEM_stage_inst_dmem_U12869 ( .A1(MEM_stage_inst_dmem_n18861), .A2(MEM_stage_inst_dmem_n15554), .ZN(MEM_stage_inst_dmem_n15529) );
NAND2_X1 MEM_stage_inst_dmem_U12868 ( .A1(MEM_stage_inst_dmem_ram_1228), .A2(MEM_stage_inst_dmem_n15553), .ZN(MEM_stage_inst_dmem_n15530) );
NAND2_X1 MEM_stage_inst_dmem_U12867 ( .A1(MEM_stage_inst_dmem_n15528), .A2(MEM_stage_inst_dmem_n15527), .ZN(MEM_stage_inst_dmem_n11528) );
NAND2_X1 MEM_stage_inst_dmem_U12866 ( .A1(MEM_stage_inst_dmem_n15116), .A2(MEM_stage_inst_dmem_n15554), .ZN(MEM_stage_inst_dmem_n15527) );
NAND2_X1 MEM_stage_inst_dmem_U12865 ( .A1(MEM_stage_inst_dmem_ram_1229), .A2(MEM_stage_inst_dmem_n15553), .ZN(MEM_stage_inst_dmem_n15528) );
NAND2_X1 MEM_stage_inst_dmem_U12864 ( .A1(MEM_stage_inst_dmem_n15526), .A2(MEM_stage_inst_dmem_n15525), .ZN(MEM_stage_inst_dmem_n11529) );
NAND2_X1 MEM_stage_inst_dmem_U12863 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n15554), .ZN(MEM_stage_inst_dmem_n15525) );
NAND2_X1 MEM_stage_inst_dmem_U12862 ( .A1(MEM_stage_inst_dmem_ram_1230), .A2(MEM_stage_inst_dmem_n15553), .ZN(MEM_stage_inst_dmem_n15526) );
NAND2_X1 MEM_stage_inst_dmem_U12861 ( .A1(MEM_stage_inst_dmem_n15524), .A2(MEM_stage_inst_dmem_n15523), .ZN(MEM_stage_inst_dmem_n11530) );
NAND2_X1 MEM_stage_inst_dmem_U12860 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n15554), .ZN(MEM_stage_inst_dmem_n15523) );
INV_X1 MEM_stage_inst_dmem_U12859 ( .A(MEM_stage_inst_dmem_n15553), .ZN(MEM_stage_inst_dmem_n15554) );
NAND2_X1 MEM_stage_inst_dmem_U12858 ( .A1(MEM_stage_inst_dmem_ram_1231), .A2(MEM_stage_inst_dmem_n15553), .ZN(MEM_stage_inst_dmem_n15524) );
NAND2_X1 MEM_stage_inst_dmem_U12857 ( .A1(MEM_stage_inst_dmem_n21039), .A2(MEM_stage_inst_dmem_n15931), .ZN(MEM_stage_inst_dmem_n15553) );
NAND2_X1 MEM_stage_inst_dmem_U12856 ( .A1(MEM_stage_inst_dmem_n15522), .A2(MEM_stage_inst_dmem_n15521), .ZN(MEM_stage_inst_dmem_n11531) );
NAND2_X1 MEM_stage_inst_dmem_U12855 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n15520), .ZN(MEM_stage_inst_dmem_n15521) );
NAND2_X1 MEM_stage_inst_dmem_U12854 ( .A1(MEM_stage_inst_dmem_ram_1232), .A2(MEM_stage_inst_dmem_n15519), .ZN(MEM_stage_inst_dmem_n15522) );
NAND2_X1 MEM_stage_inst_dmem_U12853 ( .A1(MEM_stage_inst_dmem_n15518), .A2(MEM_stage_inst_dmem_n15517), .ZN(MEM_stage_inst_dmem_n11532) );
NAND2_X1 MEM_stage_inst_dmem_U12852 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n15520), .ZN(MEM_stage_inst_dmem_n15517) );
NAND2_X1 MEM_stage_inst_dmem_U12851 ( .A1(MEM_stage_inst_dmem_ram_1233), .A2(MEM_stage_inst_dmem_n15519), .ZN(MEM_stage_inst_dmem_n15518) );
NAND2_X1 MEM_stage_inst_dmem_U12850 ( .A1(MEM_stage_inst_dmem_n15516), .A2(MEM_stage_inst_dmem_n15515), .ZN(MEM_stage_inst_dmem_n11533) );
NAND2_X1 MEM_stage_inst_dmem_U12849 ( .A1(MEM_stage_inst_dmem_n18887), .A2(MEM_stage_inst_dmem_n15520), .ZN(MEM_stage_inst_dmem_n15515) );
NAND2_X1 MEM_stage_inst_dmem_U12848 ( .A1(MEM_stage_inst_dmem_ram_1234), .A2(MEM_stage_inst_dmem_n15519), .ZN(MEM_stage_inst_dmem_n15516) );
NAND2_X1 MEM_stage_inst_dmem_U12847 ( .A1(MEM_stage_inst_dmem_n15514), .A2(MEM_stage_inst_dmem_n15513), .ZN(MEM_stage_inst_dmem_n11534) );
NAND2_X1 MEM_stage_inst_dmem_U12846 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n15520), .ZN(MEM_stage_inst_dmem_n15513) );
NAND2_X1 MEM_stage_inst_dmem_U12845 ( .A1(MEM_stage_inst_dmem_ram_1235), .A2(MEM_stage_inst_dmem_n15519), .ZN(MEM_stage_inst_dmem_n15514) );
NAND2_X1 MEM_stage_inst_dmem_U12844 ( .A1(MEM_stage_inst_dmem_n15512), .A2(MEM_stage_inst_dmem_n15511), .ZN(MEM_stage_inst_dmem_n11535) );
NAND2_X1 MEM_stage_inst_dmem_U12843 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n15520), .ZN(MEM_stage_inst_dmem_n15511) );
NAND2_X1 MEM_stage_inst_dmem_U12842 ( .A1(MEM_stage_inst_dmem_ram_1236), .A2(MEM_stage_inst_dmem_n15519), .ZN(MEM_stage_inst_dmem_n15512) );
NAND2_X1 MEM_stage_inst_dmem_U12841 ( .A1(MEM_stage_inst_dmem_n15510), .A2(MEM_stage_inst_dmem_n15509), .ZN(MEM_stage_inst_dmem_n11536) );
NAND2_X1 MEM_stage_inst_dmem_U12840 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n15520), .ZN(MEM_stage_inst_dmem_n15509) );
NAND2_X1 MEM_stage_inst_dmem_U12839 ( .A1(MEM_stage_inst_dmem_ram_1237), .A2(MEM_stage_inst_dmem_n15519), .ZN(MEM_stage_inst_dmem_n15510) );
NAND2_X1 MEM_stage_inst_dmem_U12838 ( .A1(MEM_stage_inst_dmem_n15508), .A2(MEM_stage_inst_dmem_n15507), .ZN(MEM_stage_inst_dmem_n11537) );
NAND2_X1 MEM_stage_inst_dmem_U12837 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n15520), .ZN(MEM_stage_inst_dmem_n15507) );
NAND2_X1 MEM_stage_inst_dmem_U12836 ( .A1(MEM_stage_inst_dmem_ram_1238), .A2(MEM_stage_inst_dmem_n15519), .ZN(MEM_stage_inst_dmem_n15508) );
NAND2_X1 MEM_stage_inst_dmem_U12835 ( .A1(MEM_stage_inst_dmem_n15506), .A2(MEM_stage_inst_dmem_n15505), .ZN(MEM_stage_inst_dmem_n11538) );
NAND2_X1 MEM_stage_inst_dmem_U12834 ( .A1(MEM_stage_inst_dmem_n18875), .A2(MEM_stage_inst_dmem_n15520), .ZN(MEM_stage_inst_dmem_n15505) );
NAND2_X1 MEM_stage_inst_dmem_U12833 ( .A1(MEM_stage_inst_dmem_ram_1239), .A2(MEM_stage_inst_dmem_n15519), .ZN(MEM_stage_inst_dmem_n15506) );
NAND2_X1 MEM_stage_inst_dmem_U12832 ( .A1(MEM_stage_inst_dmem_n15504), .A2(MEM_stage_inst_dmem_n15503), .ZN(MEM_stage_inst_dmem_n11539) );
NAND2_X1 MEM_stage_inst_dmem_U12831 ( .A1(MEM_stage_inst_dmem_n111), .A2(MEM_stage_inst_dmem_n15520), .ZN(MEM_stage_inst_dmem_n15503) );
NAND2_X1 MEM_stage_inst_dmem_U12830 ( .A1(MEM_stage_inst_dmem_ram_1240), .A2(MEM_stage_inst_dmem_n15519), .ZN(MEM_stage_inst_dmem_n15504) );
NAND2_X1 MEM_stage_inst_dmem_U12829 ( .A1(MEM_stage_inst_dmem_n15502), .A2(MEM_stage_inst_dmem_n15501), .ZN(MEM_stage_inst_dmem_n11540) );
NAND2_X1 MEM_stage_inst_dmem_U12828 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n15520), .ZN(MEM_stage_inst_dmem_n15501) );
NAND2_X1 MEM_stage_inst_dmem_U12827 ( .A1(MEM_stage_inst_dmem_ram_1241), .A2(MEM_stage_inst_dmem_n15519), .ZN(MEM_stage_inst_dmem_n15502) );
NAND2_X1 MEM_stage_inst_dmem_U12826 ( .A1(MEM_stage_inst_dmem_n15500), .A2(MEM_stage_inst_dmem_n15499), .ZN(MEM_stage_inst_dmem_n11541) );
NAND2_X1 MEM_stage_inst_dmem_U12825 ( .A1(MEM_stage_inst_dmem_n18867), .A2(MEM_stage_inst_dmem_n15520), .ZN(MEM_stage_inst_dmem_n15499) );
NAND2_X1 MEM_stage_inst_dmem_U12824 ( .A1(MEM_stage_inst_dmem_ram_1242), .A2(MEM_stage_inst_dmem_n15519), .ZN(MEM_stage_inst_dmem_n15500) );
NAND2_X1 MEM_stage_inst_dmem_U12823 ( .A1(MEM_stage_inst_dmem_n15498), .A2(MEM_stage_inst_dmem_n15497), .ZN(MEM_stage_inst_dmem_n11542) );
NAND2_X1 MEM_stage_inst_dmem_U12822 ( .A1(MEM_stage_inst_dmem_n18864), .A2(MEM_stage_inst_dmem_n15520), .ZN(MEM_stage_inst_dmem_n15497) );
NAND2_X1 MEM_stage_inst_dmem_U12821 ( .A1(MEM_stage_inst_dmem_ram_1243), .A2(MEM_stage_inst_dmem_n15519), .ZN(MEM_stage_inst_dmem_n15498) );
NAND2_X1 MEM_stage_inst_dmem_U12820 ( .A1(MEM_stage_inst_dmem_n15496), .A2(MEM_stage_inst_dmem_n15495), .ZN(MEM_stage_inst_dmem_n11543) );
NAND2_X1 MEM_stage_inst_dmem_U12819 ( .A1(MEM_stage_inst_dmem_n18861), .A2(MEM_stage_inst_dmem_n15520), .ZN(MEM_stage_inst_dmem_n15495) );
NAND2_X1 MEM_stage_inst_dmem_U12818 ( .A1(MEM_stage_inst_dmem_ram_1244), .A2(MEM_stage_inst_dmem_n15519), .ZN(MEM_stage_inst_dmem_n15496) );
NAND2_X1 MEM_stage_inst_dmem_U12817 ( .A1(MEM_stage_inst_dmem_n15494), .A2(MEM_stage_inst_dmem_n15493), .ZN(MEM_stage_inst_dmem_n11544) );
NAND2_X1 MEM_stage_inst_dmem_U12816 ( .A1(MEM_stage_inst_dmem_n19242), .A2(MEM_stage_inst_dmem_n15520), .ZN(MEM_stage_inst_dmem_n15493) );
NAND2_X1 MEM_stage_inst_dmem_U12815 ( .A1(MEM_stage_inst_dmem_ram_1245), .A2(MEM_stage_inst_dmem_n15519), .ZN(MEM_stage_inst_dmem_n15494) );
NAND2_X1 MEM_stage_inst_dmem_U12814 ( .A1(MEM_stage_inst_dmem_n15492), .A2(MEM_stage_inst_dmem_n15491), .ZN(MEM_stage_inst_dmem_n11545) );
NAND2_X1 MEM_stage_inst_dmem_U12813 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n15520), .ZN(MEM_stage_inst_dmem_n15491) );
NAND2_X1 MEM_stage_inst_dmem_U12812 ( .A1(MEM_stage_inst_dmem_ram_1246), .A2(MEM_stage_inst_dmem_n15519), .ZN(MEM_stage_inst_dmem_n15492) );
NAND2_X1 MEM_stage_inst_dmem_U12811 ( .A1(MEM_stage_inst_dmem_n15490), .A2(MEM_stage_inst_dmem_n15489), .ZN(MEM_stage_inst_dmem_n11546) );
NAND2_X1 MEM_stage_inst_dmem_U12810 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n15520), .ZN(MEM_stage_inst_dmem_n15489) );
INV_X1 MEM_stage_inst_dmem_U12809 ( .A(MEM_stage_inst_dmem_n15519), .ZN(MEM_stage_inst_dmem_n15520) );
NAND2_X1 MEM_stage_inst_dmem_U12808 ( .A1(MEM_stage_inst_dmem_ram_1247), .A2(MEM_stage_inst_dmem_n15519), .ZN(MEM_stage_inst_dmem_n15490) );
NAND2_X1 MEM_stage_inst_dmem_U12807 ( .A1(MEM_stage_inst_dmem_n21004), .A2(MEM_stage_inst_dmem_n15931), .ZN(MEM_stage_inst_dmem_n15519) );
NAND2_X1 MEM_stage_inst_dmem_U12806 ( .A1(MEM_stage_inst_dmem_n15488), .A2(MEM_stage_inst_dmem_n15487), .ZN(MEM_stage_inst_dmem_n11547) );
NAND2_X1 MEM_stage_inst_dmem_U12805 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n15486), .ZN(MEM_stage_inst_dmem_n15487) );
NAND2_X1 MEM_stage_inst_dmem_U12804 ( .A1(MEM_stage_inst_dmem_ram_1248), .A2(MEM_stage_inst_dmem_n15485), .ZN(MEM_stage_inst_dmem_n15488) );
NAND2_X1 MEM_stage_inst_dmem_U12803 ( .A1(MEM_stage_inst_dmem_n15484), .A2(MEM_stage_inst_dmem_n15483), .ZN(MEM_stage_inst_dmem_n11548) );
NAND2_X1 MEM_stage_inst_dmem_U12802 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n15486), .ZN(MEM_stage_inst_dmem_n15483) );
NAND2_X1 MEM_stage_inst_dmem_U12801 ( .A1(MEM_stage_inst_dmem_ram_1249), .A2(MEM_stage_inst_dmem_n15485), .ZN(MEM_stage_inst_dmem_n15484) );
NAND2_X1 MEM_stage_inst_dmem_U12800 ( .A1(MEM_stage_inst_dmem_n15482), .A2(MEM_stage_inst_dmem_n15481), .ZN(MEM_stage_inst_dmem_n11549) );
NAND2_X1 MEM_stage_inst_dmem_U12799 ( .A1(MEM_stage_inst_dmem_n18887), .A2(MEM_stage_inst_dmem_n15486), .ZN(MEM_stage_inst_dmem_n15481) );
NAND2_X1 MEM_stage_inst_dmem_U12798 ( .A1(MEM_stage_inst_dmem_ram_1250), .A2(MEM_stage_inst_dmem_n15485), .ZN(MEM_stage_inst_dmem_n15482) );
NAND2_X1 MEM_stage_inst_dmem_U12797 ( .A1(MEM_stage_inst_dmem_n15480), .A2(MEM_stage_inst_dmem_n15479), .ZN(MEM_stage_inst_dmem_n11550) );
NAND2_X1 MEM_stage_inst_dmem_U12796 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n15486), .ZN(MEM_stage_inst_dmem_n15479) );
NAND2_X1 MEM_stage_inst_dmem_U12795 ( .A1(MEM_stage_inst_dmem_ram_1251), .A2(MEM_stage_inst_dmem_n15485), .ZN(MEM_stage_inst_dmem_n15480) );
NAND2_X1 MEM_stage_inst_dmem_U12794 ( .A1(MEM_stage_inst_dmem_n15478), .A2(MEM_stage_inst_dmem_n15477), .ZN(MEM_stage_inst_dmem_n11551) );
NAND2_X1 MEM_stage_inst_dmem_U12793 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n15486), .ZN(MEM_stage_inst_dmem_n15477) );
NAND2_X1 MEM_stage_inst_dmem_U12792 ( .A1(MEM_stage_inst_dmem_ram_1252), .A2(MEM_stage_inst_dmem_n15485), .ZN(MEM_stage_inst_dmem_n15478) );
NAND2_X1 MEM_stage_inst_dmem_U12791 ( .A1(MEM_stage_inst_dmem_n15476), .A2(MEM_stage_inst_dmem_n15475), .ZN(MEM_stage_inst_dmem_n11552) );
NAND2_X1 MEM_stage_inst_dmem_U12790 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n15486), .ZN(MEM_stage_inst_dmem_n15475) );
NAND2_X1 MEM_stage_inst_dmem_U12789 ( .A1(MEM_stage_inst_dmem_ram_1253), .A2(MEM_stage_inst_dmem_n15485), .ZN(MEM_stage_inst_dmem_n15476) );
NAND2_X1 MEM_stage_inst_dmem_U12788 ( .A1(MEM_stage_inst_dmem_n15474), .A2(MEM_stage_inst_dmem_n15473), .ZN(MEM_stage_inst_dmem_n11553) );
NAND2_X1 MEM_stage_inst_dmem_U12787 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n15486), .ZN(MEM_stage_inst_dmem_n15473) );
NAND2_X1 MEM_stage_inst_dmem_U12786 ( .A1(MEM_stage_inst_dmem_ram_1254), .A2(MEM_stage_inst_dmem_n15485), .ZN(MEM_stage_inst_dmem_n15474) );
NAND2_X1 MEM_stage_inst_dmem_U12785 ( .A1(MEM_stage_inst_dmem_n15472), .A2(MEM_stage_inst_dmem_n15471), .ZN(MEM_stage_inst_dmem_n11554) );
NAND2_X1 MEM_stage_inst_dmem_U12784 ( .A1(MEM_stage_inst_dmem_n18875), .A2(MEM_stage_inst_dmem_n15486), .ZN(MEM_stage_inst_dmem_n15471) );
NAND2_X1 MEM_stage_inst_dmem_U12783 ( .A1(MEM_stage_inst_dmem_ram_1255), .A2(MEM_stage_inst_dmem_n15485), .ZN(MEM_stage_inst_dmem_n15472) );
NAND2_X1 MEM_stage_inst_dmem_U12782 ( .A1(MEM_stage_inst_dmem_n15470), .A2(MEM_stage_inst_dmem_n15469), .ZN(MEM_stage_inst_dmem_n11555) );
NAND2_X1 MEM_stage_inst_dmem_U12781 ( .A1(MEM_stage_inst_dmem_n111), .A2(MEM_stage_inst_dmem_n15486), .ZN(MEM_stage_inst_dmem_n15469) );
NAND2_X1 MEM_stage_inst_dmem_U12780 ( .A1(MEM_stage_inst_dmem_ram_1256), .A2(MEM_stage_inst_dmem_n15485), .ZN(MEM_stage_inst_dmem_n15470) );
NAND2_X1 MEM_stage_inst_dmem_U12779 ( .A1(MEM_stage_inst_dmem_n15468), .A2(MEM_stage_inst_dmem_n15467), .ZN(MEM_stage_inst_dmem_n11556) );
NAND2_X1 MEM_stage_inst_dmem_U12778 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n15486), .ZN(MEM_stage_inst_dmem_n15467) );
NAND2_X1 MEM_stage_inst_dmem_U12777 ( .A1(MEM_stage_inst_dmem_ram_1257), .A2(MEM_stage_inst_dmem_n15485), .ZN(MEM_stage_inst_dmem_n15468) );
NAND2_X1 MEM_stage_inst_dmem_U12776 ( .A1(MEM_stage_inst_dmem_n15466), .A2(MEM_stage_inst_dmem_n15465), .ZN(MEM_stage_inst_dmem_n11557) );
NAND2_X1 MEM_stage_inst_dmem_U12775 ( .A1(MEM_stage_inst_dmem_n18867), .A2(MEM_stage_inst_dmem_n15486), .ZN(MEM_stage_inst_dmem_n15465) );
NAND2_X1 MEM_stage_inst_dmem_U12774 ( .A1(MEM_stage_inst_dmem_ram_1258), .A2(MEM_stage_inst_dmem_n15485), .ZN(MEM_stage_inst_dmem_n15466) );
NAND2_X1 MEM_stage_inst_dmem_U12773 ( .A1(MEM_stage_inst_dmem_n15464), .A2(MEM_stage_inst_dmem_n15463), .ZN(MEM_stage_inst_dmem_n11558) );
NAND2_X1 MEM_stage_inst_dmem_U12772 ( .A1(MEM_stage_inst_dmem_n18864), .A2(MEM_stage_inst_dmem_n15486), .ZN(MEM_stage_inst_dmem_n15463) );
NAND2_X1 MEM_stage_inst_dmem_U12771 ( .A1(MEM_stage_inst_dmem_ram_1259), .A2(MEM_stage_inst_dmem_n15485), .ZN(MEM_stage_inst_dmem_n15464) );
NAND2_X1 MEM_stage_inst_dmem_U12770 ( .A1(MEM_stage_inst_dmem_n15462), .A2(MEM_stage_inst_dmem_n15461), .ZN(MEM_stage_inst_dmem_n11559) );
NAND2_X1 MEM_stage_inst_dmem_U12769 ( .A1(MEM_stage_inst_dmem_n18861), .A2(MEM_stage_inst_dmem_n15486), .ZN(MEM_stage_inst_dmem_n15461) );
NAND2_X1 MEM_stage_inst_dmem_U12768 ( .A1(MEM_stage_inst_dmem_ram_1260), .A2(MEM_stage_inst_dmem_n15485), .ZN(MEM_stage_inst_dmem_n15462) );
NAND2_X1 MEM_stage_inst_dmem_U12767 ( .A1(MEM_stage_inst_dmem_n15460), .A2(MEM_stage_inst_dmem_n15459), .ZN(MEM_stage_inst_dmem_n11560) );
NAND2_X1 MEM_stage_inst_dmem_U12766 ( .A1(MEM_stage_inst_dmem_n20512), .A2(MEM_stage_inst_dmem_n15486), .ZN(MEM_stage_inst_dmem_n15459) );
NAND2_X1 MEM_stage_inst_dmem_U12765 ( .A1(MEM_stage_inst_dmem_ram_1261), .A2(MEM_stage_inst_dmem_n15485), .ZN(MEM_stage_inst_dmem_n15460) );
NAND2_X1 MEM_stage_inst_dmem_U12764 ( .A1(MEM_stage_inst_dmem_n15458), .A2(MEM_stage_inst_dmem_n15457), .ZN(MEM_stage_inst_dmem_n11561) );
NAND2_X1 MEM_stage_inst_dmem_U12763 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n15486), .ZN(MEM_stage_inst_dmem_n15457) );
NAND2_X1 MEM_stage_inst_dmem_U12762 ( .A1(MEM_stage_inst_dmem_ram_1262), .A2(MEM_stage_inst_dmem_n15485), .ZN(MEM_stage_inst_dmem_n15458) );
NAND2_X1 MEM_stage_inst_dmem_U12761 ( .A1(MEM_stage_inst_dmem_n15456), .A2(MEM_stage_inst_dmem_n15455), .ZN(MEM_stage_inst_dmem_n11562) );
NAND2_X1 MEM_stage_inst_dmem_U12760 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n15486), .ZN(MEM_stage_inst_dmem_n15455) );
INV_X1 MEM_stage_inst_dmem_U12759 ( .A(MEM_stage_inst_dmem_n15485), .ZN(MEM_stage_inst_dmem_n15486) );
NAND2_X1 MEM_stage_inst_dmem_U12758 ( .A1(MEM_stage_inst_dmem_ram_1263), .A2(MEM_stage_inst_dmem_n15485), .ZN(MEM_stage_inst_dmem_n15456) );
NAND2_X1 MEM_stage_inst_dmem_U12757 ( .A1(MEM_stage_inst_dmem_n20969), .A2(MEM_stage_inst_dmem_n15931), .ZN(MEM_stage_inst_dmem_n15485) );
NAND2_X1 MEM_stage_inst_dmem_U12756 ( .A1(MEM_stage_inst_dmem_n15454), .A2(MEM_stage_inst_dmem_n15453), .ZN(MEM_stage_inst_dmem_n11563) );
NAND2_X1 MEM_stage_inst_dmem_U12755 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n15452), .ZN(MEM_stage_inst_dmem_n15453) );
NAND2_X1 MEM_stage_inst_dmem_U12754 ( .A1(MEM_stage_inst_dmem_ram_1264), .A2(MEM_stage_inst_dmem_n15451), .ZN(MEM_stage_inst_dmem_n15454) );
NAND2_X1 MEM_stage_inst_dmem_U12753 ( .A1(MEM_stage_inst_dmem_n15450), .A2(MEM_stage_inst_dmem_n15449), .ZN(MEM_stage_inst_dmem_n11564) );
NAND2_X1 MEM_stage_inst_dmem_U12752 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n15452), .ZN(MEM_stage_inst_dmem_n15449) );
NAND2_X1 MEM_stage_inst_dmem_U12751 ( .A1(MEM_stage_inst_dmem_ram_1265), .A2(MEM_stage_inst_dmem_n15451), .ZN(MEM_stage_inst_dmem_n15450) );
NAND2_X1 MEM_stage_inst_dmem_U12750 ( .A1(MEM_stage_inst_dmem_n15448), .A2(MEM_stage_inst_dmem_n15447), .ZN(MEM_stage_inst_dmem_n11565) );
NAND2_X1 MEM_stage_inst_dmem_U12749 ( .A1(MEM_stage_inst_dmem_n18887), .A2(MEM_stage_inst_dmem_n15452), .ZN(MEM_stage_inst_dmem_n15447) );
NAND2_X1 MEM_stage_inst_dmem_U12748 ( .A1(MEM_stage_inst_dmem_ram_1266), .A2(MEM_stage_inst_dmem_n15451), .ZN(MEM_stage_inst_dmem_n15448) );
NAND2_X1 MEM_stage_inst_dmem_U12747 ( .A1(MEM_stage_inst_dmem_n15446), .A2(MEM_stage_inst_dmem_n15445), .ZN(MEM_stage_inst_dmem_n11566) );
NAND2_X1 MEM_stage_inst_dmem_U12746 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n15452), .ZN(MEM_stage_inst_dmem_n15445) );
NAND2_X1 MEM_stage_inst_dmem_U12745 ( .A1(MEM_stage_inst_dmem_ram_1267), .A2(MEM_stage_inst_dmem_n15451), .ZN(MEM_stage_inst_dmem_n15446) );
NAND2_X1 MEM_stage_inst_dmem_U12744 ( .A1(MEM_stage_inst_dmem_n15444), .A2(MEM_stage_inst_dmem_n15443), .ZN(MEM_stage_inst_dmem_n11567) );
NAND2_X1 MEM_stage_inst_dmem_U12743 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n15452), .ZN(MEM_stage_inst_dmem_n15443) );
NAND2_X1 MEM_stage_inst_dmem_U12742 ( .A1(MEM_stage_inst_dmem_ram_1268), .A2(MEM_stage_inst_dmem_n15451), .ZN(MEM_stage_inst_dmem_n15444) );
NAND2_X1 MEM_stage_inst_dmem_U12741 ( .A1(MEM_stage_inst_dmem_n15442), .A2(MEM_stage_inst_dmem_n15441), .ZN(MEM_stage_inst_dmem_n11568) );
NAND2_X1 MEM_stage_inst_dmem_U12740 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n15452), .ZN(MEM_stage_inst_dmem_n15441) );
NAND2_X1 MEM_stage_inst_dmem_U12739 ( .A1(MEM_stage_inst_dmem_ram_1269), .A2(MEM_stage_inst_dmem_n15451), .ZN(MEM_stage_inst_dmem_n15442) );
NAND2_X1 MEM_stage_inst_dmem_U12738 ( .A1(MEM_stage_inst_dmem_n15440), .A2(MEM_stage_inst_dmem_n15439), .ZN(MEM_stage_inst_dmem_n11569) );
NAND2_X1 MEM_stage_inst_dmem_U12737 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n15452), .ZN(MEM_stage_inst_dmem_n15439) );
NAND2_X1 MEM_stage_inst_dmem_U12736 ( .A1(MEM_stage_inst_dmem_ram_1270), .A2(MEM_stage_inst_dmem_n15451), .ZN(MEM_stage_inst_dmem_n15440) );
NAND2_X1 MEM_stage_inst_dmem_U12735 ( .A1(MEM_stage_inst_dmem_n15438), .A2(MEM_stage_inst_dmem_n15437), .ZN(MEM_stage_inst_dmem_n11570) );
NAND2_X1 MEM_stage_inst_dmem_U12734 ( .A1(MEM_stage_inst_dmem_n18875), .A2(MEM_stage_inst_dmem_n15452), .ZN(MEM_stage_inst_dmem_n15437) );
NAND2_X1 MEM_stage_inst_dmem_U12733 ( .A1(MEM_stage_inst_dmem_ram_1271), .A2(MEM_stage_inst_dmem_n15451), .ZN(MEM_stage_inst_dmem_n15438) );
NAND2_X1 MEM_stage_inst_dmem_U12732 ( .A1(MEM_stage_inst_dmem_n15436), .A2(MEM_stage_inst_dmem_n15435), .ZN(MEM_stage_inst_dmem_n11571) );
NAND2_X1 MEM_stage_inst_dmem_U12731 ( .A1(MEM_stage_inst_dmem_n111), .A2(MEM_stage_inst_dmem_n15452), .ZN(MEM_stage_inst_dmem_n15435) );
NAND2_X1 MEM_stage_inst_dmem_U12730 ( .A1(MEM_stage_inst_dmem_ram_1272), .A2(MEM_stage_inst_dmem_n15451), .ZN(MEM_stage_inst_dmem_n15436) );
NAND2_X1 MEM_stage_inst_dmem_U12729 ( .A1(MEM_stage_inst_dmem_n15434), .A2(MEM_stage_inst_dmem_n15433), .ZN(MEM_stage_inst_dmem_n11572) );
NAND2_X1 MEM_stage_inst_dmem_U12728 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n15452), .ZN(MEM_stage_inst_dmem_n15433) );
NAND2_X1 MEM_stage_inst_dmem_U12727 ( .A1(MEM_stage_inst_dmem_ram_1273), .A2(MEM_stage_inst_dmem_n15451), .ZN(MEM_stage_inst_dmem_n15434) );
NAND2_X1 MEM_stage_inst_dmem_U12726 ( .A1(MEM_stage_inst_dmem_n15432), .A2(MEM_stage_inst_dmem_n15431), .ZN(MEM_stage_inst_dmem_n11573) );
NAND2_X1 MEM_stage_inst_dmem_U12725 ( .A1(MEM_stage_inst_dmem_n18867), .A2(MEM_stage_inst_dmem_n15452), .ZN(MEM_stage_inst_dmem_n15431) );
NAND2_X1 MEM_stage_inst_dmem_U12724 ( .A1(MEM_stage_inst_dmem_ram_1274), .A2(MEM_stage_inst_dmem_n15451), .ZN(MEM_stage_inst_dmem_n15432) );
NAND2_X1 MEM_stage_inst_dmem_U12723 ( .A1(MEM_stage_inst_dmem_n15430), .A2(MEM_stage_inst_dmem_n15429), .ZN(MEM_stage_inst_dmem_n11574) );
NAND2_X1 MEM_stage_inst_dmem_U12722 ( .A1(MEM_stage_inst_dmem_n18864), .A2(MEM_stage_inst_dmem_n15452), .ZN(MEM_stage_inst_dmem_n15429) );
NAND2_X1 MEM_stage_inst_dmem_U12721 ( .A1(MEM_stage_inst_dmem_ram_1275), .A2(MEM_stage_inst_dmem_n15451), .ZN(MEM_stage_inst_dmem_n15430) );
NAND2_X1 MEM_stage_inst_dmem_U12720 ( .A1(MEM_stage_inst_dmem_n15428), .A2(MEM_stage_inst_dmem_n15427), .ZN(MEM_stage_inst_dmem_n11575) );
NAND2_X1 MEM_stage_inst_dmem_U12719 ( .A1(MEM_stage_inst_dmem_n18861), .A2(MEM_stage_inst_dmem_n15452), .ZN(MEM_stage_inst_dmem_n15427) );
NAND2_X1 MEM_stage_inst_dmem_U12718 ( .A1(MEM_stage_inst_dmem_ram_1276), .A2(MEM_stage_inst_dmem_n15451), .ZN(MEM_stage_inst_dmem_n15428) );
NAND2_X1 MEM_stage_inst_dmem_U12717 ( .A1(MEM_stage_inst_dmem_n15426), .A2(MEM_stage_inst_dmem_n15425), .ZN(MEM_stage_inst_dmem_n11576) );
NAND2_X1 MEM_stage_inst_dmem_U12716 ( .A1(EX_pipeline_reg_out_18), .A2(MEM_stage_inst_dmem_n15452), .ZN(MEM_stage_inst_dmem_n15425) );
NAND2_X1 MEM_stage_inst_dmem_U12715 ( .A1(MEM_stage_inst_dmem_ram_1277), .A2(MEM_stage_inst_dmem_n15451), .ZN(MEM_stage_inst_dmem_n15426) );
NAND2_X1 MEM_stage_inst_dmem_U12714 ( .A1(MEM_stage_inst_dmem_n15424), .A2(MEM_stage_inst_dmem_n15423), .ZN(MEM_stage_inst_dmem_n11577) );
NAND2_X1 MEM_stage_inst_dmem_U12713 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n15452), .ZN(MEM_stage_inst_dmem_n15423) );
NAND2_X1 MEM_stage_inst_dmem_U12712 ( .A1(MEM_stage_inst_dmem_ram_1278), .A2(MEM_stage_inst_dmem_n15451), .ZN(MEM_stage_inst_dmem_n15424) );
NAND2_X1 MEM_stage_inst_dmem_U12711 ( .A1(MEM_stage_inst_dmem_n15422), .A2(MEM_stage_inst_dmem_n15421), .ZN(MEM_stage_inst_dmem_n11578) );
NAND2_X1 MEM_stage_inst_dmem_U12710 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n15452), .ZN(MEM_stage_inst_dmem_n15421) );
NAND2_X1 MEM_stage_inst_dmem_U12709 ( .A1(MEM_stage_inst_dmem_ram_1279), .A2(MEM_stage_inst_dmem_n15451), .ZN(MEM_stage_inst_dmem_n15422) );
NAND2_X1 MEM_stage_inst_dmem_U12708 ( .A1(MEM_stage_inst_dmem_n20934), .A2(MEM_stage_inst_dmem_n15931), .ZN(MEM_stage_inst_dmem_n15451) );
NOR2_X2 MEM_stage_inst_dmem_U12707 ( .A1(MEM_stage_inst_dmem_n16519), .A2(MEM_stage_inst_dmem_n19823), .ZN(MEM_stage_inst_dmem_n15931) );
NAND2_X1 MEM_stage_inst_dmem_U12706 ( .A1(MEM_stage_inst_dmem_n15420), .A2(MEM_stage_inst_dmem_n15419), .ZN(MEM_stage_inst_dmem_n11579) );
NAND2_X1 MEM_stage_inst_dmem_U12705 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n15418), .ZN(MEM_stage_inst_dmem_n15419) );
NAND2_X1 MEM_stage_inst_dmem_U12704 ( .A1(MEM_stage_inst_dmem_ram_1280), .A2(MEM_stage_inst_dmem_n15417), .ZN(MEM_stage_inst_dmem_n15420) );
NAND2_X1 MEM_stage_inst_dmem_U12703 ( .A1(MEM_stage_inst_dmem_n15416), .A2(MEM_stage_inst_dmem_n15415), .ZN(MEM_stage_inst_dmem_n11580) );
NAND2_X1 MEM_stage_inst_dmem_U12702 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n15418), .ZN(MEM_stage_inst_dmem_n15415) );
NAND2_X1 MEM_stage_inst_dmem_U12701 ( .A1(MEM_stage_inst_dmem_ram_1281), .A2(MEM_stage_inst_dmem_n15417), .ZN(MEM_stage_inst_dmem_n15416) );
NAND2_X1 MEM_stage_inst_dmem_U12700 ( .A1(MEM_stage_inst_dmem_n15414), .A2(MEM_stage_inst_dmem_n15413), .ZN(MEM_stage_inst_dmem_n11581) );
NAND2_X1 MEM_stage_inst_dmem_U12699 ( .A1(MEM_stage_inst_dmem_n18887), .A2(MEM_stage_inst_dmem_n15418), .ZN(MEM_stage_inst_dmem_n15413) );
NAND2_X1 MEM_stage_inst_dmem_U12698 ( .A1(MEM_stage_inst_dmem_ram_1282), .A2(MEM_stage_inst_dmem_n15417), .ZN(MEM_stage_inst_dmem_n15414) );
NAND2_X1 MEM_stage_inst_dmem_U12697 ( .A1(MEM_stage_inst_dmem_n15412), .A2(MEM_stage_inst_dmem_n15411), .ZN(MEM_stage_inst_dmem_n11582) );
NAND2_X1 MEM_stage_inst_dmem_U12696 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n15418), .ZN(MEM_stage_inst_dmem_n15411) );
NAND2_X1 MEM_stage_inst_dmem_U12695 ( .A1(MEM_stage_inst_dmem_ram_1283), .A2(MEM_stage_inst_dmem_n15417), .ZN(MEM_stage_inst_dmem_n15412) );
NAND2_X1 MEM_stage_inst_dmem_U12694 ( .A1(MEM_stage_inst_dmem_n15410), .A2(MEM_stage_inst_dmem_n15409), .ZN(MEM_stage_inst_dmem_n11583) );
NAND2_X1 MEM_stage_inst_dmem_U12693 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n15418), .ZN(MEM_stage_inst_dmem_n15409) );
NAND2_X1 MEM_stage_inst_dmem_U12692 ( .A1(MEM_stage_inst_dmem_ram_1284), .A2(MEM_stage_inst_dmem_n15417), .ZN(MEM_stage_inst_dmem_n15410) );
NAND2_X1 MEM_stage_inst_dmem_U12691 ( .A1(MEM_stage_inst_dmem_n15408), .A2(MEM_stage_inst_dmem_n15407), .ZN(MEM_stage_inst_dmem_n11584) );
NAND2_X1 MEM_stage_inst_dmem_U12690 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n15418), .ZN(MEM_stage_inst_dmem_n15407) );
NAND2_X1 MEM_stage_inst_dmem_U12689 ( .A1(MEM_stage_inst_dmem_ram_1285), .A2(MEM_stage_inst_dmem_n15417), .ZN(MEM_stage_inst_dmem_n15408) );
NAND2_X1 MEM_stage_inst_dmem_U12688 ( .A1(MEM_stage_inst_dmem_n15406), .A2(MEM_stage_inst_dmem_n15405), .ZN(MEM_stage_inst_dmem_n11585) );
NAND2_X1 MEM_stage_inst_dmem_U12687 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n15418), .ZN(MEM_stage_inst_dmem_n15405) );
NAND2_X1 MEM_stage_inst_dmem_U12686 ( .A1(MEM_stage_inst_dmem_ram_1286), .A2(MEM_stage_inst_dmem_n15417), .ZN(MEM_stage_inst_dmem_n15406) );
NAND2_X1 MEM_stage_inst_dmem_U12685 ( .A1(MEM_stage_inst_dmem_n15404), .A2(MEM_stage_inst_dmem_n15403), .ZN(MEM_stage_inst_dmem_n11586) );
NAND2_X1 MEM_stage_inst_dmem_U12684 ( .A1(MEM_stage_inst_dmem_n18875), .A2(MEM_stage_inst_dmem_n15418), .ZN(MEM_stage_inst_dmem_n15403) );
NAND2_X1 MEM_stage_inst_dmem_U12683 ( .A1(MEM_stage_inst_dmem_ram_1287), .A2(MEM_stage_inst_dmem_n15417), .ZN(MEM_stage_inst_dmem_n15404) );
NAND2_X1 MEM_stage_inst_dmem_U12682 ( .A1(MEM_stage_inst_dmem_n15402), .A2(MEM_stage_inst_dmem_n15401), .ZN(MEM_stage_inst_dmem_n11587) );
NAND2_X1 MEM_stage_inst_dmem_U12681 ( .A1(MEM_stage_inst_dmem_n111), .A2(MEM_stage_inst_dmem_n15418), .ZN(MEM_stage_inst_dmem_n15401) );
NAND2_X1 MEM_stage_inst_dmem_U12680 ( .A1(MEM_stage_inst_dmem_ram_1288), .A2(MEM_stage_inst_dmem_n15417), .ZN(MEM_stage_inst_dmem_n15402) );
NAND2_X1 MEM_stage_inst_dmem_U12679 ( .A1(MEM_stage_inst_dmem_n15400), .A2(MEM_stage_inst_dmem_n15399), .ZN(MEM_stage_inst_dmem_n11588) );
NAND2_X1 MEM_stage_inst_dmem_U12678 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n15418), .ZN(MEM_stage_inst_dmem_n15399) );
NAND2_X1 MEM_stage_inst_dmem_U12677 ( .A1(MEM_stage_inst_dmem_ram_1289), .A2(MEM_stage_inst_dmem_n15417), .ZN(MEM_stage_inst_dmem_n15400) );
NAND2_X1 MEM_stage_inst_dmem_U12676 ( .A1(MEM_stage_inst_dmem_n15398), .A2(MEM_stage_inst_dmem_n15397), .ZN(MEM_stage_inst_dmem_n11589) );
NAND2_X1 MEM_stage_inst_dmem_U12675 ( .A1(MEM_stage_inst_dmem_n18867), .A2(MEM_stage_inst_dmem_n15418), .ZN(MEM_stage_inst_dmem_n15397) );
NAND2_X1 MEM_stage_inst_dmem_U12674 ( .A1(MEM_stage_inst_dmem_ram_1290), .A2(MEM_stage_inst_dmem_n15417), .ZN(MEM_stage_inst_dmem_n15398) );
NAND2_X1 MEM_stage_inst_dmem_U12673 ( .A1(MEM_stage_inst_dmem_n15396), .A2(MEM_stage_inst_dmem_n15395), .ZN(MEM_stage_inst_dmem_n11590) );
NAND2_X1 MEM_stage_inst_dmem_U12672 ( .A1(MEM_stage_inst_dmem_n18864), .A2(MEM_stage_inst_dmem_n15418), .ZN(MEM_stage_inst_dmem_n15395) );
NAND2_X1 MEM_stage_inst_dmem_U12671 ( .A1(MEM_stage_inst_dmem_ram_1291), .A2(MEM_stage_inst_dmem_n15417), .ZN(MEM_stage_inst_dmem_n15396) );
NAND2_X1 MEM_stage_inst_dmem_U12670 ( .A1(MEM_stage_inst_dmem_n15394), .A2(MEM_stage_inst_dmem_n15393), .ZN(MEM_stage_inst_dmem_n11591) );
NAND2_X1 MEM_stage_inst_dmem_U12669 ( .A1(MEM_stage_inst_dmem_n18861), .A2(MEM_stage_inst_dmem_n15418), .ZN(MEM_stage_inst_dmem_n15393) );
NAND2_X1 MEM_stage_inst_dmem_U12668 ( .A1(MEM_stage_inst_dmem_ram_1292), .A2(MEM_stage_inst_dmem_n15417), .ZN(MEM_stage_inst_dmem_n15394) );
NAND2_X1 MEM_stage_inst_dmem_U12667 ( .A1(MEM_stage_inst_dmem_n15392), .A2(MEM_stage_inst_dmem_n15391), .ZN(MEM_stage_inst_dmem_n11592) );
NAND2_X1 MEM_stage_inst_dmem_U12666 ( .A1(MEM_stage_inst_dmem_n116), .A2(MEM_stage_inst_dmem_n15418), .ZN(MEM_stage_inst_dmem_n15391) );
NAND2_X1 MEM_stage_inst_dmem_U12665 ( .A1(MEM_stage_inst_dmem_ram_1293), .A2(MEM_stage_inst_dmem_n15417), .ZN(MEM_stage_inst_dmem_n15392) );
NAND2_X1 MEM_stage_inst_dmem_U12664 ( .A1(MEM_stage_inst_dmem_n15390), .A2(MEM_stage_inst_dmem_n15389), .ZN(MEM_stage_inst_dmem_n11593) );
NAND2_X1 MEM_stage_inst_dmem_U12663 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n15418), .ZN(MEM_stage_inst_dmem_n15389) );
NAND2_X1 MEM_stage_inst_dmem_U12662 ( .A1(MEM_stage_inst_dmem_ram_1294), .A2(MEM_stage_inst_dmem_n15417), .ZN(MEM_stage_inst_dmem_n15390) );
NAND2_X1 MEM_stage_inst_dmem_U12661 ( .A1(MEM_stage_inst_dmem_n15388), .A2(MEM_stage_inst_dmem_n15387), .ZN(MEM_stage_inst_dmem_n11594) );
NAND2_X1 MEM_stage_inst_dmem_U12660 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n15418), .ZN(MEM_stage_inst_dmem_n15387) );
INV_X1 MEM_stage_inst_dmem_U12659 ( .A(MEM_stage_inst_dmem_n15417), .ZN(MEM_stage_inst_dmem_n15418) );
NAND2_X1 MEM_stage_inst_dmem_U12658 ( .A1(MEM_stage_inst_dmem_ram_1295), .A2(MEM_stage_inst_dmem_n15417), .ZN(MEM_stage_inst_dmem_n15388) );
NAND2_X1 MEM_stage_inst_dmem_U12657 ( .A1(MEM_stage_inst_dmem_n21465), .A2(MEM_stage_inst_dmem_n15386), .ZN(MEM_stage_inst_dmem_n15417) );
NAND2_X1 MEM_stage_inst_dmem_U12656 ( .A1(MEM_stage_inst_dmem_n15385), .A2(MEM_stage_inst_dmem_n15384), .ZN(MEM_stage_inst_dmem_n11595) );
NAND2_X1 MEM_stage_inst_dmem_U12655 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n15383), .ZN(MEM_stage_inst_dmem_n15384) );
NAND2_X1 MEM_stage_inst_dmem_U12654 ( .A1(MEM_stage_inst_dmem_ram_1296), .A2(MEM_stage_inst_dmem_n15382), .ZN(MEM_stage_inst_dmem_n15385) );
NAND2_X1 MEM_stage_inst_dmem_U12653 ( .A1(MEM_stage_inst_dmem_n15381), .A2(MEM_stage_inst_dmem_n15380), .ZN(MEM_stage_inst_dmem_n11596) );
NAND2_X1 MEM_stage_inst_dmem_U12652 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n15383), .ZN(MEM_stage_inst_dmem_n15380) );
NAND2_X1 MEM_stage_inst_dmem_U12651 ( .A1(MEM_stage_inst_dmem_ram_1297), .A2(MEM_stage_inst_dmem_n15382), .ZN(MEM_stage_inst_dmem_n15381) );
NAND2_X1 MEM_stage_inst_dmem_U12650 ( .A1(MEM_stage_inst_dmem_n15379), .A2(MEM_stage_inst_dmem_n15378), .ZN(MEM_stage_inst_dmem_n11597) );
NAND2_X1 MEM_stage_inst_dmem_U12649 ( .A1(MEM_stage_inst_dmem_n18887), .A2(MEM_stage_inst_dmem_n15383), .ZN(MEM_stage_inst_dmem_n15378) );
NAND2_X1 MEM_stage_inst_dmem_U12648 ( .A1(MEM_stage_inst_dmem_ram_1298), .A2(MEM_stage_inst_dmem_n15382), .ZN(MEM_stage_inst_dmem_n15379) );
NAND2_X1 MEM_stage_inst_dmem_U12647 ( .A1(MEM_stage_inst_dmem_n15377), .A2(MEM_stage_inst_dmem_n15376), .ZN(MEM_stage_inst_dmem_n11598) );
NAND2_X1 MEM_stage_inst_dmem_U12646 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n15383), .ZN(MEM_stage_inst_dmem_n15376) );
NAND2_X1 MEM_stage_inst_dmem_U12645 ( .A1(MEM_stage_inst_dmem_ram_1299), .A2(MEM_stage_inst_dmem_n15382), .ZN(MEM_stage_inst_dmem_n15377) );
NAND2_X1 MEM_stage_inst_dmem_U12644 ( .A1(MEM_stage_inst_dmem_n15375), .A2(MEM_stage_inst_dmem_n15374), .ZN(MEM_stage_inst_dmem_n11599) );
NAND2_X1 MEM_stage_inst_dmem_U12643 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n15383), .ZN(MEM_stage_inst_dmem_n15374) );
NAND2_X1 MEM_stage_inst_dmem_U12642 ( .A1(MEM_stage_inst_dmem_ram_1300), .A2(MEM_stage_inst_dmem_n15382), .ZN(MEM_stage_inst_dmem_n15375) );
NAND2_X1 MEM_stage_inst_dmem_U12641 ( .A1(MEM_stage_inst_dmem_n15373), .A2(MEM_stage_inst_dmem_n15372), .ZN(MEM_stage_inst_dmem_n11600) );
NAND2_X1 MEM_stage_inst_dmem_U12640 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n15383), .ZN(MEM_stage_inst_dmem_n15372) );
NAND2_X1 MEM_stage_inst_dmem_U12639 ( .A1(MEM_stage_inst_dmem_ram_1301), .A2(MEM_stage_inst_dmem_n15382), .ZN(MEM_stage_inst_dmem_n15373) );
NAND2_X1 MEM_stage_inst_dmem_U12638 ( .A1(MEM_stage_inst_dmem_n15371), .A2(MEM_stage_inst_dmem_n15370), .ZN(MEM_stage_inst_dmem_n11601) );
NAND2_X1 MEM_stage_inst_dmem_U12637 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n15383), .ZN(MEM_stage_inst_dmem_n15370) );
NAND2_X1 MEM_stage_inst_dmem_U12636 ( .A1(MEM_stage_inst_dmem_ram_1302), .A2(MEM_stage_inst_dmem_n15382), .ZN(MEM_stage_inst_dmem_n15371) );
NAND2_X1 MEM_stage_inst_dmem_U12635 ( .A1(MEM_stage_inst_dmem_n15369), .A2(MEM_stage_inst_dmem_n15368), .ZN(MEM_stage_inst_dmem_n11602) );
NAND2_X1 MEM_stage_inst_dmem_U12634 ( .A1(MEM_stage_inst_dmem_n18875), .A2(MEM_stage_inst_dmem_n15383), .ZN(MEM_stage_inst_dmem_n15368) );
NAND2_X1 MEM_stage_inst_dmem_U12633 ( .A1(MEM_stage_inst_dmem_ram_1303), .A2(MEM_stage_inst_dmem_n15382), .ZN(MEM_stage_inst_dmem_n15369) );
NAND2_X1 MEM_stage_inst_dmem_U12632 ( .A1(MEM_stage_inst_dmem_n15367), .A2(MEM_stage_inst_dmem_n15366), .ZN(MEM_stage_inst_dmem_n11603) );
NAND2_X1 MEM_stage_inst_dmem_U12631 ( .A1(MEM_stage_inst_dmem_n111), .A2(MEM_stage_inst_dmem_n15383), .ZN(MEM_stage_inst_dmem_n15366) );
NAND2_X1 MEM_stage_inst_dmem_U12630 ( .A1(MEM_stage_inst_dmem_ram_1304), .A2(MEM_stage_inst_dmem_n15382), .ZN(MEM_stage_inst_dmem_n15367) );
NAND2_X1 MEM_stage_inst_dmem_U12629 ( .A1(MEM_stage_inst_dmem_n15365), .A2(MEM_stage_inst_dmem_n15364), .ZN(MEM_stage_inst_dmem_n11604) );
NAND2_X1 MEM_stage_inst_dmem_U12628 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n15383), .ZN(MEM_stage_inst_dmem_n15364) );
NAND2_X1 MEM_stage_inst_dmem_U12627 ( .A1(MEM_stage_inst_dmem_ram_1305), .A2(MEM_stage_inst_dmem_n15382), .ZN(MEM_stage_inst_dmem_n15365) );
NAND2_X1 MEM_stage_inst_dmem_U12626 ( .A1(MEM_stage_inst_dmem_n15363), .A2(MEM_stage_inst_dmem_n15362), .ZN(MEM_stage_inst_dmem_n11605) );
NAND2_X1 MEM_stage_inst_dmem_U12625 ( .A1(MEM_stage_inst_dmem_n18867), .A2(MEM_stage_inst_dmem_n15383), .ZN(MEM_stage_inst_dmem_n15362) );
NAND2_X1 MEM_stage_inst_dmem_U12624 ( .A1(MEM_stage_inst_dmem_ram_1306), .A2(MEM_stage_inst_dmem_n15382), .ZN(MEM_stage_inst_dmem_n15363) );
NAND2_X1 MEM_stage_inst_dmem_U12623 ( .A1(MEM_stage_inst_dmem_n15361), .A2(MEM_stage_inst_dmem_n15360), .ZN(MEM_stage_inst_dmem_n11606) );
NAND2_X1 MEM_stage_inst_dmem_U12622 ( .A1(MEM_stage_inst_dmem_n18864), .A2(MEM_stage_inst_dmem_n15383), .ZN(MEM_stage_inst_dmem_n15360) );
NAND2_X1 MEM_stage_inst_dmem_U12621 ( .A1(MEM_stage_inst_dmem_ram_1307), .A2(MEM_stage_inst_dmem_n15382), .ZN(MEM_stage_inst_dmem_n15361) );
NAND2_X1 MEM_stage_inst_dmem_U12620 ( .A1(MEM_stage_inst_dmem_n15359), .A2(MEM_stage_inst_dmem_n15358), .ZN(MEM_stage_inst_dmem_n11607) );
NAND2_X1 MEM_stage_inst_dmem_U12619 ( .A1(MEM_stage_inst_dmem_n18861), .A2(MEM_stage_inst_dmem_n15383), .ZN(MEM_stage_inst_dmem_n15358) );
NAND2_X1 MEM_stage_inst_dmem_U12618 ( .A1(MEM_stage_inst_dmem_ram_1308), .A2(MEM_stage_inst_dmem_n15382), .ZN(MEM_stage_inst_dmem_n15359) );
NAND2_X1 MEM_stage_inst_dmem_U12617 ( .A1(MEM_stage_inst_dmem_n15357), .A2(MEM_stage_inst_dmem_n15356), .ZN(MEM_stage_inst_dmem_n11608) );
NAND2_X1 MEM_stage_inst_dmem_U12616 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n15383), .ZN(MEM_stage_inst_dmem_n15356) );
NAND2_X1 MEM_stage_inst_dmem_U12615 ( .A1(MEM_stage_inst_dmem_ram_1309), .A2(MEM_stage_inst_dmem_n15382), .ZN(MEM_stage_inst_dmem_n15357) );
NAND2_X1 MEM_stage_inst_dmem_U12614 ( .A1(MEM_stage_inst_dmem_n15355), .A2(MEM_stage_inst_dmem_n15354), .ZN(MEM_stage_inst_dmem_n11609) );
NAND2_X1 MEM_stage_inst_dmem_U12613 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n15383), .ZN(MEM_stage_inst_dmem_n15354) );
NAND2_X1 MEM_stage_inst_dmem_U12612 ( .A1(MEM_stage_inst_dmem_ram_1310), .A2(MEM_stage_inst_dmem_n15382), .ZN(MEM_stage_inst_dmem_n15355) );
NAND2_X1 MEM_stage_inst_dmem_U12611 ( .A1(MEM_stage_inst_dmem_n15353), .A2(MEM_stage_inst_dmem_n15352), .ZN(MEM_stage_inst_dmem_n11610) );
NAND2_X1 MEM_stage_inst_dmem_U12610 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n15383), .ZN(MEM_stage_inst_dmem_n15352) );
INV_X1 MEM_stage_inst_dmem_U12609 ( .A(MEM_stage_inst_dmem_n15382), .ZN(MEM_stage_inst_dmem_n15383) );
NAND2_X1 MEM_stage_inst_dmem_U12608 ( .A1(MEM_stage_inst_dmem_ram_1311), .A2(MEM_stage_inst_dmem_n15382), .ZN(MEM_stage_inst_dmem_n15353) );
NAND2_X1 MEM_stage_inst_dmem_U12607 ( .A1(MEM_stage_inst_dmem_n21429), .A2(MEM_stage_inst_dmem_n15386), .ZN(MEM_stage_inst_dmem_n15382) );
NAND2_X1 MEM_stage_inst_dmem_U12606 ( .A1(MEM_stage_inst_dmem_n15351), .A2(MEM_stage_inst_dmem_n15350), .ZN(MEM_stage_inst_dmem_n11611) );
NAND2_X1 MEM_stage_inst_dmem_U12605 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n15349), .ZN(MEM_stage_inst_dmem_n15350) );
NAND2_X1 MEM_stage_inst_dmem_U12604 ( .A1(MEM_stage_inst_dmem_ram_1312), .A2(MEM_stage_inst_dmem_n15348), .ZN(MEM_stage_inst_dmem_n15351) );
NAND2_X1 MEM_stage_inst_dmem_U12603 ( .A1(MEM_stage_inst_dmem_n15347), .A2(MEM_stage_inst_dmem_n15346), .ZN(MEM_stage_inst_dmem_n11612) );
NAND2_X1 MEM_stage_inst_dmem_U12602 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n15349), .ZN(MEM_stage_inst_dmem_n15346) );
NAND2_X1 MEM_stage_inst_dmem_U12601 ( .A1(MEM_stage_inst_dmem_ram_1313), .A2(MEM_stage_inst_dmem_n15348), .ZN(MEM_stage_inst_dmem_n15347) );
NAND2_X1 MEM_stage_inst_dmem_U12600 ( .A1(MEM_stage_inst_dmem_n15345), .A2(MEM_stage_inst_dmem_n15344), .ZN(MEM_stage_inst_dmem_n11613) );
NAND2_X1 MEM_stage_inst_dmem_U12599 ( .A1(MEM_stage_inst_dmem_n18887), .A2(MEM_stage_inst_dmem_n15349), .ZN(MEM_stage_inst_dmem_n15344) );
NAND2_X1 MEM_stage_inst_dmem_U12598 ( .A1(MEM_stage_inst_dmem_ram_1314), .A2(MEM_stage_inst_dmem_n15348), .ZN(MEM_stage_inst_dmem_n15345) );
NAND2_X1 MEM_stage_inst_dmem_U12597 ( .A1(MEM_stage_inst_dmem_n15343), .A2(MEM_stage_inst_dmem_n15342), .ZN(MEM_stage_inst_dmem_n11614) );
NAND2_X1 MEM_stage_inst_dmem_U12596 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n15349), .ZN(MEM_stage_inst_dmem_n15342) );
NAND2_X1 MEM_stage_inst_dmem_U12595 ( .A1(MEM_stage_inst_dmem_ram_1315), .A2(MEM_stage_inst_dmem_n15348), .ZN(MEM_stage_inst_dmem_n15343) );
NAND2_X1 MEM_stage_inst_dmem_U12594 ( .A1(MEM_stage_inst_dmem_n15341), .A2(MEM_stage_inst_dmem_n15340), .ZN(MEM_stage_inst_dmem_n11615) );
NAND2_X1 MEM_stage_inst_dmem_U12593 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n15349), .ZN(MEM_stage_inst_dmem_n15340) );
NAND2_X1 MEM_stage_inst_dmem_U12592 ( .A1(MEM_stage_inst_dmem_ram_1316), .A2(MEM_stage_inst_dmem_n15348), .ZN(MEM_stage_inst_dmem_n15341) );
NAND2_X1 MEM_stage_inst_dmem_U12591 ( .A1(MEM_stage_inst_dmem_n15339), .A2(MEM_stage_inst_dmem_n15338), .ZN(MEM_stage_inst_dmem_n11616) );
NAND2_X1 MEM_stage_inst_dmem_U12590 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n15349), .ZN(MEM_stage_inst_dmem_n15338) );
NAND2_X1 MEM_stage_inst_dmem_U12589 ( .A1(MEM_stage_inst_dmem_ram_1317), .A2(MEM_stage_inst_dmem_n15348), .ZN(MEM_stage_inst_dmem_n15339) );
NAND2_X1 MEM_stage_inst_dmem_U12588 ( .A1(MEM_stage_inst_dmem_n15337), .A2(MEM_stage_inst_dmem_n15336), .ZN(MEM_stage_inst_dmem_n11617) );
NAND2_X1 MEM_stage_inst_dmem_U12587 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n15349), .ZN(MEM_stage_inst_dmem_n15336) );
NAND2_X1 MEM_stage_inst_dmem_U12586 ( .A1(MEM_stage_inst_dmem_ram_1318), .A2(MEM_stage_inst_dmem_n15348), .ZN(MEM_stage_inst_dmem_n15337) );
NAND2_X1 MEM_stage_inst_dmem_U12585 ( .A1(MEM_stage_inst_dmem_n15335), .A2(MEM_stage_inst_dmem_n15334), .ZN(MEM_stage_inst_dmem_n11618) );
NAND2_X1 MEM_stage_inst_dmem_U12584 ( .A1(MEM_stage_inst_dmem_n18875), .A2(MEM_stage_inst_dmem_n15349), .ZN(MEM_stage_inst_dmem_n15334) );
NAND2_X1 MEM_stage_inst_dmem_U12583 ( .A1(MEM_stage_inst_dmem_ram_1319), .A2(MEM_stage_inst_dmem_n15348), .ZN(MEM_stage_inst_dmem_n15335) );
NAND2_X1 MEM_stage_inst_dmem_U12582 ( .A1(MEM_stage_inst_dmem_n15333), .A2(MEM_stage_inst_dmem_n15332), .ZN(MEM_stage_inst_dmem_n11619) );
NAND2_X1 MEM_stage_inst_dmem_U12581 ( .A1(MEM_stage_inst_dmem_n111), .A2(MEM_stage_inst_dmem_n15349), .ZN(MEM_stage_inst_dmem_n15332) );
NAND2_X1 MEM_stage_inst_dmem_U12580 ( .A1(MEM_stage_inst_dmem_ram_1320), .A2(MEM_stage_inst_dmem_n15348), .ZN(MEM_stage_inst_dmem_n15333) );
NAND2_X1 MEM_stage_inst_dmem_U12579 ( .A1(MEM_stage_inst_dmem_n15331), .A2(MEM_stage_inst_dmem_n15330), .ZN(MEM_stage_inst_dmem_n11620) );
NAND2_X1 MEM_stage_inst_dmem_U12578 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n15349), .ZN(MEM_stage_inst_dmem_n15330) );
NAND2_X1 MEM_stage_inst_dmem_U12577 ( .A1(MEM_stage_inst_dmem_ram_1321), .A2(MEM_stage_inst_dmem_n15348), .ZN(MEM_stage_inst_dmem_n15331) );
NAND2_X1 MEM_stage_inst_dmem_U12576 ( .A1(MEM_stage_inst_dmem_n15329), .A2(MEM_stage_inst_dmem_n15328), .ZN(MEM_stage_inst_dmem_n11621) );
NAND2_X1 MEM_stage_inst_dmem_U12575 ( .A1(MEM_stage_inst_dmem_n18867), .A2(MEM_stage_inst_dmem_n15349), .ZN(MEM_stage_inst_dmem_n15328) );
NAND2_X1 MEM_stage_inst_dmem_U12574 ( .A1(MEM_stage_inst_dmem_ram_1322), .A2(MEM_stage_inst_dmem_n15348), .ZN(MEM_stage_inst_dmem_n15329) );
NAND2_X1 MEM_stage_inst_dmem_U12573 ( .A1(MEM_stage_inst_dmem_n15327), .A2(MEM_stage_inst_dmem_n15326), .ZN(MEM_stage_inst_dmem_n11622) );
NAND2_X1 MEM_stage_inst_dmem_U12572 ( .A1(MEM_stage_inst_dmem_n18864), .A2(MEM_stage_inst_dmem_n15349), .ZN(MEM_stage_inst_dmem_n15326) );
NAND2_X1 MEM_stage_inst_dmem_U12571 ( .A1(MEM_stage_inst_dmem_ram_1323), .A2(MEM_stage_inst_dmem_n15348), .ZN(MEM_stage_inst_dmem_n15327) );
NAND2_X1 MEM_stage_inst_dmem_U12570 ( .A1(MEM_stage_inst_dmem_n15325), .A2(MEM_stage_inst_dmem_n15324), .ZN(MEM_stage_inst_dmem_n11623) );
NAND2_X1 MEM_stage_inst_dmem_U12569 ( .A1(MEM_stage_inst_dmem_n18861), .A2(MEM_stage_inst_dmem_n15349), .ZN(MEM_stage_inst_dmem_n15324) );
NAND2_X1 MEM_stage_inst_dmem_U12568 ( .A1(MEM_stage_inst_dmem_ram_1324), .A2(MEM_stage_inst_dmem_n15348), .ZN(MEM_stage_inst_dmem_n15325) );
NAND2_X1 MEM_stage_inst_dmem_U12567 ( .A1(MEM_stage_inst_dmem_n15323), .A2(MEM_stage_inst_dmem_n15322), .ZN(MEM_stage_inst_dmem_n11624) );
NAND2_X1 MEM_stage_inst_dmem_U12566 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n15349), .ZN(MEM_stage_inst_dmem_n15322) );
NAND2_X1 MEM_stage_inst_dmem_U12565 ( .A1(MEM_stage_inst_dmem_ram_1325), .A2(MEM_stage_inst_dmem_n15348), .ZN(MEM_stage_inst_dmem_n15323) );
NAND2_X1 MEM_stage_inst_dmem_U12564 ( .A1(MEM_stage_inst_dmem_n15321), .A2(MEM_stage_inst_dmem_n15320), .ZN(MEM_stage_inst_dmem_n11625) );
NAND2_X1 MEM_stage_inst_dmem_U12563 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n15349), .ZN(MEM_stage_inst_dmem_n15320) );
NAND2_X1 MEM_stage_inst_dmem_U12562 ( .A1(MEM_stage_inst_dmem_ram_1326), .A2(MEM_stage_inst_dmem_n15348), .ZN(MEM_stage_inst_dmem_n15321) );
NAND2_X1 MEM_stage_inst_dmem_U12561 ( .A1(MEM_stage_inst_dmem_n15319), .A2(MEM_stage_inst_dmem_n15318), .ZN(MEM_stage_inst_dmem_n11626) );
NAND2_X1 MEM_stage_inst_dmem_U12560 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n15349), .ZN(MEM_stage_inst_dmem_n15318) );
INV_X1 MEM_stage_inst_dmem_U12559 ( .A(MEM_stage_inst_dmem_n15348), .ZN(MEM_stage_inst_dmem_n15349) );
NAND2_X1 MEM_stage_inst_dmem_U12558 ( .A1(MEM_stage_inst_dmem_ram_1327), .A2(MEM_stage_inst_dmem_n15348), .ZN(MEM_stage_inst_dmem_n15319) );
NAND2_X1 MEM_stage_inst_dmem_U12557 ( .A1(MEM_stage_inst_dmem_n21394), .A2(MEM_stage_inst_dmem_n15386), .ZN(MEM_stage_inst_dmem_n15348) );
NAND2_X1 MEM_stage_inst_dmem_U12556 ( .A1(MEM_stage_inst_dmem_n15317), .A2(MEM_stage_inst_dmem_n15316), .ZN(MEM_stage_inst_dmem_n11627) );
NAND2_X1 MEM_stage_inst_dmem_U12555 ( .A1(EX_pipeline_reg_out_5), .A2(MEM_stage_inst_dmem_n15315), .ZN(MEM_stage_inst_dmem_n15316) );
NAND2_X1 MEM_stage_inst_dmem_U12554 ( .A1(MEM_stage_inst_dmem_ram_1328), .A2(MEM_stage_inst_dmem_n15314), .ZN(MEM_stage_inst_dmem_n15317) );
NAND2_X1 MEM_stage_inst_dmem_U12553 ( .A1(MEM_stage_inst_dmem_n15313), .A2(MEM_stage_inst_dmem_n15312), .ZN(MEM_stage_inst_dmem_n11628) );
NAND2_X1 MEM_stage_inst_dmem_U12552 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n15315), .ZN(MEM_stage_inst_dmem_n15312) );
NAND2_X1 MEM_stage_inst_dmem_U12551 ( .A1(MEM_stage_inst_dmem_ram_1329), .A2(MEM_stage_inst_dmem_n15314), .ZN(MEM_stage_inst_dmem_n15313) );
NAND2_X1 MEM_stage_inst_dmem_U12550 ( .A1(MEM_stage_inst_dmem_n15311), .A2(MEM_stage_inst_dmem_n15310), .ZN(MEM_stage_inst_dmem_n11629) );
NAND2_X1 MEM_stage_inst_dmem_U12549 ( .A1(MEM_stage_inst_dmem_n18887), .A2(MEM_stage_inst_dmem_n15315), .ZN(MEM_stage_inst_dmem_n15310) );
NAND2_X1 MEM_stage_inst_dmem_U12548 ( .A1(MEM_stage_inst_dmem_ram_1330), .A2(MEM_stage_inst_dmem_n15314), .ZN(MEM_stage_inst_dmem_n15311) );
NAND2_X1 MEM_stage_inst_dmem_U12547 ( .A1(MEM_stage_inst_dmem_n15309), .A2(MEM_stage_inst_dmem_n15308), .ZN(MEM_stage_inst_dmem_n11630) );
NAND2_X1 MEM_stage_inst_dmem_U12546 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n15315), .ZN(MEM_stage_inst_dmem_n15308) );
NAND2_X1 MEM_stage_inst_dmem_U12545 ( .A1(MEM_stage_inst_dmem_ram_1331), .A2(MEM_stage_inst_dmem_n15314), .ZN(MEM_stage_inst_dmem_n15309) );
NAND2_X1 MEM_stage_inst_dmem_U12544 ( .A1(MEM_stage_inst_dmem_n15307), .A2(MEM_stage_inst_dmem_n15306), .ZN(MEM_stage_inst_dmem_n11631) );
NAND2_X1 MEM_stage_inst_dmem_U12543 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n15315), .ZN(MEM_stage_inst_dmem_n15306) );
NAND2_X1 MEM_stage_inst_dmem_U12542 ( .A1(MEM_stage_inst_dmem_ram_1332), .A2(MEM_stage_inst_dmem_n15314), .ZN(MEM_stage_inst_dmem_n15307) );
NAND2_X1 MEM_stage_inst_dmem_U12541 ( .A1(MEM_stage_inst_dmem_n15305), .A2(MEM_stage_inst_dmem_n15304), .ZN(MEM_stage_inst_dmem_n11632) );
NAND2_X1 MEM_stage_inst_dmem_U12540 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n15315), .ZN(MEM_stage_inst_dmem_n15304) );
NAND2_X1 MEM_stage_inst_dmem_U12539 ( .A1(MEM_stage_inst_dmem_ram_1333), .A2(MEM_stage_inst_dmem_n15314), .ZN(MEM_stage_inst_dmem_n15305) );
NAND2_X1 MEM_stage_inst_dmem_U12538 ( .A1(MEM_stage_inst_dmem_n15303), .A2(MEM_stage_inst_dmem_n15302), .ZN(MEM_stage_inst_dmem_n11633) );
NAND2_X1 MEM_stage_inst_dmem_U12537 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n15315), .ZN(MEM_stage_inst_dmem_n15302) );
NAND2_X1 MEM_stage_inst_dmem_U12536 ( .A1(MEM_stage_inst_dmem_ram_1334), .A2(MEM_stage_inst_dmem_n15314), .ZN(MEM_stage_inst_dmem_n15303) );
NAND2_X1 MEM_stage_inst_dmem_U12535 ( .A1(MEM_stage_inst_dmem_n15301), .A2(MEM_stage_inst_dmem_n15300), .ZN(MEM_stage_inst_dmem_n11634) );
NAND2_X1 MEM_stage_inst_dmem_U12534 ( .A1(MEM_stage_inst_dmem_n18875), .A2(MEM_stage_inst_dmem_n15315), .ZN(MEM_stage_inst_dmem_n15300) );
NAND2_X1 MEM_stage_inst_dmem_U12533 ( .A1(MEM_stage_inst_dmem_ram_1335), .A2(MEM_stage_inst_dmem_n15314), .ZN(MEM_stage_inst_dmem_n15301) );
NAND2_X1 MEM_stage_inst_dmem_U12532 ( .A1(MEM_stage_inst_dmem_n15299), .A2(MEM_stage_inst_dmem_n15298), .ZN(MEM_stage_inst_dmem_n11635) );
NAND2_X1 MEM_stage_inst_dmem_U12531 ( .A1(MEM_stage_inst_dmem_n111), .A2(MEM_stage_inst_dmem_n15315), .ZN(MEM_stage_inst_dmem_n15298) );
NAND2_X1 MEM_stage_inst_dmem_U12530 ( .A1(MEM_stage_inst_dmem_ram_1336), .A2(MEM_stage_inst_dmem_n15314), .ZN(MEM_stage_inst_dmem_n15299) );
NAND2_X1 MEM_stage_inst_dmem_U12529 ( .A1(MEM_stage_inst_dmem_n15297), .A2(MEM_stage_inst_dmem_n15296), .ZN(MEM_stage_inst_dmem_n11636) );
NAND2_X1 MEM_stage_inst_dmem_U12528 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n15315), .ZN(MEM_stage_inst_dmem_n15296) );
NAND2_X1 MEM_stage_inst_dmem_U12527 ( .A1(MEM_stage_inst_dmem_ram_1337), .A2(MEM_stage_inst_dmem_n15314), .ZN(MEM_stage_inst_dmem_n15297) );
NAND2_X1 MEM_stage_inst_dmem_U12526 ( .A1(MEM_stage_inst_dmem_n15295), .A2(MEM_stage_inst_dmem_n15294), .ZN(MEM_stage_inst_dmem_n11637) );
NAND2_X1 MEM_stage_inst_dmem_U12525 ( .A1(MEM_stage_inst_dmem_n18867), .A2(MEM_stage_inst_dmem_n15315), .ZN(MEM_stage_inst_dmem_n15294) );
NAND2_X1 MEM_stage_inst_dmem_U12524 ( .A1(MEM_stage_inst_dmem_ram_1338), .A2(MEM_stage_inst_dmem_n15314), .ZN(MEM_stage_inst_dmem_n15295) );
NAND2_X1 MEM_stage_inst_dmem_U12523 ( .A1(MEM_stage_inst_dmem_n15293), .A2(MEM_stage_inst_dmem_n15292), .ZN(MEM_stage_inst_dmem_n11638) );
NAND2_X1 MEM_stage_inst_dmem_U12522 ( .A1(MEM_stage_inst_dmem_n18864), .A2(MEM_stage_inst_dmem_n15315), .ZN(MEM_stage_inst_dmem_n15292) );
NAND2_X1 MEM_stage_inst_dmem_U12521 ( .A1(MEM_stage_inst_dmem_ram_1339), .A2(MEM_stage_inst_dmem_n15314), .ZN(MEM_stage_inst_dmem_n15293) );
NAND2_X1 MEM_stage_inst_dmem_U12520 ( .A1(MEM_stage_inst_dmem_n15291), .A2(MEM_stage_inst_dmem_n15290), .ZN(MEM_stage_inst_dmem_n11639) );
NAND2_X1 MEM_stage_inst_dmem_U12519 ( .A1(MEM_stage_inst_dmem_n18861), .A2(MEM_stage_inst_dmem_n15315), .ZN(MEM_stage_inst_dmem_n15290) );
NAND2_X1 MEM_stage_inst_dmem_U12518 ( .A1(MEM_stage_inst_dmem_ram_1340), .A2(MEM_stage_inst_dmem_n15314), .ZN(MEM_stage_inst_dmem_n15291) );
NAND2_X1 MEM_stage_inst_dmem_U12517 ( .A1(MEM_stage_inst_dmem_n15289), .A2(MEM_stage_inst_dmem_n15288), .ZN(MEM_stage_inst_dmem_n11640) );
NAND2_X1 MEM_stage_inst_dmem_U12516 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n15315), .ZN(MEM_stage_inst_dmem_n15288) );
NAND2_X1 MEM_stage_inst_dmem_U12515 ( .A1(MEM_stage_inst_dmem_ram_1341), .A2(MEM_stage_inst_dmem_n15314), .ZN(MEM_stage_inst_dmem_n15289) );
NAND2_X1 MEM_stage_inst_dmem_U12514 ( .A1(MEM_stage_inst_dmem_n15287), .A2(MEM_stage_inst_dmem_n15286), .ZN(MEM_stage_inst_dmem_n11641) );
NAND2_X1 MEM_stage_inst_dmem_U12513 ( .A1(EX_pipeline_reg_out_19), .A2(MEM_stage_inst_dmem_n15315), .ZN(MEM_stage_inst_dmem_n15286) );
NAND2_X1 MEM_stage_inst_dmem_U12512 ( .A1(MEM_stage_inst_dmem_ram_1342), .A2(MEM_stage_inst_dmem_n15314), .ZN(MEM_stage_inst_dmem_n15287) );
NAND2_X1 MEM_stage_inst_dmem_U12511 ( .A1(MEM_stage_inst_dmem_n15285), .A2(MEM_stage_inst_dmem_n15284), .ZN(MEM_stage_inst_dmem_n11642) );
NAND2_X1 MEM_stage_inst_dmem_U12510 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n15315), .ZN(MEM_stage_inst_dmem_n15284) );
INV_X1 MEM_stage_inst_dmem_U12509 ( .A(MEM_stage_inst_dmem_n15314), .ZN(MEM_stage_inst_dmem_n15315) );
NAND2_X1 MEM_stage_inst_dmem_U12508 ( .A1(MEM_stage_inst_dmem_ram_1343), .A2(MEM_stage_inst_dmem_n15314), .ZN(MEM_stage_inst_dmem_n15285) );
NAND2_X1 MEM_stage_inst_dmem_U12507 ( .A1(MEM_stage_inst_dmem_n21359), .A2(MEM_stage_inst_dmem_n15386), .ZN(MEM_stage_inst_dmem_n15314) );
NAND2_X1 MEM_stage_inst_dmem_U12506 ( .A1(MEM_stage_inst_dmem_n15283), .A2(MEM_stage_inst_dmem_n15282), .ZN(MEM_stage_inst_dmem_n11643) );
NAND2_X1 MEM_stage_inst_dmem_U12505 ( .A1(MEM_stage_inst_dmem_n20551), .A2(MEM_stage_inst_dmem_n15281), .ZN(MEM_stage_inst_dmem_n15282) );
NAND2_X1 MEM_stage_inst_dmem_U12504 ( .A1(MEM_stage_inst_dmem_ram_1344), .A2(MEM_stage_inst_dmem_n15280), .ZN(MEM_stage_inst_dmem_n15283) );
NAND2_X1 MEM_stage_inst_dmem_U12503 ( .A1(MEM_stage_inst_dmem_n15279), .A2(MEM_stage_inst_dmem_n15278), .ZN(MEM_stage_inst_dmem_n11644) );
NAND2_X1 MEM_stage_inst_dmem_U12502 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n15281), .ZN(MEM_stage_inst_dmem_n15278) );
NAND2_X1 MEM_stage_inst_dmem_U12501 ( .A1(MEM_stage_inst_dmem_ram_1345), .A2(MEM_stage_inst_dmem_n15280), .ZN(MEM_stage_inst_dmem_n15279) );
NAND2_X1 MEM_stage_inst_dmem_U12500 ( .A1(MEM_stage_inst_dmem_n15277), .A2(MEM_stage_inst_dmem_n15276), .ZN(MEM_stage_inst_dmem_n11645) );
NAND2_X1 MEM_stage_inst_dmem_U12499 ( .A1(MEM_stage_inst_dmem_n18887), .A2(MEM_stage_inst_dmem_n15281), .ZN(MEM_stage_inst_dmem_n15276) );
NAND2_X1 MEM_stage_inst_dmem_U12498 ( .A1(MEM_stage_inst_dmem_ram_1346), .A2(MEM_stage_inst_dmem_n15280), .ZN(MEM_stage_inst_dmem_n15277) );
NAND2_X1 MEM_stage_inst_dmem_U12497 ( .A1(MEM_stage_inst_dmem_n15275), .A2(MEM_stage_inst_dmem_n15274), .ZN(MEM_stage_inst_dmem_n11646) );
NAND2_X1 MEM_stage_inst_dmem_U12496 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n15281), .ZN(MEM_stage_inst_dmem_n15274) );
NAND2_X1 MEM_stage_inst_dmem_U12495 ( .A1(MEM_stage_inst_dmem_ram_1347), .A2(MEM_stage_inst_dmem_n15280), .ZN(MEM_stage_inst_dmem_n15275) );
NAND2_X1 MEM_stage_inst_dmem_U12494 ( .A1(MEM_stage_inst_dmem_n15273), .A2(MEM_stage_inst_dmem_n15272), .ZN(MEM_stage_inst_dmem_n11647) );
NAND2_X1 MEM_stage_inst_dmem_U12493 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n15281), .ZN(MEM_stage_inst_dmem_n15272) );
NAND2_X1 MEM_stage_inst_dmem_U12492 ( .A1(MEM_stage_inst_dmem_ram_1348), .A2(MEM_stage_inst_dmem_n15280), .ZN(MEM_stage_inst_dmem_n15273) );
NAND2_X1 MEM_stage_inst_dmem_U12491 ( .A1(MEM_stage_inst_dmem_n15271), .A2(MEM_stage_inst_dmem_n15270), .ZN(MEM_stage_inst_dmem_n11648) );
NAND2_X1 MEM_stage_inst_dmem_U12490 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n15281), .ZN(MEM_stage_inst_dmem_n15270) );
NAND2_X1 MEM_stage_inst_dmem_U12489 ( .A1(MEM_stage_inst_dmem_ram_1349), .A2(MEM_stage_inst_dmem_n15280), .ZN(MEM_stage_inst_dmem_n15271) );
NAND2_X1 MEM_stage_inst_dmem_U12488 ( .A1(MEM_stage_inst_dmem_n15269), .A2(MEM_stage_inst_dmem_n15268), .ZN(MEM_stage_inst_dmem_n11649) );
NAND2_X1 MEM_stage_inst_dmem_U12487 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n15281), .ZN(MEM_stage_inst_dmem_n15268) );
NAND2_X1 MEM_stage_inst_dmem_U12486 ( .A1(MEM_stage_inst_dmem_ram_1350), .A2(MEM_stage_inst_dmem_n15280), .ZN(MEM_stage_inst_dmem_n15269) );
NAND2_X1 MEM_stage_inst_dmem_U12485 ( .A1(MEM_stage_inst_dmem_n15267), .A2(MEM_stage_inst_dmem_n15266), .ZN(MEM_stage_inst_dmem_n11650) );
NAND2_X1 MEM_stage_inst_dmem_U12484 ( .A1(MEM_stage_inst_dmem_n18875), .A2(MEM_stage_inst_dmem_n15281), .ZN(MEM_stage_inst_dmem_n15266) );
NAND2_X1 MEM_stage_inst_dmem_U12483 ( .A1(MEM_stage_inst_dmem_ram_1351), .A2(MEM_stage_inst_dmem_n15280), .ZN(MEM_stage_inst_dmem_n15267) );
NAND2_X1 MEM_stage_inst_dmem_U12482 ( .A1(MEM_stage_inst_dmem_n15265), .A2(MEM_stage_inst_dmem_n15264), .ZN(MEM_stage_inst_dmem_n11651) );
NAND2_X1 MEM_stage_inst_dmem_U12481 ( .A1(MEM_stage_inst_dmem_n111), .A2(MEM_stage_inst_dmem_n15281), .ZN(MEM_stage_inst_dmem_n15264) );
NAND2_X1 MEM_stage_inst_dmem_U12480 ( .A1(MEM_stage_inst_dmem_ram_1352), .A2(MEM_stage_inst_dmem_n15280), .ZN(MEM_stage_inst_dmem_n15265) );
NAND2_X1 MEM_stage_inst_dmem_U12479 ( .A1(MEM_stage_inst_dmem_n15263), .A2(MEM_stage_inst_dmem_n15262), .ZN(MEM_stage_inst_dmem_n11652) );
NAND2_X1 MEM_stage_inst_dmem_U12478 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n15281), .ZN(MEM_stage_inst_dmem_n15262) );
NAND2_X1 MEM_stage_inst_dmem_U12477 ( .A1(MEM_stage_inst_dmem_ram_1353), .A2(MEM_stage_inst_dmem_n15280), .ZN(MEM_stage_inst_dmem_n15263) );
NAND2_X1 MEM_stage_inst_dmem_U12476 ( .A1(MEM_stage_inst_dmem_n15261), .A2(MEM_stage_inst_dmem_n15260), .ZN(MEM_stage_inst_dmem_n11653) );
NAND2_X1 MEM_stage_inst_dmem_U12475 ( .A1(MEM_stage_inst_dmem_n18867), .A2(MEM_stage_inst_dmem_n15281), .ZN(MEM_stage_inst_dmem_n15260) );
NAND2_X1 MEM_stage_inst_dmem_U12474 ( .A1(MEM_stage_inst_dmem_ram_1354), .A2(MEM_stage_inst_dmem_n15280), .ZN(MEM_stage_inst_dmem_n15261) );
NAND2_X1 MEM_stage_inst_dmem_U12473 ( .A1(MEM_stage_inst_dmem_n15259), .A2(MEM_stage_inst_dmem_n15258), .ZN(MEM_stage_inst_dmem_n11654) );
NAND2_X1 MEM_stage_inst_dmem_U12472 ( .A1(MEM_stage_inst_dmem_n18864), .A2(MEM_stage_inst_dmem_n15281), .ZN(MEM_stage_inst_dmem_n15258) );
NAND2_X1 MEM_stage_inst_dmem_U12471 ( .A1(MEM_stage_inst_dmem_ram_1355), .A2(MEM_stage_inst_dmem_n15280), .ZN(MEM_stage_inst_dmem_n15259) );
NAND2_X1 MEM_stage_inst_dmem_U12470 ( .A1(MEM_stage_inst_dmem_n15257), .A2(MEM_stage_inst_dmem_n15256), .ZN(MEM_stage_inst_dmem_n11655) );
NAND2_X1 MEM_stage_inst_dmem_U12469 ( .A1(MEM_stage_inst_dmem_n18861), .A2(MEM_stage_inst_dmem_n15281), .ZN(MEM_stage_inst_dmem_n15256) );
NAND2_X1 MEM_stage_inst_dmem_U12468 ( .A1(MEM_stage_inst_dmem_ram_1356), .A2(MEM_stage_inst_dmem_n15280), .ZN(MEM_stage_inst_dmem_n15257) );
NAND2_X1 MEM_stage_inst_dmem_U12467 ( .A1(MEM_stage_inst_dmem_n15255), .A2(MEM_stage_inst_dmem_n15254), .ZN(MEM_stage_inst_dmem_n11656) );
NAND2_X1 MEM_stage_inst_dmem_U12466 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n15281), .ZN(MEM_stage_inst_dmem_n15254) );
NAND2_X1 MEM_stage_inst_dmem_U12465 ( .A1(MEM_stage_inst_dmem_ram_1357), .A2(MEM_stage_inst_dmem_n15280), .ZN(MEM_stage_inst_dmem_n15255) );
NAND2_X1 MEM_stage_inst_dmem_U12464 ( .A1(MEM_stage_inst_dmem_n15253), .A2(MEM_stage_inst_dmem_n15252), .ZN(MEM_stage_inst_dmem_n11657) );
NAND2_X1 MEM_stage_inst_dmem_U12463 ( .A1(MEM_stage_inst_dmem_n20509), .A2(MEM_stage_inst_dmem_n15281), .ZN(MEM_stage_inst_dmem_n15252) );
NAND2_X1 MEM_stage_inst_dmem_U12462 ( .A1(MEM_stage_inst_dmem_ram_1358), .A2(MEM_stage_inst_dmem_n15280), .ZN(MEM_stage_inst_dmem_n15253) );
NAND2_X1 MEM_stage_inst_dmem_U12461 ( .A1(MEM_stage_inst_dmem_n15251), .A2(MEM_stage_inst_dmem_n15250), .ZN(MEM_stage_inst_dmem_n11658) );
NAND2_X1 MEM_stage_inst_dmem_U12460 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n15281), .ZN(MEM_stage_inst_dmem_n15250) );
INV_X1 MEM_stage_inst_dmem_U12459 ( .A(MEM_stage_inst_dmem_n15280), .ZN(MEM_stage_inst_dmem_n15281) );
NAND2_X1 MEM_stage_inst_dmem_U12458 ( .A1(MEM_stage_inst_dmem_ram_1359), .A2(MEM_stage_inst_dmem_n15280), .ZN(MEM_stage_inst_dmem_n15251) );
NAND2_X1 MEM_stage_inst_dmem_U12457 ( .A1(MEM_stage_inst_dmem_n21319), .A2(MEM_stage_inst_dmem_n15386), .ZN(MEM_stage_inst_dmem_n15280) );
NAND2_X1 MEM_stage_inst_dmem_U12456 ( .A1(MEM_stage_inst_dmem_n15249), .A2(MEM_stage_inst_dmem_n15248), .ZN(MEM_stage_inst_dmem_n11659) );
NAND2_X1 MEM_stage_inst_dmem_U12455 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n15247), .ZN(MEM_stage_inst_dmem_n15248) );
NAND2_X1 MEM_stage_inst_dmem_U12454 ( .A1(MEM_stage_inst_dmem_ram_1360), .A2(MEM_stage_inst_dmem_n15246), .ZN(MEM_stage_inst_dmem_n15249) );
NAND2_X1 MEM_stage_inst_dmem_U12453 ( .A1(MEM_stage_inst_dmem_n15245), .A2(MEM_stage_inst_dmem_n15244), .ZN(MEM_stage_inst_dmem_n11660) );
NAND2_X1 MEM_stage_inst_dmem_U12452 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n15247), .ZN(MEM_stage_inst_dmem_n15244) );
NAND2_X1 MEM_stage_inst_dmem_U12451 ( .A1(MEM_stage_inst_dmem_ram_1361), .A2(MEM_stage_inst_dmem_n15246), .ZN(MEM_stage_inst_dmem_n15245) );
NAND2_X1 MEM_stage_inst_dmem_U12450 ( .A1(MEM_stage_inst_dmem_n15243), .A2(MEM_stage_inst_dmem_n15242), .ZN(MEM_stage_inst_dmem_n11661) );
NAND2_X1 MEM_stage_inst_dmem_U12449 ( .A1(MEM_stage_inst_dmem_n18887), .A2(MEM_stage_inst_dmem_n15247), .ZN(MEM_stage_inst_dmem_n15242) );
NAND2_X1 MEM_stage_inst_dmem_U12448 ( .A1(MEM_stage_inst_dmem_ram_1362), .A2(MEM_stage_inst_dmem_n15246), .ZN(MEM_stage_inst_dmem_n15243) );
NAND2_X1 MEM_stage_inst_dmem_U12447 ( .A1(MEM_stage_inst_dmem_n15241), .A2(MEM_stage_inst_dmem_n15240), .ZN(MEM_stage_inst_dmem_n11662) );
NAND2_X1 MEM_stage_inst_dmem_U12446 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n15247), .ZN(MEM_stage_inst_dmem_n15240) );
NAND2_X1 MEM_stage_inst_dmem_U12445 ( .A1(MEM_stage_inst_dmem_ram_1363), .A2(MEM_stage_inst_dmem_n15246), .ZN(MEM_stage_inst_dmem_n15241) );
NAND2_X1 MEM_stage_inst_dmem_U12444 ( .A1(MEM_stage_inst_dmem_n15239), .A2(MEM_stage_inst_dmem_n15238), .ZN(MEM_stage_inst_dmem_n11663) );
NAND2_X1 MEM_stage_inst_dmem_U12443 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n15247), .ZN(MEM_stage_inst_dmem_n15238) );
NAND2_X1 MEM_stage_inst_dmem_U12442 ( .A1(MEM_stage_inst_dmem_ram_1364), .A2(MEM_stage_inst_dmem_n15246), .ZN(MEM_stage_inst_dmem_n15239) );
NAND2_X1 MEM_stage_inst_dmem_U12441 ( .A1(MEM_stage_inst_dmem_n15237), .A2(MEM_stage_inst_dmem_n15236), .ZN(MEM_stage_inst_dmem_n11664) );
NAND2_X1 MEM_stage_inst_dmem_U12440 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n15247), .ZN(MEM_stage_inst_dmem_n15236) );
NAND2_X1 MEM_stage_inst_dmem_U12439 ( .A1(MEM_stage_inst_dmem_ram_1365), .A2(MEM_stage_inst_dmem_n15246), .ZN(MEM_stage_inst_dmem_n15237) );
NAND2_X1 MEM_stage_inst_dmem_U12438 ( .A1(MEM_stage_inst_dmem_n15235), .A2(MEM_stage_inst_dmem_n15234), .ZN(MEM_stage_inst_dmem_n11665) );
NAND2_X1 MEM_stage_inst_dmem_U12437 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n15247), .ZN(MEM_stage_inst_dmem_n15234) );
NAND2_X1 MEM_stage_inst_dmem_U12436 ( .A1(MEM_stage_inst_dmem_ram_1366), .A2(MEM_stage_inst_dmem_n15246), .ZN(MEM_stage_inst_dmem_n15235) );
NAND2_X1 MEM_stage_inst_dmem_U12435 ( .A1(MEM_stage_inst_dmem_n15233), .A2(MEM_stage_inst_dmem_n15232), .ZN(MEM_stage_inst_dmem_n11666) );
NAND2_X1 MEM_stage_inst_dmem_U12434 ( .A1(MEM_stage_inst_dmem_n18875), .A2(MEM_stage_inst_dmem_n15247), .ZN(MEM_stage_inst_dmem_n15232) );
NAND2_X1 MEM_stage_inst_dmem_U12433 ( .A1(MEM_stage_inst_dmem_ram_1367), .A2(MEM_stage_inst_dmem_n15246), .ZN(MEM_stage_inst_dmem_n15233) );
NAND2_X1 MEM_stage_inst_dmem_U12432 ( .A1(MEM_stage_inst_dmem_n15231), .A2(MEM_stage_inst_dmem_n15230), .ZN(MEM_stage_inst_dmem_n11667) );
NAND2_X1 MEM_stage_inst_dmem_U12431 ( .A1(MEM_stage_inst_dmem_n111), .A2(MEM_stage_inst_dmem_n15247), .ZN(MEM_stage_inst_dmem_n15230) );
NAND2_X1 MEM_stage_inst_dmem_U12430 ( .A1(MEM_stage_inst_dmem_ram_1368), .A2(MEM_stage_inst_dmem_n15246), .ZN(MEM_stage_inst_dmem_n15231) );
NAND2_X1 MEM_stage_inst_dmem_U12429 ( .A1(MEM_stage_inst_dmem_n15229), .A2(MEM_stage_inst_dmem_n15228), .ZN(MEM_stage_inst_dmem_n11668) );
NAND2_X1 MEM_stage_inst_dmem_U12428 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n15247), .ZN(MEM_stage_inst_dmem_n15228) );
NAND2_X1 MEM_stage_inst_dmem_U12427 ( .A1(MEM_stage_inst_dmem_ram_1369), .A2(MEM_stage_inst_dmem_n15246), .ZN(MEM_stage_inst_dmem_n15229) );
NAND2_X1 MEM_stage_inst_dmem_U12426 ( .A1(MEM_stage_inst_dmem_n15227), .A2(MEM_stage_inst_dmem_n15226), .ZN(MEM_stage_inst_dmem_n11669) );
NAND2_X1 MEM_stage_inst_dmem_U12425 ( .A1(MEM_stage_inst_dmem_n18867), .A2(MEM_stage_inst_dmem_n15247), .ZN(MEM_stage_inst_dmem_n15226) );
NAND2_X1 MEM_stage_inst_dmem_U12424 ( .A1(MEM_stage_inst_dmem_ram_1370), .A2(MEM_stage_inst_dmem_n15246), .ZN(MEM_stage_inst_dmem_n15227) );
NAND2_X1 MEM_stage_inst_dmem_U12423 ( .A1(MEM_stage_inst_dmem_n15225), .A2(MEM_stage_inst_dmem_n15224), .ZN(MEM_stage_inst_dmem_n11670) );
NAND2_X1 MEM_stage_inst_dmem_U12422 ( .A1(MEM_stage_inst_dmem_n18864), .A2(MEM_stage_inst_dmem_n15247), .ZN(MEM_stage_inst_dmem_n15224) );
NAND2_X1 MEM_stage_inst_dmem_U12421 ( .A1(MEM_stage_inst_dmem_ram_1371), .A2(MEM_stage_inst_dmem_n15246), .ZN(MEM_stage_inst_dmem_n15225) );
NAND2_X1 MEM_stage_inst_dmem_U12420 ( .A1(MEM_stage_inst_dmem_n15223), .A2(MEM_stage_inst_dmem_n15222), .ZN(MEM_stage_inst_dmem_n11671) );
NAND2_X1 MEM_stage_inst_dmem_U12419 ( .A1(MEM_stage_inst_dmem_n18861), .A2(MEM_stage_inst_dmem_n15247), .ZN(MEM_stage_inst_dmem_n15222) );
NAND2_X1 MEM_stage_inst_dmem_U12418 ( .A1(MEM_stage_inst_dmem_ram_1372), .A2(MEM_stage_inst_dmem_n15246), .ZN(MEM_stage_inst_dmem_n15223) );
NAND2_X1 MEM_stage_inst_dmem_U12417 ( .A1(MEM_stage_inst_dmem_n15221), .A2(MEM_stage_inst_dmem_n15220), .ZN(MEM_stage_inst_dmem_n11672) );
NAND2_X1 MEM_stage_inst_dmem_U12416 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n15247), .ZN(MEM_stage_inst_dmem_n15220) );
NAND2_X1 MEM_stage_inst_dmem_U12415 ( .A1(MEM_stage_inst_dmem_ram_1373), .A2(MEM_stage_inst_dmem_n15246), .ZN(MEM_stage_inst_dmem_n15221) );
NAND2_X1 MEM_stage_inst_dmem_U12414 ( .A1(MEM_stage_inst_dmem_n15219), .A2(MEM_stage_inst_dmem_n15218), .ZN(MEM_stage_inst_dmem_n11673) );
NAND2_X1 MEM_stage_inst_dmem_U12413 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n15247), .ZN(MEM_stage_inst_dmem_n15218) );
NAND2_X1 MEM_stage_inst_dmem_U12412 ( .A1(MEM_stage_inst_dmem_ram_1374), .A2(MEM_stage_inst_dmem_n15246), .ZN(MEM_stage_inst_dmem_n15219) );
NAND2_X1 MEM_stage_inst_dmem_U12411 ( .A1(MEM_stage_inst_dmem_n15217), .A2(MEM_stage_inst_dmem_n15216), .ZN(MEM_stage_inst_dmem_n11674) );
NAND2_X1 MEM_stage_inst_dmem_U12410 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n15247), .ZN(MEM_stage_inst_dmem_n15216) );
INV_X1 MEM_stage_inst_dmem_U12409 ( .A(MEM_stage_inst_dmem_n15246), .ZN(MEM_stage_inst_dmem_n15247) );
NAND2_X1 MEM_stage_inst_dmem_U12408 ( .A1(MEM_stage_inst_dmem_ram_1375), .A2(MEM_stage_inst_dmem_n15246), .ZN(MEM_stage_inst_dmem_n15217) );
NAND2_X1 MEM_stage_inst_dmem_U12407 ( .A1(MEM_stage_inst_dmem_n21284), .A2(MEM_stage_inst_dmem_n15386), .ZN(MEM_stage_inst_dmem_n15246) );
NAND2_X1 MEM_stage_inst_dmem_U12406 ( .A1(MEM_stage_inst_dmem_n15215), .A2(MEM_stage_inst_dmem_n15214), .ZN(MEM_stage_inst_dmem_n11675) );
NAND2_X1 MEM_stage_inst_dmem_U12405 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n15213), .ZN(MEM_stage_inst_dmem_n15214) );
NAND2_X1 MEM_stage_inst_dmem_U12404 ( .A1(MEM_stage_inst_dmem_ram_1376), .A2(MEM_stage_inst_dmem_n15212), .ZN(MEM_stage_inst_dmem_n15215) );
NAND2_X1 MEM_stage_inst_dmem_U12403 ( .A1(MEM_stage_inst_dmem_n15211), .A2(MEM_stage_inst_dmem_n15210), .ZN(MEM_stage_inst_dmem_n11676) );
NAND2_X1 MEM_stage_inst_dmem_U12402 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n15213), .ZN(MEM_stage_inst_dmem_n15210) );
NAND2_X1 MEM_stage_inst_dmem_U12401 ( .A1(MEM_stage_inst_dmem_ram_1377), .A2(MEM_stage_inst_dmem_n15212), .ZN(MEM_stage_inst_dmem_n15211) );
NAND2_X1 MEM_stage_inst_dmem_U12400 ( .A1(MEM_stage_inst_dmem_n15209), .A2(MEM_stage_inst_dmem_n15208), .ZN(MEM_stage_inst_dmem_n11677) );
NAND2_X1 MEM_stage_inst_dmem_U12399 ( .A1(MEM_stage_inst_dmem_n18887), .A2(MEM_stage_inst_dmem_n15213), .ZN(MEM_stage_inst_dmem_n15208) );
NAND2_X1 MEM_stage_inst_dmem_U12398 ( .A1(MEM_stage_inst_dmem_ram_1378), .A2(MEM_stage_inst_dmem_n15212), .ZN(MEM_stage_inst_dmem_n15209) );
NAND2_X1 MEM_stage_inst_dmem_U12397 ( .A1(MEM_stage_inst_dmem_n15207), .A2(MEM_stage_inst_dmem_n15206), .ZN(MEM_stage_inst_dmem_n11678) );
NAND2_X1 MEM_stage_inst_dmem_U12396 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n15213), .ZN(MEM_stage_inst_dmem_n15206) );
NAND2_X1 MEM_stage_inst_dmem_U12395 ( .A1(MEM_stage_inst_dmem_ram_1379), .A2(MEM_stage_inst_dmem_n15212), .ZN(MEM_stage_inst_dmem_n15207) );
NAND2_X1 MEM_stage_inst_dmem_U12394 ( .A1(MEM_stage_inst_dmem_n15205), .A2(MEM_stage_inst_dmem_n15204), .ZN(MEM_stage_inst_dmem_n11679) );
NAND2_X1 MEM_stage_inst_dmem_U12393 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n15213), .ZN(MEM_stage_inst_dmem_n15204) );
NAND2_X1 MEM_stage_inst_dmem_U12392 ( .A1(MEM_stage_inst_dmem_ram_1380), .A2(MEM_stage_inst_dmem_n15212), .ZN(MEM_stage_inst_dmem_n15205) );
NAND2_X1 MEM_stage_inst_dmem_U12391 ( .A1(MEM_stage_inst_dmem_n15203), .A2(MEM_stage_inst_dmem_n15202), .ZN(MEM_stage_inst_dmem_n11680) );
NAND2_X1 MEM_stage_inst_dmem_U12390 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n15213), .ZN(MEM_stage_inst_dmem_n15202) );
NAND2_X1 MEM_stage_inst_dmem_U12389 ( .A1(MEM_stage_inst_dmem_ram_1381), .A2(MEM_stage_inst_dmem_n15212), .ZN(MEM_stage_inst_dmem_n15203) );
NAND2_X1 MEM_stage_inst_dmem_U12388 ( .A1(MEM_stage_inst_dmem_n15201), .A2(MEM_stage_inst_dmem_n15200), .ZN(MEM_stage_inst_dmem_n11681) );
NAND2_X1 MEM_stage_inst_dmem_U12387 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n15213), .ZN(MEM_stage_inst_dmem_n15200) );
NAND2_X1 MEM_stage_inst_dmem_U12386 ( .A1(MEM_stage_inst_dmem_ram_1382), .A2(MEM_stage_inst_dmem_n15212), .ZN(MEM_stage_inst_dmem_n15201) );
NAND2_X1 MEM_stage_inst_dmem_U12385 ( .A1(MEM_stage_inst_dmem_n15199), .A2(MEM_stage_inst_dmem_n15198), .ZN(MEM_stage_inst_dmem_n11682) );
NAND2_X1 MEM_stage_inst_dmem_U12384 ( .A1(MEM_stage_inst_dmem_n18875), .A2(MEM_stage_inst_dmem_n15213), .ZN(MEM_stage_inst_dmem_n15198) );
NAND2_X1 MEM_stage_inst_dmem_U12383 ( .A1(MEM_stage_inst_dmem_ram_1383), .A2(MEM_stage_inst_dmem_n15212), .ZN(MEM_stage_inst_dmem_n15199) );
NAND2_X1 MEM_stage_inst_dmem_U12382 ( .A1(MEM_stage_inst_dmem_n15197), .A2(MEM_stage_inst_dmem_n15196), .ZN(MEM_stage_inst_dmem_n11683) );
NAND2_X1 MEM_stage_inst_dmem_U12381 ( .A1(MEM_stage_inst_dmem_n111), .A2(MEM_stage_inst_dmem_n15213), .ZN(MEM_stage_inst_dmem_n15196) );
NAND2_X1 MEM_stage_inst_dmem_U12380 ( .A1(MEM_stage_inst_dmem_ram_1384), .A2(MEM_stage_inst_dmem_n15212), .ZN(MEM_stage_inst_dmem_n15197) );
NAND2_X1 MEM_stage_inst_dmem_U12379 ( .A1(MEM_stage_inst_dmem_n15195), .A2(MEM_stage_inst_dmem_n15194), .ZN(MEM_stage_inst_dmem_n11684) );
NAND2_X1 MEM_stage_inst_dmem_U12378 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n15213), .ZN(MEM_stage_inst_dmem_n15194) );
NAND2_X1 MEM_stage_inst_dmem_U12377 ( .A1(MEM_stage_inst_dmem_ram_1385), .A2(MEM_stage_inst_dmem_n15212), .ZN(MEM_stage_inst_dmem_n15195) );
NAND2_X1 MEM_stage_inst_dmem_U12376 ( .A1(MEM_stage_inst_dmem_n15193), .A2(MEM_stage_inst_dmem_n15192), .ZN(MEM_stage_inst_dmem_n11685) );
NAND2_X1 MEM_stage_inst_dmem_U12375 ( .A1(MEM_stage_inst_dmem_n18867), .A2(MEM_stage_inst_dmem_n15213), .ZN(MEM_stage_inst_dmem_n15192) );
NAND2_X1 MEM_stage_inst_dmem_U12374 ( .A1(MEM_stage_inst_dmem_ram_1386), .A2(MEM_stage_inst_dmem_n15212), .ZN(MEM_stage_inst_dmem_n15193) );
NAND2_X1 MEM_stage_inst_dmem_U12373 ( .A1(MEM_stage_inst_dmem_n15191), .A2(MEM_stage_inst_dmem_n15190), .ZN(MEM_stage_inst_dmem_n11686) );
NAND2_X1 MEM_stage_inst_dmem_U12372 ( .A1(MEM_stage_inst_dmem_n18864), .A2(MEM_stage_inst_dmem_n15213), .ZN(MEM_stage_inst_dmem_n15190) );
NAND2_X1 MEM_stage_inst_dmem_U12371 ( .A1(MEM_stage_inst_dmem_ram_1387), .A2(MEM_stage_inst_dmem_n15212), .ZN(MEM_stage_inst_dmem_n15191) );
NAND2_X1 MEM_stage_inst_dmem_U12370 ( .A1(MEM_stage_inst_dmem_n15189), .A2(MEM_stage_inst_dmem_n15188), .ZN(MEM_stage_inst_dmem_n11687) );
NAND2_X1 MEM_stage_inst_dmem_U12369 ( .A1(MEM_stage_inst_dmem_n18861), .A2(MEM_stage_inst_dmem_n15213), .ZN(MEM_stage_inst_dmem_n15188) );
NAND2_X1 MEM_stage_inst_dmem_U12368 ( .A1(MEM_stage_inst_dmem_ram_1388), .A2(MEM_stage_inst_dmem_n15212), .ZN(MEM_stage_inst_dmem_n15189) );
NAND2_X1 MEM_stage_inst_dmem_U12367 ( .A1(MEM_stage_inst_dmem_n15187), .A2(MEM_stage_inst_dmem_n15186), .ZN(MEM_stage_inst_dmem_n11688) );
NAND2_X1 MEM_stage_inst_dmem_U12366 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n15213), .ZN(MEM_stage_inst_dmem_n15186) );
NAND2_X1 MEM_stage_inst_dmem_U12365 ( .A1(MEM_stage_inst_dmem_ram_1389), .A2(MEM_stage_inst_dmem_n15212), .ZN(MEM_stage_inst_dmem_n15187) );
NAND2_X1 MEM_stage_inst_dmem_U12364 ( .A1(MEM_stage_inst_dmem_n15185), .A2(MEM_stage_inst_dmem_n15184), .ZN(MEM_stage_inst_dmem_n11689) );
NAND2_X1 MEM_stage_inst_dmem_U12363 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n15213), .ZN(MEM_stage_inst_dmem_n15184) );
NAND2_X1 MEM_stage_inst_dmem_U12362 ( .A1(MEM_stage_inst_dmem_ram_1390), .A2(MEM_stage_inst_dmem_n15212), .ZN(MEM_stage_inst_dmem_n15185) );
NAND2_X1 MEM_stage_inst_dmem_U12361 ( .A1(MEM_stage_inst_dmem_n15183), .A2(MEM_stage_inst_dmem_n15182), .ZN(MEM_stage_inst_dmem_n11690) );
NAND2_X1 MEM_stage_inst_dmem_U12360 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n15213), .ZN(MEM_stage_inst_dmem_n15182) );
INV_X1 MEM_stage_inst_dmem_U12359 ( .A(MEM_stage_inst_dmem_n15212), .ZN(MEM_stage_inst_dmem_n15213) );
NAND2_X1 MEM_stage_inst_dmem_U12358 ( .A1(MEM_stage_inst_dmem_ram_1391), .A2(MEM_stage_inst_dmem_n15212), .ZN(MEM_stage_inst_dmem_n15183) );
NAND2_X1 MEM_stage_inst_dmem_U12357 ( .A1(MEM_stage_inst_dmem_n21249), .A2(MEM_stage_inst_dmem_n15386), .ZN(MEM_stage_inst_dmem_n15212) );
NAND2_X1 MEM_stage_inst_dmem_U12356 ( .A1(MEM_stage_inst_dmem_n15181), .A2(MEM_stage_inst_dmem_n15180), .ZN(MEM_stage_inst_dmem_n11691) );
NAND2_X1 MEM_stage_inst_dmem_U12355 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n15179), .ZN(MEM_stage_inst_dmem_n15180) );
NAND2_X1 MEM_stage_inst_dmem_U12354 ( .A1(MEM_stage_inst_dmem_ram_1392), .A2(MEM_stage_inst_dmem_n15178), .ZN(MEM_stage_inst_dmem_n15181) );
NAND2_X1 MEM_stage_inst_dmem_U12353 ( .A1(MEM_stage_inst_dmem_n15177), .A2(MEM_stage_inst_dmem_n15176), .ZN(MEM_stage_inst_dmem_n11692) );
NAND2_X1 MEM_stage_inst_dmem_U12352 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n15179), .ZN(MEM_stage_inst_dmem_n15176) );
NAND2_X1 MEM_stage_inst_dmem_U12351 ( .A1(MEM_stage_inst_dmem_ram_1393), .A2(MEM_stage_inst_dmem_n15178), .ZN(MEM_stage_inst_dmem_n15177) );
NAND2_X1 MEM_stage_inst_dmem_U12350 ( .A1(MEM_stage_inst_dmem_n15175), .A2(MEM_stage_inst_dmem_n15174), .ZN(MEM_stage_inst_dmem_n11693) );
NAND2_X1 MEM_stage_inst_dmem_U12349 ( .A1(MEM_stage_inst_dmem_n18887), .A2(MEM_stage_inst_dmem_n15179), .ZN(MEM_stage_inst_dmem_n15174) );
BUF_X1 MEM_stage_inst_dmem_U12348 ( .A(MEM_stage_inst_dmem_n113), .Z(MEM_stage_inst_dmem_n18887) );
NAND2_X1 MEM_stage_inst_dmem_U12347 ( .A1(MEM_stage_inst_dmem_ram_1394), .A2(MEM_stage_inst_dmem_n15178), .ZN(MEM_stage_inst_dmem_n15175) );
NAND2_X1 MEM_stage_inst_dmem_U12346 ( .A1(MEM_stage_inst_dmem_n15173), .A2(MEM_stage_inst_dmem_n15172), .ZN(MEM_stage_inst_dmem_n11694) );
NAND2_X1 MEM_stage_inst_dmem_U12345 ( .A1(MEM_stage_inst_dmem_n21506), .A2(MEM_stage_inst_dmem_n15179), .ZN(MEM_stage_inst_dmem_n15172) );
NAND2_X1 MEM_stage_inst_dmem_U12344 ( .A1(MEM_stage_inst_dmem_ram_1395), .A2(MEM_stage_inst_dmem_n15178), .ZN(MEM_stage_inst_dmem_n15173) );
NAND2_X1 MEM_stage_inst_dmem_U12343 ( .A1(MEM_stage_inst_dmem_n15171), .A2(MEM_stage_inst_dmem_n15170), .ZN(MEM_stage_inst_dmem_n11695) );
NAND2_X1 MEM_stage_inst_dmem_U12342 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n15179), .ZN(MEM_stage_inst_dmem_n15170) );
NAND2_X1 MEM_stage_inst_dmem_U12341 ( .A1(MEM_stage_inst_dmem_ram_1396), .A2(MEM_stage_inst_dmem_n15178), .ZN(MEM_stage_inst_dmem_n15171) );
NAND2_X1 MEM_stage_inst_dmem_U12340 ( .A1(MEM_stage_inst_dmem_n15169), .A2(MEM_stage_inst_dmem_n15168), .ZN(MEM_stage_inst_dmem_n11696) );
NAND2_X1 MEM_stage_inst_dmem_U12339 ( .A1(MEM_stage_inst_dmem_n21508), .A2(MEM_stage_inst_dmem_n15179), .ZN(MEM_stage_inst_dmem_n15168) );
NAND2_X1 MEM_stage_inst_dmem_U12338 ( .A1(MEM_stage_inst_dmem_ram_1397), .A2(MEM_stage_inst_dmem_n15178), .ZN(MEM_stage_inst_dmem_n15169) );
NAND2_X1 MEM_stage_inst_dmem_U12337 ( .A1(MEM_stage_inst_dmem_n15167), .A2(MEM_stage_inst_dmem_n15166), .ZN(MEM_stage_inst_dmem_n11697) );
NAND2_X1 MEM_stage_inst_dmem_U12336 ( .A1(MEM_stage_inst_dmem_n18878), .A2(MEM_stage_inst_dmem_n15179), .ZN(MEM_stage_inst_dmem_n15166) );
BUF_X2 MEM_stage_inst_dmem_U12335 ( .A(MEM_stage_inst_dmem_n20533), .Z(MEM_stage_inst_dmem_n18878) );
NAND2_X1 MEM_stage_inst_dmem_U12334 ( .A1(MEM_stage_inst_dmem_ram_1398), .A2(MEM_stage_inst_dmem_n15178), .ZN(MEM_stage_inst_dmem_n15167) );
NAND2_X1 MEM_stage_inst_dmem_U12333 ( .A1(MEM_stage_inst_dmem_n15165), .A2(MEM_stage_inst_dmem_n15164), .ZN(MEM_stage_inst_dmem_n11698) );
NAND2_X1 MEM_stage_inst_dmem_U12332 ( .A1(MEM_stage_inst_dmem_n18875), .A2(MEM_stage_inst_dmem_n15179), .ZN(MEM_stage_inst_dmem_n15164) );
BUF_X1 MEM_stage_inst_dmem_U12331 ( .A(MEM_stage_inst_dmem_n18), .Z(MEM_stage_inst_dmem_n18875) );
NAND2_X1 MEM_stage_inst_dmem_U12330 ( .A1(MEM_stage_inst_dmem_ram_1399), .A2(MEM_stage_inst_dmem_n15178), .ZN(MEM_stage_inst_dmem_n15165) );
NAND2_X1 MEM_stage_inst_dmem_U12329 ( .A1(MEM_stage_inst_dmem_n15163), .A2(MEM_stage_inst_dmem_n15162), .ZN(MEM_stage_inst_dmem_n11699) );
NAND2_X1 MEM_stage_inst_dmem_U12328 ( .A1(MEM_stage_inst_dmem_n20527), .A2(MEM_stage_inst_dmem_n15179), .ZN(MEM_stage_inst_dmem_n15162) );
NAND2_X1 MEM_stage_inst_dmem_U12326 ( .A1(MEM_stage_inst_dmem_ram_1400), .A2(MEM_stage_inst_dmem_n15178), .ZN(MEM_stage_inst_dmem_n15163) );
NAND2_X1 MEM_stage_inst_dmem_U12325 ( .A1(MEM_stage_inst_dmem_n15161), .A2(MEM_stage_inst_dmem_n15160), .ZN(MEM_stage_inst_dmem_n11700) );
NAND2_X1 MEM_stage_inst_dmem_U12324 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n15179), .ZN(MEM_stage_inst_dmem_n15160) );
BUF_X1 MEM_stage_inst_dmem_U12323 ( .A(MEM_stage_inst_dmem_n20524), .Z(MEM_stage_inst_dmem_n19251) );
NAND2_X1 MEM_stage_inst_dmem_U12322 ( .A1(MEM_stage_inst_dmem_ram_1401), .A2(MEM_stage_inst_dmem_n15178), .ZN(MEM_stage_inst_dmem_n15161) );
NAND2_X1 MEM_stage_inst_dmem_U12321 ( .A1(MEM_stage_inst_dmem_n15159), .A2(MEM_stage_inst_dmem_n15158), .ZN(MEM_stage_inst_dmem_n11701) );
NAND2_X1 MEM_stage_inst_dmem_U12320 ( .A1(MEM_stage_inst_dmem_n18867), .A2(MEM_stage_inst_dmem_n15179), .ZN(MEM_stage_inst_dmem_n15158) );
BUF_X1 MEM_stage_inst_dmem_U12319 ( .A(MEM_stage_inst_dmem_n102), .Z(MEM_stage_inst_dmem_n18867) );
NAND2_X1 MEM_stage_inst_dmem_U12318 ( .A1(MEM_stage_inst_dmem_ram_1402), .A2(MEM_stage_inst_dmem_n15178), .ZN(MEM_stage_inst_dmem_n15159) );
NAND2_X1 MEM_stage_inst_dmem_U12317 ( .A1(MEM_stage_inst_dmem_n15157), .A2(MEM_stage_inst_dmem_n15156), .ZN(MEM_stage_inst_dmem_n11702) );
NAND2_X1 MEM_stage_inst_dmem_U12316 ( .A1(MEM_stage_inst_dmem_n18864), .A2(MEM_stage_inst_dmem_n15179), .ZN(MEM_stage_inst_dmem_n15156) );
NAND2_X1 MEM_stage_inst_dmem_U12315 ( .A1(MEM_stage_inst_dmem_ram_1403), .A2(MEM_stage_inst_dmem_n15178), .ZN(MEM_stage_inst_dmem_n15157) );
NAND2_X1 MEM_stage_inst_dmem_U12314 ( .A1(MEM_stage_inst_dmem_n15155), .A2(MEM_stage_inst_dmem_n15154), .ZN(MEM_stage_inst_dmem_n11703) );
NAND2_X1 MEM_stage_inst_dmem_U12313 ( .A1(MEM_stage_inst_dmem_n18861), .A2(MEM_stage_inst_dmem_n15179), .ZN(MEM_stage_inst_dmem_n15154) );
NAND2_X1 MEM_stage_inst_dmem_U12312 ( .A1(MEM_stage_inst_dmem_ram_1404), .A2(MEM_stage_inst_dmem_n15178), .ZN(MEM_stage_inst_dmem_n15155) );
NAND2_X1 MEM_stage_inst_dmem_U12311 ( .A1(MEM_stage_inst_dmem_n15153), .A2(MEM_stage_inst_dmem_n15152), .ZN(MEM_stage_inst_dmem_n11704) );
NAND2_X1 MEM_stage_inst_dmem_U12310 ( .A1(MEM_stage_inst_dmem_n15116), .A2(MEM_stage_inst_dmem_n15179), .ZN(MEM_stage_inst_dmem_n15152) );
NAND2_X1 MEM_stage_inst_dmem_U12309 ( .A1(MEM_stage_inst_dmem_ram_1405), .A2(MEM_stage_inst_dmem_n15178), .ZN(MEM_stage_inst_dmem_n15153) );
NAND2_X1 MEM_stage_inst_dmem_U12308 ( .A1(MEM_stage_inst_dmem_n15151), .A2(MEM_stage_inst_dmem_n15150), .ZN(MEM_stage_inst_dmem_n11705) );
NAND2_X1 MEM_stage_inst_dmem_U12307 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n15179), .ZN(MEM_stage_inst_dmem_n15150) );
NAND2_X1 MEM_stage_inst_dmem_U12306 ( .A1(MEM_stage_inst_dmem_ram_1406), .A2(MEM_stage_inst_dmem_n15178), .ZN(MEM_stage_inst_dmem_n15151) );
NAND2_X1 MEM_stage_inst_dmem_U12305 ( .A1(MEM_stage_inst_dmem_n15149), .A2(MEM_stage_inst_dmem_n15148), .ZN(MEM_stage_inst_dmem_n11706) );
NAND2_X1 MEM_stage_inst_dmem_U12304 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n15179), .ZN(MEM_stage_inst_dmem_n15148) );
INV_X1 MEM_stage_inst_dmem_U12303 ( .A(MEM_stage_inst_dmem_n15178), .ZN(MEM_stage_inst_dmem_n15179) );
NAND2_X1 MEM_stage_inst_dmem_U12302 ( .A1(MEM_stage_inst_dmem_ram_1407), .A2(MEM_stage_inst_dmem_n15178), .ZN(MEM_stage_inst_dmem_n15149) );
NAND2_X1 MEM_stage_inst_dmem_U12301 ( .A1(MEM_stage_inst_dmem_n21214), .A2(MEM_stage_inst_dmem_n15386), .ZN(MEM_stage_inst_dmem_n15178) );
NAND2_X1 MEM_stage_inst_dmem_U12300 ( .A1(MEM_stage_inst_dmem_n15147), .A2(MEM_stage_inst_dmem_n15146), .ZN(MEM_stage_inst_dmem_n11707) );
NAND2_X1 MEM_stage_inst_dmem_U12299 ( .A1(MEM_stage_inst_dmem_n15145), .A2(MEM_stage_inst_dmem_n15144), .ZN(MEM_stage_inst_dmem_n15146) );
NAND2_X1 MEM_stage_inst_dmem_U12298 ( .A1(MEM_stage_inst_dmem_ram_1408), .A2(MEM_stage_inst_dmem_n15143), .ZN(MEM_stage_inst_dmem_n15147) );
NAND2_X1 MEM_stage_inst_dmem_U12297 ( .A1(MEM_stage_inst_dmem_n15142), .A2(MEM_stage_inst_dmem_n15141), .ZN(MEM_stage_inst_dmem_n11708) );
NAND2_X1 MEM_stage_inst_dmem_U12296 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n15144), .ZN(MEM_stage_inst_dmem_n15141) );
NAND2_X1 MEM_stage_inst_dmem_U12295 ( .A1(MEM_stage_inst_dmem_ram_1409), .A2(MEM_stage_inst_dmem_n15143), .ZN(MEM_stage_inst_dmem_n15142) );
NAND2_X1 MEM_stage_inst_dmem_U12294 ( .A1(MEM_stage_inst_dmem_n15140), .A2(MEM_stage_inst_dmem_n15139), .ZN(MEM_stage_inst_dmem_n11709) );
NAND2_X1 MEM_stage_inst_dmem_U12293 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n15144), .ZN(MEM_stage_inst_dmem_n15139) );
NAND2_X1 MEM_stage_inst_dmem_U12292 ( .A1(MEM_stage_inst_dmem_ram_1410), .A2(MEM_stage_inst_dmem_n15143), .ZN(MEM_stage_inst_dmem_n15140) );
NAND2_X1 MEM_stage_inst_dmem_U12291 ( .A1(MEM_stage_inst_dmem_n15138), .A2(MEM_stage_inst_dmem_n15137), .ZN(MEM_stage_inst_dmem_n11710) );
NAND2_X1 MEM_stage_inst_dmem_U12290 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n15144), .ZN(MEM_stage_inst_dmem_n15137) );
NAND2_X1 MEM_stage_inst_dmem_U12289 ( .A1(MEM_stage_inst_dmem_ram_1411), .A2(MEM_stage_inst_dmem_n15143), .ZN(MEM_stage_inst_dmem_n15138) );
NAND2_X1 MEM_stage_inst_dmem_U12288 ( .A1(MEM_stage_inst_dmem_n15136), .A2(MEM_stage_inst_dmem_n15135), .ZN(MEM_stage_inst_dmem_n11711) );
NAND2_X1 MEM_stage_inst_dmem_U12287 ( .A1(MEM_stage_inst_dmem_n16368), .A2(MEM_stage_inst_dmem_n15144), .ZN(MEM_stage_inst_dmem_n15135) );
NAND2_X1 MEM_stage_inst_dmem_U12286 ( .A1(MEM_stage_inst_dmem_ram_1412), .A2(MEM_stage_inst_dmem_n15143), .ZN(MEM_stage_inst_dmem_n15136) );
NAND2_X1 MEM_stage_inst_dmem_U12285 ( .A1(MEM_stage_inst_dmem_n15134), .A2(MEM_stage_inst_dmem_n15133), .ZN(MEM_stage_inst_dmem_n11712) );
NAND2_X1 MEM_stage_inst_dmem_U12284 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n15144), .ZN(MEM_stage_inst_dmem_n15133) );
NAND2_X1 MEM_stage_inst_dmem_U12283 ( .A1(MEM_stage_inst_dmem_ram_1413), .A2(MEM_stage_inst_dmem_n15143), .ZN(MEM_stage_inst_dmem_n15134) );
NAND2_X1 MEM_stage_inst_dmem_U12282 ( .A1(MEM_stage_inst_dmem_n15132), .A2(MEM_stage_inst_dmem_n15131), .ZN(MEM_stage_inst_dmem_n11713) );
NAND2_X1 MEM_stage_inst_dmem_U12281 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n15144), .ZN(MEM_stage_inst_dmem_n15131) );
NAND2_X1 MEM_stage_inst_dmem_U12280 ( .A1(MEM_stage_inst_dmem_ram_1414), .A2(MEM_stage_inst_dmem_n15143), .ZN(MEM_stage_inst_dmem_n15132) );
NAND2_X1 MEM_stage_inst_dmem_U12279 ( .A1(MEM_stage_inst_dmem_n15130), .A2(MEM_stage_inst_dmem_n15129), .ZN(MEM_stage_inst_dmem_n11714) );
NAND2_X1 MEM_stage_inst_dmem_U12278 ( .A1(MEM_stage_inst_dmem_n16361), .A2(MEM_stage_inst_dmem_n15144), .ZN(MEM_stage_inst_dmem_n15129) );
NAND2_X1 MEM_stage_inst_dmem_U12277 ( .A1(MEM_stage_inst_dmem_ram_1415), .A2(MEM_stage_inst_dmem_n15143), .ZN(MEM_stage_inst_dmem_n15130) );
NAND2_X1 MEM_stage_inst_dmem_U12276 ( .A1(MEM_stage_inst_dmem_n15128), .A2(MEM_stage_inst_dmem_n15127), .ZN(MEM_stage_inst_dmem_n11715) );
NAND2_X1 MEM_stage_inst_dmem_U12275 ( .A1(MEM_stage_inst_dmem_n13883), .A2(MEM_stage_inst_dmem_n15144), .ZN(MEM_stage_inst_dmem_n15127) );
NAND2_X1 MEM_stage_inst_dmem_U12274 ( .A1(MEM_stage_inst_dmem_ram_1416), .A2(MEM_stage_inst_dmem_n15143), .ZN(MEM_stage_inst_dmem_n15128) );
NAND2_X1 MEM_stage_inst_dmem_U12273 ( .A1(MEM_stage_inst_dmem_n15126), .A2(MEM_stage_inst_dmem_n15125), .ZN(MEM_stage_inst_dmem_n11716) );
NAND2_X1 MEM_stage_inst_dmem_U12272 ( .A1(MEM_stage_inst_dmem_n19251), .A2(MEM_stage_inst_dmem_n15144), .ZN(MEM_stage_inst_dmem_n15125) );
NAND2_X1 MEM_stage_inst_dmem_U12271 ( .A1(MEM_stage_inst_dmem_ram_1417), .A2(MEM_stage_inst_dmem_n15143), .ZN(MEM_stage_inst_dmem_n15126) );
NAND2_X1 MEM_stage_inst_dmem_U12270 ( .A1(MEM_stage_inst_dmem_n15124), .A2(MEM_stage_inst_dmem_n15123), .ZN(MEM_stage_inst_dmem_n11717) );
NAND2_X1 MEM_stage_inst_dmem_U12269 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n15144), .ZN(MEM_stage_inst_dmem_n15123) );
NAND2_X1 MEM_stage_inst_dmem_U12268 ( .A1(MEM_stage_inst_dmem_ram_1418), .A2(MEM_stage_inst_dmem_n15143), .ZN(MEM_stage_inst_dmem_n15124) );
NAND2_X1 MEM_stage_inst_dmem_U12267 ( .A1(MEM_stage_inst_dmem_n15122), .A2(MEM_stage_inst_dmem_n15121), .ZN(MEM_stage_inst_dmem_n11718) );
NAND2_X1 MEM_stage_inst_dmem_U12266 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n15144), .ZN(MEM_stage_inst_dmem_n15121) );
NAND2_X1 MEM_stage_inst_dmem_U12265 ( .A1(MEM_stage_inst_dmem_ram_1419), .A2(MEM_stage_inst_dmem_n15143), .ZN(MEM_stage_inst_dmem_n15122) );
NAND2_X1 MEM_stage_inst_dmem_U12264 ( .A1(MEM_stage_inst_dmem_n15120), .A2(MEM_stage_inst_dmem_n15119), .ZN(MEM_stage_inst_dmem_n11719) );
NAND2_X1 MEM_stage_inst_dmem_U12263 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n15144), .ZN(MEM_stage_inst_dmem_n15119) );
NAND2_X1 MEM_stage_inst_dmem_U12262 ( .A1(MEM_stage_inst_dmem_ram_1420), .A2(MEM_stage_inst_dmem_n15143), .ZN(MEM_stage_inst_dmem_n15120) );
NAND2_X1 MEM_stage_inst_dmem_U12261 ( .A1(MEM_stage_inst_dmem_n15118), .A2(MEM_stage_inst_dmem_n15117), .ZN(MEM_stage_inst_dmem_n11720) );
NAND2_X1 MEM_stage_inst_dmem_U12260 ( .A1(MEM_stage_inst_dmem_n15116), .A2(MEM_stage_inst_dmem_n15144), .ZN(MEM_stage_inst_dmem_n15117) );
NAND2_X1 MEM_stage_inst_dmem_U12259 ( .A1(MEM_stage_inst_dmem_ram_1421), .A2(MEM_stage_inst_dmem_n15143), .ZN(MEM_stage_inst_dmem_n15118) );
NAND2_X1 MEM_stage_inst_dmem_U12258 ( .A1(MEM_stage_inst_dmem_n15115), .A2(MEM_stage_inst_dmem_n15114), .ZN(MEM_stage_inst_dmem_n11721) );
NAND2_X1 MEM_stage_inst_dmem_U12257 ( .A1(MEM_stage_inst_dmem_n15113), .A2(MEM_stage_inst_dmem_n15144), .ZN(MEM_stage_inst_dmem_n15114) );
NAND2_X1 MEM_stage_inst_dmem_U12256 ( .A1(MEM_stage_inst_dmem_ram_1422), .A2(MEM_stage_inst_dmem_n15143), .ZN(MEM_stage_inst_dmem_n15115) );
NAND2_X1 MEM_stage_inst_dmem_U12255 ( .A1(MEM_stage_inst_dmem_n15112), .A2(MEM_stage_inst_dmem_n15111), .ZN(MEM_stage_inst_dmem_n11722) );
NAND2_X1 MEM_stage_inst_dmem_U12254 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n15144), .ZN(MEM_stage_inst_dmem_n15111) );
INV_X1 MEM_stage_inst_dmem_U12253 ( .A(MEM_stage_inst_dmem_n15143), .ZN(MEM_stage_inst_dmem_n15144) );
NAND2_X1 MEM_stage_inst_dmem_U12252 ( .A1(MEM_stage_inst_dmem_ram_1423), .A2(MEM_stage_inst_dmem_n15143), .ZN(MEM_stage_inst_dmem_n15112) );
NAND2_X1 MEM_stage_inst_dmem_U12251 ( .A1(MEM_stage_inst_dmem_n21179), .A2(MEM_stage_inst_dmem_n15386), .ZN(MEM_stage_inst_dmem_n15143) );
NAND2_X1 MEM_stage_inst_dmem_U12250 ( .A1(MEM_stage_inst_dmem_n15109), .A2(MEM_stage_inst_dmem_n15108), .ZN(MEM_stage_inst_dmem_n11723) );
NAND2_X1 MEM_stage_inst_dmem_U12249 ( .A1(MEM_stage_inst_dmem_n15145), .A2(MEM_stage_inst_dmem_n15107), .ZN(MEM_stage_inst_dmem_n15108) );
NAND2_X1 MEM_stage_inst_dmem_U12248 ( .A1(MEM_stage_inst_dmem_ram_1424), .A2(MEM_stage_inst_dmem_n15106), .ZN(MEM_stage_inst_dmem_n15109) );
NAND2_X1 MEM_stage_inst_dmem_U12247 ( .A1(MEM_stage_inst_dmem_n15105), .A2(MEM_stage_inst_dmem_n15104), .ZN(MEM_stage_inst_dmem_n11724) );
NAND2_X1 MEM_stage_inst_dmem_U12246 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n15107), .ZN(MEM_stage_inst_dmem_n15104) );
NAND2_X1 MEM_stage_inst_dmem_U12245 ( .A1(MEM_stage_inst_dmem_ram_1425), .A2(MEM_stage_inst_dmem_n15106), .ZN(MEM_stage_inst_dmem_n15105) );
NAND2_X1 MEM_stage_inst_dmem_U12244 ( .A1(MEM_stage_inst_dmem_n15103), .A2(MEM_stage_inst_dmem_n15102), .ZN(MEM_stage_inst_dmem_n11725) );
NAND2_X1 MEM_stage_inst_dmem_U12243 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n15107), .ZN(MEM_stage_inst_dmem_n15102) );
NAND2_X1 MEM_stage_inst_dmem_U12242 ( .A1(MEM_stage_inst_dmem_ram_1426), .A2(MEM_stage_inst_dmem_n15106), .ZN(MEM_stage_inst_dmem_n15103) );
NAND2_X1 MEM_stage_inst_dmem_U12241 ( .A1(MEM_stage_inst_dmem_n15101), .A2(MEM_stage_inst_dmem_n15100), .ZN(MEM_stage_inst_dmem_n11726) );
NAND2_X1 MEM_stage_inst_dmem_U12240 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n15107), .ZN(MEM_stage_inst_dmem_n15100) );
NAND2_X1 MEM_stage_inst_dmem_U12239 ( .A1(MEM_stage_inst_dmem_ram_1427), .A2(MEM_stage_inst_dmem_n15106), .ZN(MEM_stage_inst_dmem_n15101) );
NAND2_X1 MEM_stage_inst_dmem_U12238 ( .A1(MEM_stage_inst_dmem_n15099), .A2(MEM_stage_inst_dmem_n15098), .ZN(MEM_stage_inst_dmem_n11727) );
NAND2_X1 MEM_stage_inst_dmem_U12237 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n15107), .ZN(MEM_stage_inst_dmem_n15098) );
NAND2_X1 MEM_stage_inst_dmem_U12236 ( .A1(MEM_stage_inst_dmem_ram_1428), .A2(MEM_stage_inst_dmem_n15106), .ZN(MEM_stage_inst_dmem_n15099) );
NAND2_X1 MEM_stage_inst_dmem_U12235 ( .A1(MEM_stage_inst_dmem_n15097), .A2(MEM_stage_inst_dmem_n15096), .ZN(MEM_stage_inst_dmem_n11728) );
NAND2_X1 MEM_stage_inst_dmem_U12234 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n15107), .ZN(MEM_stage_inst_dmem_n15096) );
NAND2_X1 MEM_stage_inst_dmem_U12233 ( .A1(MEM_stage_inst_dmem_ram_1429), .A2(MEM_stage_inst_dmem_n15106), .ZN(MEM_stage_inst_dmem_n15097) );
NAND2_X1 MEM_stage_inst_dmem_U12232 ( .A1(MEM_stage_inst_dmem_n15095), .A2(MEM_stage_inst_dmem_n15094), .ZN(MEM_stage_inst_dmem_n11729) );
NAND2_X1 MEM_stage_inst_dmem_U12231 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n15107), .ZN(MEM_stage_inst_dmem_n15094) );
NAND2_X1 MEM_stage_inst_dmem_U12230 ( .A1(MEM_stage_inst_dmem_ram_1430), .A2(MEM_stage_inst_dmem_n15106), .ZN(MEM_stage_inst_dmem_n15095) );
NAND2_X1 MEM_stage_inst_dmem_U12229 ( .A1(MEM_stage_inst_dmem_n15093), .A2(MEM_stage_inst_dmem_n15092), .ZN(MEM_stage_inst_dmem_n11730) );
NAND2_X1 MEM_stage_inst_dmem_U12228 ( .A1(MEM_stage_inst_dmem_n112), .A2(MEM_stage_inst_dmem_n15107), .ZN(MEM_stage_inst_dmem_n15092) );
NAND2_X1 MEM_stage_inst_dmem_U12227 ( .A1(MEM_stage_inst_dmem_ram_1431), .A2(MEM_stage_inst_dmem_n15106), .ZN(MEM_stage_inst_dmem_n15093) );
NAND2_X1 MEM_stage_inst_dmem_U12226 ( .A1(MEM_stage_inst_dmem_n15091), .A2(MEM_stage_inst_dmem_n15090), .ZN(MEM_stage_inst_dmem_n11731) );
NAND2_X1 MEM_stage_inst_dmem_U12225 ( .A1(MEM_stage_inst_dmem_n13051), .A2(MEM_stage_inst_dmem_n15107), .ZN(MEM_stage_inst_dmem_n15090) );
NAND2_X1 MEM_stage_inst_dmem_U12224 ( .A1(MEM_stage_inst_dmem_ram_1432), .A2(MEM_stage_inst_dmem_n15106), .ZN(MEM_stage_inst_dmem_n15091) );
NAND2_X1 MEM_stage_inst_dmem_U12223 ( .A1(MEM_stage_inst_dmem_n15089), .A2(MEM_stage_inst_dmem_n15088), .ZN(MEM_stage_inst_dmem_n11732) );
NAND2_X1 MEM_stage_inst_dmem_U12222 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n15107), .ZN(MEM_stage_inst_dmem_n15088) );
NAND2_X1 MEM_stage_inst_dmem_U12221 ( .A1(MEM_stage_inst_dmem_ram_1433), .A2(MEM_stage_inst_dmem_n15106), .ZN(MEM_stage_inst_dmem_n15089) );
NAND2_X1 MEM_stage_inst_dmem_U12220 ( .A1(MEM_stage_inst_dmem_n15087), .A2(MEM_stage_inst_dmem_n15086), .ZN(MEM_stage_inst_dmem_n11733) );
NAND2_X1 MEM_stage_inst_dmem_U12219 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n15107), .ZN(MEM_stage_inst_dmem_n15086) );
NAND2_X1 MEM_stage_inst_dmem_U12218 ( .A1(MEM_stage_inst_dmem_ram_1434), .A2(MEM_stage_inst_dmem_n15106), .ZN(MEM_stage_inst_dmem_n15087) );
NAND2_X1 MEM_stage_inst_dmem_U12217 ( .A1(MEM_stage_inst_dmem_n15085), .A2(MEM_stage_inst_dmem_n15084), .ZN(MEM_stage_inst_dmem_n11734) );
NAND2_X1 MEM_stage_inst_dmem_U12216 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n15107), .ZN(MEM_stage_inst_dmem_n15084) );
NAND2_X1 MEM_stage_inst_dmem_U12215 ( .A1(MEM_stage_inst_dmem_ram_1435), .A2(MEM_stage_inst_dmem_n15106), .ZN(MEM_stage_inst_dmem_n15085) );
NAND2_X1 MEM_stage_inst_dmem_U12214 ( .A1(MEM_stage_inst_dmem_n15083), .A2(MEM_stage_inst_dmem_n15082), .ZN(MEM_stage_inst_dmem_n11735) );
NAND2_X1 MEM_stage_inst_dmem_U12213 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n15107), .ZN(MEM_stage_inst_dmem_n15082) );
NAND2_X1 MEM_stage_inst_dmem_U12212 ( .A1(MEM_stage_inst_dmem_ram_1436), .A2(MEM_stage_inst_dmem_n15106), .ZN(MEM_stage_inst_dmem_n15083) );
NAND2_X1 MEM_stage_inst_dmem_U12211 ( .A1(MEM_stage_inst_dmem_n15081), .A2(MEM_stage_inst_dmem_n15080), .ZN(MEM_stage_inst_dmem_n11736) );
NAND2_X1 MEM_stage_inst_dmem_U12210 ( .A1(MEM_stage_inst_dmem_n15116), .A2(MEM_stage_inst_dmem_n15107), .ZN(MEM_stage_inst_dmem_n15080) );
NAND2_X1 MEM_stage_inst_dmem_U12209 ( .A1(MEM_stage_inst_dmem_ram_1437), .A2(MEM_stage_inst_dmem_n15106), .ZN(MEM_stage_inst_dmem_n15081) );
NAND2_X1 MEM_stage_inst_dmem_U12208 ( .A1(MEM_stage_inst_dmem_n15079), .A2(MEM_stage_inst_dmem_n15078), .ZN(MEM_stage_inst_dmem_n11737) );
NAND2_X1 MEM_stage_inst_dmem_U12207 ( .A1(MEM_stage_inst_dmem_n15113), .A2(MEM_stage_inst_dmem_n15107), .ZN(MEM_stage_inst_dmem_n15078) );
NAND2_X1 MEM_stage_inst_dmem_U12206 ( .A1(MEM_stage_inst_dmem_ram_1438), .A2(MEM_stage_inst_dmem_n15106), .ZN(MEM_stage_inst_dmem_n15079) );
NAND2_X1 MEM_stage_inst_dmem_U12205 ( .A1(MEM_stage_inst_dmem_n15077), .A2(MEM_stage_inst_dmem_n15076), .ZN(MEM_stage_inst_dmem_n11738) );
NAND2_X1 MEM_stage_inst_dmem_U12204 ( .A1(MEM_stage_inst_dmem_n16343), .A2(MEM_stage_inst_dmem_n15107), .ZN(MEM_stage_inst_dmem_n15076) );
INV_X1 MEM_stage_inst_dmem_U12203 ( .A(MEM_stage_inst_dmem_n15106), .ZN(MEM_stage_inst_dmem_n15107) );
NAND2_X1 MEM_stage_inst_dmem_U12202 ( .A1(MEM_stage_inst_dmem_ram_1439), .A2(MEM_stage_inst_dmem_n15106), .ZN(MEM_stage_inst_dmem_n15077) );
NAND2_X1 MEM_stage_inst_dmem_U12201 ( .A1(MEM_stage_inst_dmem_n21144), .A2(MEM_stage_inst_dmem_n15386), .ZN(MEM_stage_inst_dmem_n15106) );
NAND2_X1 MEM_stage_inst_dmem_U12200 ( .A1(MEM_stage_inst_dmem_n15075), .A2(MEM_stage_inst_dmem_n15074), .ZN(MEM_stage_inst_dmem_n11739) );
NAND2_X1 MEM_stage_inst_dmem_U12199 ( .A1(MEM_stage_inst_dmem_n15145), .A2(MEM_stage_inst_dmem_n15073), .ZN(MEM_stage_inst_dmem_n15074) );
NAND2_X1 MEM_stage_inst_dmem_U12198 ( .A1(MEM_stage_inst_dmem_ram_1440), .A2(MEM_stage_inst_dmem_n15072), .ZN(MEM_stage_inst_dmem_n15075) );
NAND2_X1 MEM_stage_inst_dmem_U12197 ( .A1(MEM_stage_inst_dmem_n15071), .A2(MEM_stage_inst_dmem_n15070), .ZN(MEM_stage_inst_dmem_n11740) );
NAND2_X1 MEM_stage_inst_dmem_U12196 ( .A1(EX_pipeline_reg_out_6), .A2(MEM_stage_inst_dmem_n15073), .ZN(MEM_stage_inst_dmem_n15070) );
NAND2_X1 MEM_stage_inst_dmem_U12195 ( .A1(MEM_stage_inst_dmem_ram_1441), .A2(MEM_stage_inst_dmem_n15072), .ZN(MEM_stage_inst_dmem_n15071) );
NAND2_X1 MEM_stage_inst_dmem_U12194 ( .A1(MEM_stage_inst_dmem_n15069), .A2(MEM_stage_inst_dmem_n15068), .ZN(MEM_stage_inst_dmem_n11741) );
NAND2_X1 MEM_stage_inst_dmem_U12193 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n15073), .ZN(MEM_stage_inst_dmem_n15068) );
NAND2_X1 MEM_stage_inst_dmem_U12192 ( .A1(MEM_stage_inst_dmem_ram_1442), .A2(MEM_stage_inst_dmem_n15072), .ZN(MEM_stage_inst_dmem_n15069) );
NAND2_X1 MEM_stage_inst_dmem_U12191 ( .A1(MEM_stage_inst_dmem_n15067), .A2(MEM_stage_inst_dmem_n15066), .ZN(MEM_stage_inst_dmem_n11742) );
NAND2_X1 MEM_stage_inst_dmem_U12190 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n15073), .ZN(MEM_stage_inst_dmem_n15066) );
NAND2_X1 MEM_stage_inst_dmem_U12189 ( .A1(MEM_stage_inst_dmem_ram_1443), .A2(MEM_stage_inst_dmem_n15072), .ZN(MEM_stage_inst_dmem_n15067) );
NAND2_X1 MEM_stage_inst_dmem_U12188 ( .A1(MEM_stage_inst_dmem_n15065), .A2(MEM_stage_inst_dmem_n15064), .ZN(MEM_stage_inst_dmem_n11743) );
NAND2_X1 MEM_stage_inst_dmem_U12187 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n15073), .ZN(MEM_stage_inst_dmem_n15064) );
NAND2_X1 MEM_stage_inst_dmem_U12186 ( .A1(MEM_stage_inst_dmem_ram_1444), .A2(MEM_stage_inst_dmem_n15072), .ZN(MEM_stage_inst_dmem_n15065) );
NAND2_X1 MEM_stage_inst_dmem_U12185 ( .A1(MEM_stage_inst_dmem_n15063), .A2(MEM_stage_inst_dmem_n15062), .ZN(MEM_stage_inst_dmem_n11744) );
NAND2_X1 MEM_stage_inst_dmem_U12184 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n15073), .ZN(MEM_stage_inst_dmem_n15062) );
NAND2_X1 MEM_stage_inst_dmem_U12183 ( .A1(MEM_stage_inst_dmem_ram_1445), .A2(MEM_stage_inst_dmem_n15072), .ZN(MEM_stage_inst_dmem_n15063) );
NAND2_X1 MEM_stage_inst_dmem_U12182 ( .A1(MEM_stage_inst_dmem_n15061), .A2(MEM_stage_inst_dmem_n15060), .ZN(MEM_stage_inst_dmem_n11745) );
NAND2_X1 MEM_stage_inst_dmem_U12181 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n15073), .ZN(MEM_stage_inst_dmem_n15060) );
NAND2_X1 MEM_stage_inst_dmem_U12180 ( .A1(MEM_stage_inst_dmem_ram_1446), .A2(MEM_stage_inst_dmem_n15072), .ZN(MEM_stage_inst_dmem_n15061) );
NAND2_X1 MEM_stage_inst_dmem_U12179 ( .A1(MEM_stage_inst_dmem_n15059), .A2(MEM_stage_inst_dmem_n15058), .ZN(MEM_stage_inst_dmem_n11746) );
NAND2_X1 MEM_stage_inst_dmem_U12178 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n15073), .ZN(MEM_stage_inst_dmem_n15058) );
NAND2_X1 MEM_stage_inst_dmem_U12177 ( .A1(MEM_stage_inst_dmem_ram_1447), .A2(MEM_stage_inst_dmem_n15072), .ZN(MEM_stage_inst_dmem_n15059) );
NAND2_X1 MEM_stage_inst_dmem_U12176 ( .A1(MEM_stage_inst_dmem_n15057), .A2(MEM_stage_inst_dmem_n15056), .ZN(MEM_stage_inst_dmem_n11747) );
NAND2_X1 MEM_stage_inst_dmem_U12175 ( .A1(MEM_stage_inst_dmem_n111), .A2(MEM_stage_inst_dmem_n15073), .ZN(MEM_stage_inst_dmem_n15056) );
NAND2_X1 MEM_stage_inst_dmem_U12174 ( .A1(MEM_stage_inst_dmem_ram_1448), .A2(MEM_stage_inst_dmem_n15072), .ZN(MEM_stage_inst_dmem_n15057) );
NAND2_X1 MEM_stage_inst_dmem_U12173 ( .A1(MEM_stage_inst_dmem_n15055), .A2(MEM_stage_inst_dmem_n15054), .ZN(MEM_stage_inst_dmem_n11748) );
NAND2_X1 MEM_stage_inst_dmem_U12172 ( .A1(MEM_stage_inst_dmem_n19251), .A2(MEM_stage_inst_dmem_n15073), .ZN(MEM_stage_inst_dmem_n15054) );
NAND2_X1 MEM_stage_inst_dmem_U12171 ( .A1(MEM_stage_inst_dmem_ram_1449), .A2(MEM_stage_inst_dmem_n15072), .ZN(MEM_stage_inst_dmem_n15055) );
NAND2_X1 MEM_stage_inst_dmem_U12170 ( .A1(MEM_stage_inst_dmem_n15053), .A2(MEM_stage_inst_dmem_n15052), .ZN(MEM_stage_inst_dmem_n11749) );
NAND2_X1 MEM_stage_inst_dmem_U12169 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n15073), .ZN(MEM_stage_inst_dmem_n15052) );
NAND2_X1 MEM_stage_inst_dmem_U12168 ( .A1(MEM_stage_inst_dmem_ram_1450), .A2(MEM_stage_inst_dmem_n15072), .ZN(MEM_stage_inst_dmem_n15053) );
NAND2_X1 MEM_stage_inst_dmem_U12167 ( .A1(MEM_stage_inst_dmem_n15051), .A2(MEM_stage_inst_dmem_n15050), .ZN(MEM_stage_inst_dmem_n11750) );
NAND2_X1 MEM_stage_inst_dmem_U12166 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n15073), .ZN(MEM_stage_inst_dmem_n15050) );
NAND2_X1 MEM_stage_inst_dmem_U12165 ( .A1(MEM_stage_inst_dmem_ram_1451), .A2(MEM_stage_inst_dmem_n15072), .ZN(MEM_stage_inst_dmem_n15051) );
NAND2_X1 MEM_stage_inst_dmem_U12164 ( .A1(MEM_stage_inst_dmem_n15049), .A2(MEM_stage_inst_dmem_n15048), .ZN(MEM_stage_inst_dmem_n11751) );
NAND2_X1 MEM_stage_inst_dmem_U12163 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n15073), .ZN(MEM_stage_inst_dmem_n15048) );
NAND2_X1 MEM_stage_inst_dmem_U12162 ( .A1(MEM_stage_inst_dmem_ram_1452), .A2(MEM_stage_inst_dmem_n15072), .ZN(MEM_stage_inst_dmem_n15049) );
NAND2_X1 MEM_stage_inst_dmem_U12161 ( .A1(MEM_stage_inst_dmem_n15047), .A2(MEM_stage_inst_dmem_n15046), .ZN(MEM_stage_inst_dmem_n11752) );
NAND2_X1 MEM_stage_inst_dmem_U12160 ( .A1(MEM_stage_inst_dmem_n15116), .A2(MEM_stage_inst_dmem_n15073), .ZN(MEM_stage_inst_dmem_n15046) );
NAND2_X1 MEM_stage_inst_dmem_U12159 ( .A1(MEM_stage_inst_dmem_ram_1453), .A2(MEM_stage_inst_dmem_n15072), .ZN(MEM_stage_inst_dmem_n15047) );
NAND2_X1 MEM_stage_inst_dmem_U12158 ( .A1(MEM_stage_inst_dmem_n15045), .A2(MEM_stage_inst_dmem_n15044), .ZN(MEM_stage_inst_dmem_n11753) );
NAND2_X1 MEM_stage_inst_dmem_U12157 ( .A1(MEM_stage_inst_dmem_n15113), .A2(MEM_stage_inst_dmem_n15073), .ZN(MEM_stage_inst_dmem_n15044) );
NAND2_X1 MEM_stage_inst_dmem_U12156 ( .A1(MEM_stage_inst_dmem_ram_1454), .A2(MEM_stage_inst_dmem_n15072), .ZN(MEM_stage_inst_dmem_n15045) );
NAND2_X1 MEM_stage_inst_dmem_U12155 ( .A1(MEM_stage_inst_dmem_n15043), .A2(MEM_stage_inst_dmem_n15042), .ZN(MEM_stage_inst_dmem_n11754) );
NAND2_X1 MEM_stage_inst_dmem_U12154 ( .A1(MEM_stage_inst_dmem_n14693), .A2(MEM_stage_inst_dmem_n15073), .ZN(MEM_stage_inst_dmem_n15042) );
INV_X1 MEM_stage_inst_dmem_U12153 ( .A(MEM_stage_inst_dmem_n15072), .ZN(MEM_stage_inst_dmem_n15073) );
NAND2_X1 MEM_stage_inst_dmem_U12152 ( .A1(MEM_stage_inst_dmem_ram_1455), .A2(MEM_stage_inst_dmem_n15072), .ZN(MEM_stage_inst_dmem_n15043) );
NAND2_X1 MEM_stage_inst_dmem_U12151 ( .A1(MEM_stage_inst_dmem_n21109), .A2(MEM_stage_inst_dmem_n15386), .ZN(MEM_stage_inst_dmem_n15072) );
NAND2_X1 MEM_stage_inst_dmem_U12150 ( .A1(MEM_stage_inst_dmem_n15041), .A2(MEM_stage_inst_dmem_n15040), .ZN(MEM_stage_inst_dmem_n11755) );
NAND2_X1 MEM_stage_inst_dmem_U12149 ( .A1(MEM_stage_inst_dmem_n15145), .A2(MEM_stage_inst_dmem_n15039), .ZN(MEM_stage_inst_dmem_n15040) );
NAND2_X1 MEM_stage_inst_dmem_U12148 ( .A1(MEM_stage_inst_dmem_ram_1456), .A2(MEM_stage_inst_dmem_n15038), .ZN(MEM_stage_inst_dmem_n15041) );
NAND2_X1 MEM_stage_inst_dmem_U12147 ( .A1(MEM_stage_inst_dmem_n15037), .A2(MEM_stage_inst_dmem_n15036), .ZN(MEM_stage_inst_dmem_n11756) );
NAND2_X1 MEM_stage_inst_dmem_U12146 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n15039), .ZN(MEM_stage_inst_dmem_n15036) );
NAND2_X1 MEM_stage_inst_dmem_U12145 ( .A1(MEM_stage_inst_dmem_ram_1457), .A2(MEM_stage_inst_dmem_n15038), .ZN(MEM_stage_inst_dmem_n15037) );
NAND2_X1 MEM_stage_inst_dmem_U12144 ( .A1(MEM_stage_inst_dmem_n15035), .A2(MEM_stage_inst_dmem_n15034), .ZN(MEM_stage_inst_dmem_n11757) );
NAND2_X1 MEM_stage_inst_dmem_U12143 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n15039), .ZN(MEM_stage_inst_dmem_n15034) );
NAND2_X1 MEM_stage_inst_dmem_U12142 ( .A1(MEM_stage_inst_dmem_ram_1458), .A2(MEM_stage_inst_dmem_n15038), .ZN(MEM_stage_inst_dmem_n15035) );
NAND2_X1 MEM_stage_inst_dmem_U12141 ( .A1(MEM_stage_inst_dmem_n15033), .A2(MEM_stage_inst_dmem_n15032), .ZN(MEM_stage_inst_dmem_n11758) );
NAND2_X1 MEM_stage_inst_dmem_U12140 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n15039), .ZN(MEM_stage_inst_dmem_n15032) );
NAND2_X1 MEM_stage_inst_dmem_U12139 ( .A1(MEM_stage_inst_dmem_ram_1459), .A2(MEM_stage_inst_dmem_n15038), .ZN(MEM_stage_inst_dmem_n15033) );
NAND2_X1 MEM_stage_inst_dmem_U12138 ( .A1(MEM_stage_inst_dmem_n15031), .A2(MEM_stage_inst_dmem_n15030), .ZN(MEM_stage_inst_dmem_n11759) );
NAND2_X1 MEM_stage_inst_dmem_U12137 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n15039), .ZN(MEM_stage_inst_dmem_n15030) );
NAND2_X1 MEM_stage_inst_dmem_U12136 ( .A1(MEM_stage_inst_dmem_ram_1460), .A2(MEM_stage_inst_dmem_n15038), .ZN(MEM_stage_inst_dmem_n15031) );
NAND2_X1 MEM_stage_inst_dmem_U12135 ( .A1(MEM_stage_inst_dmem_n15029), .A2(MEM_stage_inst_dmem_n15028), .ZN(MEM_stage_inst_dmem_n11760) );
NAND2_X1 MEM_stage_inst_dmem_U12134 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n15039), .ZN(MEM_stage_inst_dmem_n15028) );
NAND2_X1 MEM_stage_inst_dmem_U12133 ( .A1(MEM_stage_inst_dmem_ram_1461), .A2(MEM_stage_inst_dmem_n15038), .ZN(MEM_stage_inst_dmem_n15029) );
NAND2_X1 MEM_stage_inst_dmem_U12132 ( .A1(MEM_stage_inst_dmem_n15027), .A2(MEM_stage_inst_dmem_n15026), .ZN(MEM_stage_inst_dmem_n11761) );
NAND2_X1 MEM_stage_inst_dmem_U12131 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n15039), .ZN(MEM_stage_inst_dmem_n15026) );
NAND2_X1 MEM_stage_inst_dmem_U12130 ( .A1(MEM_stage_inst_dmem_ram_1462), .A2(MEM_stage_inst_dmem_n15038), .ZN(MEM_stage_inst_dmem_n15027) );
NAND2_X1 MEM_stage_inst_dmem_U12129 ( .A1(MEM_stage_inst_dmem_n15025), .A2(MEM_stage_inst_dmem_n15024), .ZN(MEM_stage_inst_dmem_n11762) );
NAND2_X1 MEM_stage_inst_dmem_U12128 ( .A1(MEM_stage_inst_dmem_n112), .A2(MEM_stage_inst_dmem_n15039), .ZN(MEM_stage_inst_dmem_n15024) );
NAND2_X1 MEM_stage_inst_dmem_U12127 ( .A1(MEM_stage_inst_dmem_ram_1463), .A2(MEM_stage_inst_dmem_n15038), .ZN(MEM_stage_inst_dmem_n15025) );
NAND2_X1 MEM_stage_inst_dmem_U12126 ( .A1(MEM_stage_inst_dmem_n15023), .A2(MEM_stage_inst_dmem_n15022), .ZN(MEM_stage_inst_dmem_n11763) );
NAND2_X1 MEM_stage_inst_dmem_U12125 ( .A1(MEM_stage_inst_dmem_n21335), .A2(MEM_stage_inst_dmem_n15039), .ZN(MEM_stage_inst_dmem_n15022) );
NAND2_X1 MEM_stage_inst_dmem_U12124 ( .A1(MEM_stage_inst_dmem_ram_1464), .A2(MEM_stage_inst_dmem_n15038), .ZN(MEM_stage_inst_dmem_n15023) );
NAND2_X1 MEM_stage_inst_dmem_U12123 ( .A1(MEM_stage_inst_dmem_n15021), .A2(MEM_stage_inst_dmem_n15020), .ZN(MEM_stage_inst_dmem_n11764) );
NAND2_X1 MEM_stage_inst_dmem_U12122 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n15039), .ZN(MEM_stage_inst_dmem_n15020) );
NAND2_X1 MEM_stage_inst_dmem_U12121 ( .A1(MEM_stage_inst_dmem_ram_1465), .A2(MEM_stage_inst_dmem_n15038), .ZN(MEM_stage_inst_dmem_n15021) );
NAND2_X1 MEM_stage_inst_dmem_U12120 ( .A1(MEM_stage_inst_dmem_n15019), .A2(MEM_stage_inst_dmem_n15018), .ZN(MEM_stage_inst_dmem_n11765) );
NAND2_X1 MEM_stage_inst_dmem_U12119 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n15039), .ZN(MEM_stage_inst_dmem_n15018) );
NAND2_X1 MEM_stage_inst_dmem_U12118 ( .A1(MEM_stage_inst_dmem_ram_1466), .A2(MEM_stage_inst_dmem_n15038), .ZN(MEM_stage_inst_dmem_n15019) );
NAND2_X1 MEM_stage_inst_dmem_U12117 ( .A1(MEM_stage_inst_dmem_n15017), .A2(MEM_stage_inst_dmem_n15016), .ZN(MEM_stage_inst_dmem_n11766) );
NAND2_X1 MEM_stage_inst_dmem_U12116 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n15039), .ZN(MEM_stage_inst_dmem_n15016) );
NAND2_X1 MEM_stage_inst_dmem_U12115 ( .A1(MEM_stage_inst_dmem_ram_1467), .A2(MEM_stage_inst_dmem_n15038), .ZN(MEM_stage_inst_dmem_n15017) );
NAND2_X1 MEM_stage_inst_dmem_U12114 ( .A1(MEM_stage_inst_dmem_n15015), .A2(MEM_stage_inst_dmem_n15014), .ZN(MEM_stage_inst_dmem_n11767) );
NAND2_X1 MEM_stage_inst_dmem_U12113 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n15039), .ZN(MEM_stage_inst_dmem_n15014) );
NAND2_X1 MEM_stage_inst_dmem_U12112 ( .A1(MEM_stage_inst_dmem_ram_1468), .A2(MEM_stage_inst_dmem_n15038), .ZN(MEM_stage_inst_dmem_n15015) );
NAND2_X1 MEM_stage_inst_dmem_U12111 ( .A1(MEM_stage_inst_dmem_n15013), .A2(MEM_stage_inst_dmem_n15012), .ZN(MEM_stage_inst_dmem_n11768) );
NAND2_X1 MEM_stage_inst_dmem_U12110 ( .A1(MEM_stage_inst_dmem_n15116), .A2(MEM_stage_inst_dmem_n15039), .ZN(MEM_stage_inst_dmem_n15012) );
NAND2_X1 MEM_stage_inst_dmem_U12109 ( .A1(MEM_stage_inst_dmem_ram_1469), .A2(MEM_stage_inst_dmem_n15038), .ZN(MEM_stage_inst_dmem_n15013) );
NAND2_X1 MEM_stage_inst_dmem_U12108 ( .A1(MEM_stage_inst_dmem_n15011), .A2(MEM_stage_inst_dmem_n15010), .ZN(MEM_stage_inst_dmem_n11769) );
NAND2_X1 MEM_stage_inst_dmem_U12107 ( .A1(MEM_stage_inst_dmem_n15113), .A2(MEM_stage_inst_dmem_n15039), .ZN(MEM_stage_inst_dmem_n15010) );
NAND2_X1 MEM_stage_inst_dmem_U12106 ( .A1(MEM_stage_inst_dmem_ram_1470), .A2(MEM_stage_inst_dmem_n15038), .ZN(MEM_stage_inst_dmem_n15011) );
NAND2_X1 MEM_stage_inst_dmem_U12105 ( .A1(MEM_stage_inst_dmem_n15009), .A2(MEM_stage_inst_dmem_n15008), .ZN(MEM_stage_inst_dmem_n11770) );
NAND2_X1 MEM_stage_inst_dmem_U12104 ( .A1(MEM_stage_inst_dmem_n15110), .A2(MEM_stage_inst_dmem_n15039), .ZN(MEM_stage_inst_dmem_n15008) );
INV_X1 MEM_stage_inst_dmem_U12103 ( .A(MEM_stage_inst_dmem_n15038), .ZN(MEM_stage_inst_dmem_n15039) );
NAND2_X1 MEM_stage_inst_dmem_U12102 ( .A1(MEM_stage_inst_dmem_ram_1471), .A2(MEM_stage_inst_dmem_n15038), .ZN(MEM_stage_inst_dmem_n15009) );
NAND2_X1 MEM_stage_inst_dmem_U12101 ( .A1(MEM_stage_inst_dmem_n21074), .A2(MEM_stage_inst_dmem_n15386), .ZN(MEM_stage_inst_dmem_n15038) );
NAND2_X1 MEM_stage_inst_dmem_U12100 ( .A1(MEM_stage_inst_dmem_n15007), .A2(MEM_stage_inst_dmem_n15006), .ZN(MEM_stage_inst_dmem_n11771) );
NAND2_X1 MEM_stage_inst_dmem_U12099 ( .A1(MEM_stage_inst_dmem_n15145), .A2(MEM_stage_inst_dmem_n15005), .ZN(MEM_stage_inst_dmem_n15006) );
NAND2_X1 MEM_stage_inst_dmem_U12098 ( .A1(MEM_stage_inst_dmem_ram_1472), .A2(MEM_stage_inst_dmem_n15004), .ZN(MEM_stage_inst_dmem_n15007) );
NAND2_X1 MEM_stage_inst_dmem_U12097 ( .A1(MEM_stage_inst_dmem_n15003), .A2(MEM_stage_inst_dmem_n15002), .ZN(MEM_stage_inst_dmem_n11772) );
NAND2_X1 MEM_stage_inst_dmem_U12096 ( .A1(MEM_stage_inst_dmem_n20547), .A2(MEM_stage_inst_dmem_n15005), .ZN(MEM_stage_inst_dmem_n15002) );
NAND2_X1 MEM_stage_inst_dmem_U12095 ( .A1(MEM_stage_inst_dmem_ram_1473), .A2(MEM_stage_inst_dmem_n15004), .ZN(MEM_stage_inst_dmem_n15003) );
NAND2_X1 MEM_stage_inst_dmem_U12094 ( .A1(MEM_stage_inst_dmem_n15001), .A2(MEM_stage_inst_dmem_n15000), .ZN(MEM_stage_inst_dmem_n11773) );
NAND2_X1 MEM_stage_inst_dmem_U12093 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n15005), .ZN(MEM_stage_inst_dmem_n15000) );
NAND2_X1 MEM_stage_inst_dmem_U12092 ( .A1(MEM_stage_inst_dmem_ram_1474), .A2(MEM_stage_inst_dmem_n15004), .ZN(MEM_stage_inst_dmem_n15001) );
NAND2_X1 MEM_stage_inst_dmem_U12091 ( .A1(MEM_stage_inst_dmem_n14999), .A2(MEM_stage_inst_dmem_n14998), .ZN(MEM_stage_inst_dmem_n11774) );
NAND2_X1 MEM_stage_inst_dmem_U12090 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n15005), .ZN(MEM_stage_inst_dmem_n14998) );
NAND2_X1 MEM_stage_inst_dmem_U12089 ( .A1(MEM_stage_inst_dmem_ram_1475), .A2(MEM_stage_inst_dmem_n15004), .ZN(MEM_stage_inst_dmem_n14999) );
NAND2_X1 MEM_stage_inst_dmem_U12088 ( .A1(MEM_stage_inst_dmem_n14997), .A2(MEM_stage_inst_dmem_n14996), .ZN(MEM_stage_inst_dmem_n11775) );
NAND2_X1 MEM_stage_inst_dmem_U12087 ( .A1(MEM_stage_inst_dmem_n16368), .A2(MEM_stage_inst_dmem_n15005), .ZN(MEM_stage_inst_dmem_n14996) );
NAND2_X1 MEM_stage_inst_dmem_U12086 ( .A1(MEM_stage_inst_dmem_ram_1476), .A2(MEM_stage_inst_dmem_n15004), .ZN(MEM_stage_inst_dmem_n14997) );
NAND2_X1 MEM_stage_inst_dmem_U12085 ( .A1(MEM_stage_inst_dmem_n14995), .A2(MEM_stage_inst_dmem_n14994), .ZN(MEM_stage_inst_dmem_n11776) );
NAND2_X1 MEM_stage_inst_dmem_U12084 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n15005), .ZN(MEM_stage_inst_dmem_n14994) );
NAND2_X1 MEM_stage_inst_dmem_U12083 ( .A1(MEM_stage_inst_dmem_ram_1477), .A2(MEM_stage_inst_dmem_n15004), .ZN(MEM_stage_inst_dmem_n14995) );
NAND2_X1 MEM_stage_inst_dmem_U12082 ( .A1(MEM_stage_inst_dmem_n14993), .A2(MEM_stage_inst_dmem_n14992), .ZN(MEM_stage_inst_dmem_n11777) );
NAND2_X1 MEM_stage_inst_dmem_U12081 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n15005), .ZN(MEM_stage_inst_dmem_n14992) );
NAND2_X1 MEM_stage_inst_dmem_U12080 ( .A1(MEM_stage_inst_dmem_ram_1478), .A2(MEM_stage_inst_dmem_n15004), .ZN(MEM_stage_inst_dmem_n14993) );
NAND2_X1 MEM_stage_inst_dmem_U12079 ( .A1(MEM_stage_inst_dmem_n14991), .A2(MEM_stage_inst_dmem_n14990), .ZN(MEM_stage_inst_dmem_n11778) );
NAND2_X1 MEM_stage_inst_dmem_U12078 ( .A1(MEM_stage_inst_dmem_n16361), .A2(MEM_stage_inst_dmem_n15005), .ZN(MEM_stage_inst_dmem_n14990) );
NAND2_X1 MEM_stage_inst_dmem_U12077 ( .A1(MEM_stage_inst_dmem_ram_1479), .A2(MEM_stage_inst_dmem_n15004), .ZN(MEM_stage_inst_dmem_n14991) );
NAND2_X1 MEM_stage_inst_dmem_U12076 ( .A1(MEM_stage_inst_dmem_n14989), .A2(MEM_stage_inst_dmem_n14988), .ZN(MEM_stage_inst_dmem_n11779) );
NAND2_X1 MEM_stage_inst_dmem_U12075 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n15005), .ZN(MEM_stage_inst_dmem_n14988) );
NAND2_X1 MEM_stage_inst_dmem_U12074 ( .A1(MEM_stage_inst_dmem_ram_1480), .A2(MEM_stage_inst_dmem_n15004), .ZN(MEM_stage_inst_dmem_n14989) );
NAND2_X1 MEM_stage_inst_dmem_U12073 ( .A1(MEM_stage_inst_dmem_n14987), .A2(MEM_stage_inst_dmem_n14986), .ZN(MEM_stage_inst_dmem_n11780) );
NAND2_X1 MEM_stage_inst_dmem_U12072 ( .A1(MEM_stage_inst_dmem_n19251), .A2(MEM_stage_inst_dmem_n15005), .ZN(MEM_stage_inst_dmem_n14986) );
NAND2_X1 MEM_stage_inst_dmem_U12071 ( .A1(MEM_stage_inst_dmem_ram_1481), .A2(MEM_stage_inst_dmem_n15004), .ZN(MEM_stage_inst_dmem_n14987) );
NAND2_X1 MEM_stage_inst_dmem_U12070 ( .A1(MEM_stage_inst_dmem_n14985), .A2(MEM_stage_inst_dmem_n14984), .ZN(MEM_stage_inst_dmem_n11781) );
NAND2_X1 MEM_stage_inst_dmem_U12069 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n15005), .ZN(MEM_stage_inst_dmem_n14984) );
NAND2_X1 MEM_stage_inst_dmem_U12068 ( .A1(MEM_stage_inst_dmem_ram_1482), .A2(MEM_stage_inst_dmem_n15004), .ZN(MEM_stage_inst_dmem_n14985) );
NAND2_X1 MEM_stage_inst_dmem_U12067 ( .A1(MEM_stage_inst_dmem_n14983), .A2(MEM_stage_inst_dmem_n14982), .ZN(MEM_stage_inst_dmem_n11782) );
NAND2_X1 MEM_stage_inst_dmem_U12066 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n15005), .ZN(MEM_stage_inst_dmem_n14982) );
NAND2_X1 MEM_stage_inst_dmem_U12065 ( .A1(MEM_stage_inst_dmem_ram_1483), .A2(MEM_stage_inst_dmem_n15004), .ZN(MEM_stage_inst_dmem_n14983) );
NAND2_X1 MEM_stage_inst_dmem_U12064 ( .A1(MEM_stage_inst_dmem_n14981), .A2(MEM_stage_inst_dmem_n14980), .ZN(MEM_stage_inst_dmem_n11783) );
NAND2_X1 MEM_stage_inst_dmem_U12063 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n15005), .ZN(MEM_stage_inst_dmem_n14980) );
NAND2_X1 MEM_stage_inst_dmem_U12062 ( .A1(MEM_stage_inst_dmem_ram_1484), .A2(MEM_stage_inst_dmem_n15004), .ZN(MEM_stage_inst_dmem_n14981) );
NAND2_X1 MEM_stage_inst_dmem_U12061 ( .A1(MEM_stage_inst_dmem_n14979), .A2(MEM_stage_inst_dmem_n14978), .ZN(MEM_stage_inst_dmem_n11784) );
NAND2_X1 MEM_stage_inst_dmem_U12060 ( .A1(MEM_stage_inst_dmem_n15116), .A2(MEM_stage_inst_dmem_n15005), .ZN(MEM_stage_inst_dmem_n14978) );
NAND2_X1 MEM_stage_inst_dmem_U12059 ( .A1(MEM_stage_inst_dmem_ram_1485), .A2(MEM_stage_inst_dmem_n15004), .ZN(MEM_stage_inst_dmem_n14979) );
NAND2_X1 MEM_stage_inst_dmem_U12058 ( .A1(MEM_stage_inst_dmem_n14977), .A2(MEM_stage_inst_dmem_n14976), .ZN(MEM_stage_inst_dmem_n11785) );
NAND2_X1 MEM_stage_inst_dmem_U12057 ( .A1(MEM_stage_inst_dmem_n15113), .A2(MEM_stage_inst_dmem_n15005), .ZN(MEM_stage_inst_dmem_n14976) );
NAND2_X1 MEM_stage_inst_dmem_U12056 ( .A1(MEM_stage_inst_dmem_ram_1486), .A2(MEM_stage_inst_dmem_n15004), .ZN(MEM_stage_inst_dmem_n14977) );
NAND2_X1 MEM_stage_inst_dmem_U12055 ( .A1(MEM_stage_inst_dmem_n14975), .A2(MEM_stage_inst_dmem_n14974), .ZN(MEM_stage_inst_dmem_n11786) );
NAND2_X1 MEM_stage_inst_dmem_U12054 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n15005), .ZN(MEM_stage_inst_dmem_n14974) );
INV_X1 MEM_stage_inst_dmem_U12053 ( .A(MEM_stage_inst_dmem_n15004), .ZN(MEM_stage_inst_dmem_n15005) );
NAND2_X1 MEM_stage_inst_dmem_U12052 ( .A1(MEM_stage_inst_dmem_ram_1487), .A2(MEM_stage_inst_dmem_n15004), .ZN(MEM_stage_inst_dmem_n14975) );
NAND2_X1 MEM_stage_inst_dmem_U12051 ( .A1(MEM_stage_inst_dmem_n21039), .A2(MEM_stage_inst_dmem_n15386), .ZN(MEM_stage_inst_dmem_n15004) );
NAND2_X1 MEM_stage_inst_dmem_U12050 ( .A1(MEM_stage_inst_dmem_n14973), .A2(MEM_stage_inst_dmem_n14972), .ZN(MEM_stage_inst_dmem_n11787) );
NAND2_X1 MEM_stage_inst_dmem_U12049 ( .A1(MEM_stage_inst_dmem_n15145), .A2(MEM_stage_inst_dmem_n14971), .ZN(MEM_stage_inst_dmem_n14972) );
NAND2_X1 MEM_stage_inst_dmem_U12048 ( .A1(MEM_stage_inst_dmem_ram_1488), .A2(MEM_stage_inst_dmem_n14970), .ZN(MEM_stage_inst_dmem_n14973) );
NAND2_X1 MEM_stage_inst_dmem_U12047 ( .A1(MEM_stage_inst_dmem_n14969), .A2(MEM_stage_inst_dmem_n14968), .ZN(MEM_stage_inst_dmem_n11788) );
NAND2_X1 MEM_stage_inst_dmem_U12046 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n14971), .ZN(MEM_stage_inst_dmem_n14968) );
NAND2_X1 MEM_stage_inst_dmem_U12045 ( .A1(MEM_stage_inst_dmem_ram_1489), .A2(MEM_stage_inst_dmem_n14970), .ZN(MEM_stage_inst_dmem_n14969) );
NAND2_X1 MEM_stage_inst_dmem_U12044 ( .A1(MEM_stage_inst_dmem_n14967), .A2(MEM_stage_inst_dmem_n14966), .ZN(MEM_stage_inst_dmem_n11789) );
NAND2_X1 MEM_stage_inst_dmem_U12043 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n14971), .ZN(MEM_stage_inst_dmem_n14966) );
NAND2_X1 MEM_stage_inst_dmem_U12042 ( .A1(MEM_stage_inst_dmem_ram_1490), .A2(MEM_stage_inst_dmem_n14970), .ZN(MEM_stage_inst_dmem_n14967) );
NAND2_X1 MEM_stage_inst_dmem_U12041 ( .A1(MEM_stage_inst_dmem_n14965), .A2(MEM_stage_inst_dmem_n14964), .ZN(MEM_stage_inst_dmem_n11790) );
NAND2_X1 MEM_stage_inst_dmem_U12040 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n14971), .ZN(MEM_stage_inst_dmem_n14964) );
NAND2_X1 MEM_stage_inst_dmem_U12039 ( .A1(MEM_stage_inst_dmem_ram_1491), .A2(MEM_stage_inst_dmem_n14970), .ZN(MEM_stage_inst_dmem_n14965) );
NAND2_X1 MEM_stage_inst_dmem_U12038 ( .A1(MEM_stage_inst_dmem_n14963), .A2(MEM_stage_inst_dmem_n14962), .ZN(MEM_stage_inst_dmem_n11791) );
NAND2_X1 MEM_stage_inst_dmem_U12037 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n14971), .ZN(MEM_stage_inst_dmem_n14962) );
NAND2_X1 MEM_stage_inst_dmem_U12036 ( .A1(MEM_stage_inst_dmem_ram_1492), .A2(MEM_stage_inst_dmem_n14970), .ZN(MEM_stage_inst_dmem_n14963) );
NAND2_X1 MEM_stage_inst_dmem_U12035 ( .A1(MEM_stage_inst_dmem_n14961), .A2(MEM_stage_inst_dmem_n14960), .ZN(MEM_stage_inst_dmem_n11792) );
NAND2_X1 MEM_stage_inst_dmem_U12034 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n14971), .ZN(MEM_stage_inst_dmem_n14960) );
NAND2_X1 MEM_stage_inst_dmem_U12033 ( .A1(MEM_stage_inst_dmem_ram_1493), .A2(MEM_stage_inst_dmem_n14970), .ZN(MEM_stage_inst_dmem_n14961) );
NAND2_X1 MEM_stage_inst_dmem_U12032 ( .A1(MEM_stage_inst_dmem_n14959), .A2(MEM_stage_inst_dmem_n14958), .ZN(MEM_stage_inst_dmem_n11793) );
NAND2_X1 MEM_stage_inst_dmem_U12031 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n14971), .ZN(MEM_stage_inst_dmem_n14958) );
NAND2_X1 MEM_stage_inst_dmem_U12030 ( .A1(MEM_stage_inst_dmem_ram_1494), .A2(MEM_stage_inst_dmem_n14970), .ZN(MEM_stage_inst_dmem_n14959) );
NAND2_X1 MEM_stage_inst_dmem_U12029 ( .A1(MEM_stage_inst_dmem_n14957), .A2(MEM_stage_inst_dmem_n14956), .ZN(MEM_stage_inst_dmem_n11794) );
NAND2_X1 MEM_stage_inst_dmem_U12028 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n14971), .ZN(MEM_stage_inst_dmem_n14956) );
NAND2_X1 MEM_stage_inst_dmem_U12027 ( .A1(MEM_stage_inst_dmem_ram_1495), .A2(MEM_stage_inst_dmem_n14970), .ZN(MEM_stage_inst_dmem_n14957) );
NAND2_X1 MEM_stage_inst_dmem_U12026 ( .A1(MEM_stage_inst_dmem_n14955), .A2(MEM_stage_inst_dmem_n14954), .ZN(MEM_stage_inst_dmem_n11795) );
NAND2_X1 MEM_stage_inst_dmem_U12025 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n14971), .ZN(MEM_stage_inst_dmem_n14954) );
NAND2_X1 MEM_stage_inst_dmem_U12024 ( .A1(MEM_stage_inst_dmem_ram_1496), .A2(MEM_stage_inst_dmem_n14970), .ZN(MEM_stage_inst_dmem_n14955) );
NAND2_X1 MEM_stage_inst_dmem_U12023 ( .A1(MEM_stage_inst_dmem_n14953), .A2(MEM_stage_inst_dmem_n14952), .ZN(MEM_stage_inst_dmem_n11796) );
NAND2_X1 MEM_stage_inst_dmem_U12022 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n14971), .ZN(MEM_stage_inst_dmem_n14952) );
NAND2_X1 MEM_stage_inst_dmem_U12021 ( .A1(MEM_stage_inst_dmem_ram_1497), .A2(MEM_stage_inst_dmem_n14970), .ZN(MEM_stage_inst_dmem_n14953) );
NAND2_X1 MEM_stage_inst_dmem_U12020 ( .A1(MEM_stage_inst_dmem_n14951), .A2(MEM_stage_inst_dmem_n14950), .ZN(MEM_stage_inst_dmem_n11797) );
NAND2_X1 MEM_stage_inst_dmem_U12019 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n14971), .ZN(MEM_stage_inst_dmem_n14950) );
NAND2_X1 MEM_stage_inst_dmem_U12018 ( .A1(MEM_stage_inst_dmem_ram_1498), .A2(MEM_stage_inst_dmem_n14970), .ZN(MEM_stage_inst_dmem_n14951) );
NAND2_X1 MEM_stage_inst_dmem_U12017 ( .A1(MEM_stage_inst_dmem_n14949), .A2(MEM_stage_inst_dmem_n14948), .ZN(MEM_stage_inst_dmem_n11798) );
NAND2_X1 MEM_stage_inst_dmem_U12016 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n14971), .ZN(MEM_stage_inst_dmem_n14948) );
NAND2_X1 MEM_stage_inst_dmem_U12015 ( .A1(MEM_stage_inst_dmem_ram_1499), .A2(MEM_stage_inst_dmem_n14970), .ZN(MEM_stage_inst_dmem_n14949) );
NAND2_X1 MEM_stage_inst_dmem_U12014 ( .A1(MEM_stage_inst_dmem_n14947), .A2(MEM_stage_inst_dmem_n14946), .ZN(MEM_stage_inst_dmem_n11799) );
NAND2_X1 MEM_stage_inst_dmem_U12013 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n14971), .ZN(MEM_stage_inst_dmem_n14946) );
NAND2_X1 MEM_stage_inst_dmem_U12012 ( .A1(MEM_stage_inst_dmem_ram_1500), .A2(MEM_stage_inst_dmem_n14970), .ZN(MEM_stage_inst_dmem_n14947) );
NAND2_X1 MEM_stage_inst_dmem_U12011 ( .A1(MEM_stage_inst_dmem_n14945), .A2(MEM_stage_inst_dmem_n14944), .ZN(MEM_stage_inst_dmem_n11800) );
NAND2_X1 MEM_stage_inst_dmem_U12010 ( .A1(MEM_stage_inst_dmem_n15116), .A2(MEM_stage_inst_dmem_n14971), .ZN(MEM_stage_inst_dmem_n14944) );
NAND2_X1 MEM_stage_inst_dmem_U12009 ( .A1(MEM_stage_inst_dmem_ram_1501), .A2(MEM_stage_inst_dmem_n14970), .ZN(MEM_stage_inst_dmem_n14945) );
NAND2_X1 MEM_stage_inst_dmem_U12008 ( .A1(MEM_stage_inst_dmem_n14943), .A2(MEM_stage_inst_dmem_n14942), .ZN(MEM_stage_inst_dmem_n11801) );
NAND2_X1 MEM_stage_inst_dmem_U12007 ( .A1(MEM_stage_inst_dmem_n15113), .A2(MEM_stage_inst_dmem_n14971), .ZN(MEM_stage_inst_dmem_n14942) );
NAND2_X1 MEM_stage_inst_dmem_U12006 ( .A1(MEM_stage_inst_dmem_ram_1502), .A2(MEM_stage_inst_dmem_n14970), .ZN(MEM_stage_inst_dmem_n14943) );
NAND2_X1 MEM_stage_inst_dmem_U12005 ( .A1(MEM_stage_inst_dmem_n14941), .A2(MEM_stage_inst_dmem_n14940), .ZN(MEM_stage_inst_dmem_n11802) );
NAND2_X1 MEM_stage_inst_dmem_U12004 ( .A1(MEM_stage_inst_dmem_n16343), .A2(MEM_stage_inst_dmem_n14971), .ZN(MEM_stage_inst_dmem_n14940) );
INV_X1 MEM_stage_inst_dmem_U12003 ( .A(MEM_stage_inst_dmem_n14970), .ZN(MEM_stage_inst_dmem_n14971) );
NAND2_X1 MEM_stage_inst_dmem_U12002 ( .A1(MEM_stage_inst_dmem_ram_1503), .A2(MEM_stage_inst_dmem_n14970), .ZN(MEM_stage_inst_dmem_n14941) );
NAND2_X1 MEM_stage_inst_dmem_U12001 ( .A1(MEM_stage_inst_dmem_n21004), .A2(MEM_stage_inst_dmem_n15386), .ZN(MEM_stage_inst_dmem_n14970) );
NAND2_X1 MEM_stage_inst_dmem_U12000 ( .A1(MEM_stage_inst_dmem_n14939), .A2(MEM_stage_inst_dmem_n14938), .ZN(MEM_stage_inst_dmem_n11803) );
NAND2_X1 MEM_stage_inst_dmem_U11999 ( .A1(MEM_stage_inst_dmem_n15145), .A2(MEM_stage_inst_dmem_n14937), .ZN(MEM_stage_inst_dmem_n14938) );
NAND2_X1 MEM_stage_inst_dmem_U11998 ( .A1(MEM_stage_inst_dmem_ram_1504), .A2(MEM_stage_inst_dmem_n14936), .ZN(MEM_stage_inst_dmem_n14939) );
NAND2_X1 MEM_stage_inst_dmem_U11997 ( .A1(MEM_stage_inst_dmem_n14935), .A2(MEM_stage_inst_dmem_n14934), .ZN(MEM_stage_inst_dmem_n11804) );
NAND2_X1 MEM_stage_inst_dmem_U11996 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n14937), .ZN(MEM_stage_inst_dmem_n14934) );
NAND2_X1 MEM_stage_inst_dmem_U11995 ( .A1(MEM_stage_inst_dmem_ram_1505), .A2(MEM_stage_inst_dmem_n14936), .ZN(MEM_stage_inst_dmem_n14935) );
NAND2_X1 MEM_stage_inst_dmem_U11994 ( .A1(MEM_stage_inst_dmem_n14933), .A2(MEM_stage_inst_dmem_n14932), .ZN(MEM_stage_inst_dmem_n11805) );
NAND2_X1 MEM_stage_inst_dmem_U11993 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n14937), .ZN(MEM_stage_inst_dmem_n14932) );
NAND2_X1 MEM_stage_inst_dmem_U11992 ( .A1(MEM_stage_inst_dmem_ram_1506), .A2(MEM_stage_inst_dmem_n14936), .ZN(MEM_stage_inst_dmem_n14933) );
NAND2_X1 MEM_stage_inst_dmem_U11991 ( .A1(MEM_stage_inst_dmem_n14931), .A2(MEM_stage_inst_dmem_n14930), .ZN(MEM_stage_inst_dmem_n11806) );
NAND2_X1 MEM_stage_inst_dmem_U11990 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n14937), .ZN(MEM_stage_inst_dmem_n14930) );
NAND2_X1 MEM_stage_inst_dmem_U11989 ( .A1(MEM_stage_inst_dmem_ram_1507), .A2(MEM_stage_inst_dmem_n14936), .ZN(MEM_stage_inst_dmem_n14931) );
NAND2_X1 MEM_stage_inst_dmem_U11988 ( .A1(MEM_stage_inst_dmem_n14929), .A2(MEM_stage_inst_dmem_n14928), .ZN(MEM_stage_inst_dmem_n11807) );
NAND2_X1 MEM_stage_inst_dmem_U11987 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n14937), .ZN(MEM_stage_inst_dmem_n14928) );
NAND2_X1 MEM_stage_inst_dmem_U11986 ( .A1(MEM_stage_inst_dmem_ram_1508), .A2(MEM_stage_inst_dmem_n14936), .ZN(MEM_stage_inst_dmem_n14929) );
NAND2_X1 MEM_stage_inst_dmem_U11985 ( .A1(MEM_stage_inst_dmem_n14927), .A2(MEM_stage_inst_dmem_n14926), .ZN(MEM_stage_inst_dmem_n11808) );
NAND2_X1 MEM_stage_inst_dmem_U11984 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n14937), .ZN(MEM_stage_inst_dmem_n14926) );
NAND2_X1 MEM_stage_inst_dmem_U11983 ( .A1(MEM_stage_inst_dmem_ram_1509), .A2(MEM_stage_inst_dmem_n14936), .ZN(MEM_stage_inst_dmem_n14927) );
NAND2_X1 MEM_stage_inst_dmem_U11982 ( .A1(MEM_stage_inst_dmem_n14925), .A2(MEM_stage_inst_dmem_n14924), .ZN(MEM_stage_inst_dmem_n11809) );
NAND2_X1 MEM_stage_inst_dmem_U11981 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n14937), .ZN(MEM_stage_inst_dmem_n14924) );
NAND2_X1 MEM_stage_inst_dmem_U11980 ( .A1(MEM_stage_inst_dmem_ram_1510), .A2(MEM_stage_inst_dmem_n14936), .ZN(MEM_stage_inst_dmem_n14925) );
NAND2_X1 MEM_stage_inst_dmem_U11979 ( .A1(MEM_stage_inst_dmem_n14923), .A2(MEM_stage_inst_dmem_n14922), .ZN(MEM_stage_inst_dmem_n11810) );
NAND2_X1 MEM_stage_inst_dmem_U11978 ( .A1(MEM_stage_inst_dmem_n16361), .A2(MEM_stage_inst_dmem_n14937), .ZN(MEM_stage_inst_dmem_n14922) );
NAND2_X1 MEM_stage_inst_dmem_U11977 ( .A1(MEM_stage_inst_dmem_ram_1511), .A2(MEM_stage_inst_dmem_n14936), .ZN(MEM_stage_inst_dmem_n14923) );
NAND2_X1 MEM_stage_inst_dmem_U11976 ( .A1(MEM_stage_inst_dmem_n14921), .A2(MEM_stage_inst_dmem_n14920), .ZN(MEM_stage_inst_dmem_n11811) );
NAND2_X1 MEM_stage_inst_dmem_U11975 ( .A1(MEM_stage_inst_dmem_n18013), .A2(MEM_stage_inst_dmem_n14937), .ZN(MEM_stage_inst_dmem_n14920) );
NAND2_X1 MEM_stage_inst_dmem_U11974 ( .A1(MEM_stage_inst_dmem_ram_1512), .A2(MEM_stage_inst_dmem_n14936), .ZN(MEM_stage_inst_dmem_n14921) );
NAND2_X1 MEM_stage_inst_dmem_U11973 ( .A1(MEM_stage_inst_dmem_n14919), .A2(MEM_stage_inst_dmem_n14918), .ZN(MEM_stage_inst_dmem_n11812) );
NAND2_X1 MEM_stage_inst_dmem_U11972 ( .A1(MEM_stage_inst_dmem_n19251), .A2(MEM_stage_inst_dmem_n14937), .ZN(MEM_stage_inst_dmem_n14918) );
NAND2_X1 MEM_stage_inst_dmem_U11971 ( .A1(MEM_stage_inst_dmem_ram_1513), .A2(MEM_stage_inst_dmem_n14936), .ZN(MEM_stage_inst_dmem_n14919) );
NAND2_X1 MEM_stage_inst_dmem_U11970 ( .A1(MEM_stage_inst_dmem_n14917), .A2(MEM_stage_inst_dmem_n14916), .ZN(MEM_stage_inst_dmem_n11813) );
NAND2_X1 MEM_stage_inst_dmem_U11969 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n14937), .ZN(MEM_stage_inst_dmem_n14916) );
NAND2_X1 MEM_stage_inst_dmem_U11968 ( .A1(MEM_stage_inst_dmem_ram_1514), .A2(MEM_stage_inst_dmem_n14936), .ZN(MEM_stage_inst_dmem_n14917) );
NAND2_X1 MEM_stage_inst_dmem_U11967 ( .A1(MEM_stage_inst_dmem_n14915), .A2(MEM_stage_inst_dmem_n14914), .ZN(MEM_stage_inst_dmem_n11814) );
NAND2_X1 MEM_stage_inst_dmem_U11966 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n14937), .ZN(MEM_stage_inst_dmem_n14914) );
NAND2_X1 MEM_stage_inst_dmem_U11965 ( .A1(MEM_stage_inst_dmem_ram_1515), .A2(MEM_stage_inst_dmem_n14936), .ZN(MEM_stage_inst_dmem_n14915) );
NAND2_X1 MEM_stage_inst_dmem_U11964 ( .A1(MEM_stage_inst_dmem_n14913), .A2(MEM_stage_inst_dmem_n14912), .ZN(MEM_stage_inst_dmem_n11815) );
NAND2_X1 MEM_stage_inst_dmem_U11963 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n14937), .ZN(MEM_stage_inst_dmem_n14912) );
NAND2_X1 MEM_stage_inst_dmem_U11962 ( .A1(MEM_stage_inst_dmem_ram_1516), .A2(MEM_stage_inst_dmem_n14936), .ZN(MEM_stage_inst_dmem_n14913) );
NAND2_X1 MEM_stage_inst_dmem_U11961 ( .A1(MEM_stage_inst_dmem_n14911), .A2(MEM_stage_inst_dmem_n14910), .ZN(MEM_stage_inst_dmem_n11816) );
NAND2_X1 MEM_stage_inst_dmem_U11960 ( .A1(MEM_stage_inst_dmem_n15116), .A2(MEM_stage_inst_dmem_n14937), .ZN(MEM_stage_inst_dmem_n14910) );
NAND2_X1 MEM_stage_inst_dmem_U11959 ( .A1(MEM_stage_inst_dmem_ram_1517), .A2(MEM_stage_inst_dmem_n14936), .ZN(MEM_stage_inst_dmem_n14911) );
NAND2_X1 MEM_stage_inst_dmem_U11958 ( .A1(MEM_stage_inst_dmem_n14909), .A2(MEM_stage_inst_dmem_n14908), .ZN(MEM_stage_inst_dmem_n11817) );
NAND2_X1 MEM_stage_inst_dmem_U11957 ( .A1(MEM_stage_inst_dmem_n15113), .A2(MEM_stage_inst_dmem_n14937), .ZN(MEM_stage_inst_dmem_n14908) );
NAND2_X1 MEM_stage_inst_dmem_U11956 ( .A1(MEM_stage_inst_dmem_ram_1518), .A2(MEM_stage_inst_dmem_n14936), .ZN(MEM_stage_inst_dmem_n14909) );
NAND2_X1 MEM_stage_inst_dmem_U11955 ( .A1(MEM_stage_inst_dmem_n14907), .A2(MEM_stage_inst_dmem_n14906), .ZN(MEM_stage_inst_dmem_n11818) );
NAND2_X1 MEM_stage_inst_dmem_U11954 ( .A1(MEM_stage_inst_dmem_n14693), .A2(MEM_stage_inst_dmem_n14937), .ZN(MEM_stage_inst_dmem_n14906) );
NAND2_X1 MEM_stage_inst_dmem_U11953 ( .A1(MEM_stage_inst_dmem_ram_1519), .A2(MEM_stage_inst_dmem_n14936), .ZN(MEM_stage_inst_dmem_n14907) );
NAND2_X1 MEM_stage_inst_dmem_U11952 ( .A1(MEM_stage_inst_dmem_n20969), .A2(MEM_stage_inst_dmem_n15386), .ZN(MEM_stage_inst_dmem_n14936) );
NAND2_X1 MEM_stage_inst_dmem_U11951 ( .A1(MEM_stage_inst_dmem_n14905), .A2(MEM_stage_inst_dmem_n14904), .ZN(MEM_stage_inst_dmem_n11819) );
NAND2_X1 MEM_stage_inst_dmem_U11950 ( .A1(MEM_stage_inst_dmem_n15145), .A2(MEM_stage_inst_dmem_n14903), .ZN(MEM_stage_inst_dmem_n14904) );
NAND2_X1 MEM_stage_inst_dmem_U11949 ( .A1(MEM_stage_inst_dmem_ram_1520), .A2(MEM_stage_inst_dmem_n14902), .ZN(MEM_stage_inst_dmem_n14905) );
NAND2_X1 MEM_stage_inst_dmem_U11948 ( .A1(MEM_stage_inst_dmem_n14901), .A2(MEM_stage_inst_dmem_n14900), .ZN(MEM_stage_inst_dmem_n11820) );
NAND2_X1 MEM_stage_inst_dmem_U11947 ( .A1(MEM_stage_inst_dmem_n109), .A2(MEM_stage_inst_dmem_n14903), .ZN(MEM_stage_inst_dmem_n14900) );
NAND2_X1 MEM_stage_inst_dmem_U11946 ( .A1(MEM_stage_inst_dmem_ram_1521), .A2(MEM_stage_inst_dmem_n14902), .ZN(MEM_stage_inst_dmem_n14901) );
NAND2_X1 MEM_stage_inst_dmem_U11945 ( .A1(MEM_stage_inst_dmem_n14899), .A2(MEM_stage_inst_dmem_n14898), .ZN(MEM_stage_inst_dmem_n11821) );
NAND2_X1 MEM_stage_inst_dmem_U11944 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n14903), .ZN(MEM_stage_inst_dmem_n14898) );
NAND2_X1 MEM_stage_inst_dmem_U11943 ( .A1(MEM_stage_inst_dmem_ram_1522), .A2(MEM_stage_inst_dmem_n14902), .ZN(MEM_stage_inst_dmem_n14899) );
NAND2_X1 MEM_stage_inst_dmem_U11942 ( .A1(MEM_stage_inst_dmem_n14897), .A2(MEM_stage_inst_dmem_n14896), .ZN(MEM_stage_inst_dmem_n11822) );
NAND2_X1 MEM_stage_inst_dmem_U11941 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n14903), .ZN(MEM_stage_inst_dmem_n14896) );
NAND2_X1 MEM_stage_inst_dmem_U11940 ( .A1(MEM_stage_inst_dmem_ram_1523), .A2(MEM_stage_inst_dmem_n14902), .ZN(MEM_stage_inst_dmem_n14897) );
NAND2_X1 MEM_stage_inst_dmem_U11939 ( .A1(MEM_stage_inst_dmem_n14895), .A2(MEM_stage_inst_dmem_n14894), .ZN(MEM_stage_inst_dmem_n11823) );
NAND2_X1 MEM_stage_inst_dmem_U11938 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n14903), .ZN(MEM_stage_inst_dmem_n14894) );
NAND2_X1 MEM_stage_inst_dmem_U11937 ( .A1(MEM_stage_inst_dmem_ram_1524), .A2(MEM_stage_inst_dmem_n14902), .ZN(MEM_stage_inst_dmem_n14895) );
NAND2_X1 MEM_stage_inst_dmem_U11936 ( .A1(MEM_stage_inst_dmem_n14893), .A2(MEM_stage_inst_dmem_n14892), .ZN(MEM_stage_inst_dmem_n11824) );
NAND2_X1 MEM_stage_inst_dmem_U11935 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n14903), .ZN(MEM_stage_inst_dmem_n14892) );
NAND2_X1 MEM_stage_inst_dmem_U11934 ( .A1(MEM_stage_inst_dmem_ram_1525), .A2(MEM_stage_inst_dmem_n14902), .ZN(MEM_stage_inst_dmem_n14893) );
NAND2_X1 MEM_stage_inst_dmem_U11933 ( .A1(MEM_stage_inst_dmem_n14891), .A2(MEM_stage_inst_dmem_n14890), .ZN(MEM_stage_inst_dmem_n11825) );
NAND2_X1 MEM_stage_inst_dmem_U11932 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n14903), .ZN(MEM_stage_inst_dmem_n14890) );
NAND2_X1 MEM_stage_inst_dmem_U11931 ( .A1(MEM_stage_inst_dmem_ram_1526), .A2(MEM_stage_inst_dmem_n14902), .ZN(MEM_stage_inst_dmem_n14891) );
NAND2_X1 MEM_stage_inst_dmem_U11930 ( .A1(MEM_stage_inst_dmem_n14889), .A2(MEM_stage_inst_dmem_n14888), .ZN(MEM_stage_inst_dmem_n11826) );
NAND2_X1 MEM_stage_inst_dmem_U11929 ( .A1(MEM_stage_inst_dmem_n112), .A2(MEM_stage_inst_dmem_n14903), .ZN(MEM_stage_inst_dmem_n14888) );
NAND2_X1 MEM_stage_inst_dmem_U11928 ( .A1(MEM_stage_inst_dmem_ram_1527), .A2(MEM_stage_inst_dmem_n14902), .ZN(MEM_stage_inst_dmem_n14889) );
NAND2_X1 MEM_stage_inst_dmem_U11927 ( .A1(MEM_stage_inst_dmem_n14887), .A2(MEM_stage_inst_dmem_n14886), .ZN(MEM_stage_inst_dmem_n11827) );
NAND2_X1 MEM_stage_inst_dmem_U11926 ( .A1(EX_pipeline_reg_out_13), .A2(MEM_stage_inst_dmem_n14903), .ZN(MEM_stage_inst_dmem_n14886) );
NAND2_X1 MEM_stage_inst_dmem_U11925 ( .A1(MEM_stage_inst_dmem_ram_1528), .A2(MEM_stage_inst_dmem_n14902), .ZN(MEM_stage_inst_dmem_n14887) );
NAND2_X1 MEM_stage_inst_dmem_U11924 ( .A1(MEM_stage_inst_dmem_n14885), .A2(MEM_stage_inst_dmem_n14884), .ZN(MEM_stage_inst_dmem_n11828) );
NAND2_X1 MEM_stage_inst_dmem_U11923 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n14903), .ZN(MEM_stage_inst_dmem_n14884) );
NAND2_X1 MEM_stage_inst_dmem_U11922 ( .A1(MEM_stage_inst_dmem_ram_1529), .A2(MEM_stage_inst_dmem_n14902), .ZN(MEM_stage_inst_dmem_n14885) );
NAND2_X1 MEM_stage_inst_dmem_U11921 ( .A1(MEM_stage_inst_dmem_n14883), .A2(MEM_stage_inst_dmem_n14882), .ZN(MEM_stage_inst_dmem_n11829) );
NAND2_X1 MEM_stage_inst_dmem_U11920 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n14903), .ZN(MEM_stage_inst_dmem_n14882) );
NAND2_X1 MEM_stage_inst_dmem_U11919 ( .A1(MEM_stage_inst_dmem_ram_1530), .A2(MEM_stage_inst_dmem_n14902), .ZN(MEM_stage_inst_dmem_n14883) );
NAND2_X1 MEM_stage_inst_dmem_U11918 ( .A1(MEM_stage_inst_dmem_n14881), .A2(MEM_stage_inst_dmem_n14880), .ZN(MEM_stage_inst_dmem_n11830) );
NAND2_X1 MEM_stage_inst_dmem_U11917 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n14903), .ZN(MEM_stage_inst_dmem_n14880) );
NAND2_X1 MEM_stage_inst_dmem_U11916 ( .A1(MEM_stage_inst_dmem_ram_1531), .A2(MEM_stage_inst_dmem_n14902), .ZN(MEM_stage_inst_dmem_n14881) );
NAND2_X1 MEM_stage_inst_dmem_U11915 ( .A1(MEM_stage_inst_dmem_n14879), .A2(MEM_stage_inst_dmem_n14878), .ZN(MEM_stage_inst_dmem_n11831) );
NAND2_X1 MEM_stage_inst_dmem_U11914 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n14903), .ZN(MEM_stage_inst_dmem_n14878) );
NAND2_X1 MEM_stage_inst_dmem_U11913 ( .A1(MEM_stage_inst_dmem_ram_1532), .A2(MEM_stage_inst_dmem_n14902), .ZN(MEM_stage_inst_dmem_n14879) );
NAND2_X1 MEM_stage_inst_dmem_U11912 ( .A1(MEM_stage_inst_dmem_n14877), .A2(MEM_stage_inst_dmem_n14876), .ZN(MEM_stage_inst_dmem_n11832) );
NAND2_X1 MEM_stage_inst_dmem_U11911 ( .A1(MEM_stage_inst_dmem_n15116), .A2(MEM_stage_inst_dmem_n14903), .ZN(MEM_stage_inst_dmem_n14876) );
NAND2_X1 MEM_stage_inst_dmem_U11910 ( .A1(MEM_stage_inst_dmem_ram_1533), .A2(MEM_stage_inst_dmem_n14902), .ZN(MEM_stage_inst_dmem_n14877) );
NAND2_X1 MEM_stage_inst_dmem_U11909 ( .A1(MEM_stage_inst_dmem_n14875), .A2(MEM_stage_inst_dmem_n14874), .ZN(MEM_stage_inst_dmem_n11833) );
NAND2_X1 MEM_stage_inst_dmem_U11908 ( .A1(MEM_stage_inst_dmem_n15113), .A2(MEM_stage_inst_dmem_n14903), .ZN(MEM_stage_inst_dmem_n14874) );
NAND2_X1 MEM_stage_inst_dmem_U11907 ( .A1(MEM_stage_inst_dmem_ram_1534), .A2(MEM_stage_inst_dmem_n14902), .ZN(MEM_stage_inst_dmem_n14875) );
NAND2_X1 MEM_stage_inst_dmem_U11906 ( .A1(MEM_stage_inst_dmem_n14873), .A2(MEM_stage_inst_dmem_n14872), .ZN(MEM_stage_inst_dmem_n11834) );
NAND2_X1 MEM_stage_inst_dmem_U11905 ( .A1(MEM_stage_inst_dmem_n15110), .A2(MEM_stage_inst_dmem_n14903), .ZN(MEM_stage_inst_dmem_n14872) );
INV_X1 MEM_stage_inst_dmem_U11904 ( .A(MEM_stage_inst_dmem_n14902), .ZN(MEM_stage_inst_dmem_n14903) );
NAND2_X1 MEM_stage_inst_dmem_U11903 ( .A1(MEM_stage_inst_dmem_ram_1535), .A2(MEM_stage_inst_dmem_n14902), .ZN(MEM_stage_inst_dmem_n14873) );
NAND2_X1 MEM_stage_inst_dmem_U11902 ( .A1(MEM_stage_inst_dmem_n20934), .A2(MEM_stage_inst_dmem_n15386), .ZN(MEM_stage_inst_dmem_n14902) );
NOR2_X2 MEM_stage_inst_dmem_U11901 ( .A1(MEM_stage_inst_dmem_n15968), .A2(MEM_stage_inst_dmem_n19823), .ZN(MEM_stage_inst_dmem_n15386) );
NAND2_X1 MEM_stage_inst_dmem_U11900 ( .A1(EX_pipeline_reg_out_27), .A2(MEM_stage_inst_dmem_n15967), .ZN(MEM_stage_inst_dmem_n19823) );
NAND2_X1 MEM_stage_inst_dmem_U11899 ( .A1(MEM_stage_inst_dmem_n14871), .A2(MEM_stage_inst_dmem_n14870), .ZN(MEM_stage_inst_dmem_n11835) );
NAND2_X1 MEM_stage_inst_dmem_U11898 ( .A1(MEM_stage_inst_dmem_n15145), .A2(MEM_stage_inst_dmem_n14869), .ZN(MEM_stage_inst_dmem_n14870) );
NAND2_X1 MEM_stage_inst_dmem_U11897 ( .A1(MEM_stage_inst_dmem_ram_512), .A2(MEM_stage_inst_dmem_n14868), .ZN(MEM_stage_inst_dmem_n14871) );
NAND2_X1 MEM_stage_inst_dmem_U11896 ( .A1(MEM_stage_inst_dmem_n14867), .A2(MEM_stage_inst_dmem_n14866), .ZN(MEM_stage_inst_dmem_n11836) );
NAND2_X1 MEM_stage_inst_dmem_U11895 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n14869), .ZN(MEM_stage_inst_dmem_n14866) );
NAND2_X1 MEM_stage_inst_dmem_U11894 ( .A1(MEM_stage_inst_dmem_ram_513), .A2(MEM_stage_inst_dmem_n14868), .ZN(MEM_stage_inst_dmem_n14867) );
NAND2_X1 MEM_stage_inst_dmem_U11893 ( .A1(MEM_stage_inst_dmem_n14865), .A2(MEM_stage_inst_dmem_n14864), .ZN(MEM_stage_inst_dmem_n11837) );
NAND2_X1 MEM_stage_inst_dmem_U11892 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n14869), .ZN(MEM_stage_inst_dmem_n14864) );
NAND2_X1 MEM_stage_inst_dmem_U11891 ( .A1(MEM_stage_inst_dmem_ram_514), .A2(MEM_stage_inst_dmem_n14868), .ZN(MEM_stage_inst_dmem_n14865) );
NAND2_X1 MEM_stage_inst_dmem_U11890 ( .A1(MEM_stage_inst_dmem_n14863), .A2(MEM_stage_inst_dmem_n14862), .ZN(MEM_stage_inst_dmem_n11838) );
NAND2_X1 MEM_stage_inst_dmem_U11889 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n14869), .ZN(MEM_stage_inst_dmem_n14862) );
NAND2_X1 MEM_stage_inst_dmem_U11888 ( .A1(MEM_stage_inst_dmem_ram_515), .A2(MEM_stage_inst_dmem_n14868), .ZN(MEM_stage_inst_dmem_n14863) );
NAND2_X1 MEM_stage_inst_dmem_U11887 ( .A1(MEM_stage_inst_dmem_n14861), .A2(MEM_stage_inst_dmem_n14860), .ZN(MEM_stage_inst_dmem_n11839) );
NAND2_X1 MEM_stage_inst_dmem_U11886 ( .A1(MEM_stage_inst_dmem_n16368), .A2(MEM_stage_inst_dmem_n14869), .ZN(MEM_stage_inst_dmem_n14860) );
NAND2_X1 MEM_stage_inst_dmem_U11885 ( .A1(MEM_stage_inst_dmem_ram_516), .A2(MEM_stage_inst_dmem_n14868), .ZN(MEM_stage_inst_dmem_n14861) );
NAND2_X1 MEM_stage_inst_dmem_U11884 ( .A1(MEM_stage_inst_dmem_n14859), .A2(MEM_stage_inst_dmem_n14858), .ZN(MEM_stage_inst_dmem_n11840) );
NAND2_X1 MEM_stage_inst_dmem_U11883 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n14869), .ZN(MEM_stage_inst_dmem_n14858) );
NAND2_X1 MEM_stage_inst_dmem_U11882 ( .A1(MEM_stage_inst_dmem_ram_517), .A2(MEM_stage_inst_dmem_n14868), .ZN(MEM_stage_inst_dmem_n14859) );
NAND2_X1 MEM_stage_inst_dmem_U11881 ( .A1(MEM_stage_inst_dmem_n14857), .A2(MEM_stage_inst_dmem_n14856), .ZN(MEM_stage_inst_dmem_n11841) );
NAND2_X1 MEM_stage_inst_dmem_U11880 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n14869), .ZN(MEM_stage_inst_dmem_n14856) );
NAND2_X1 MEM_stage_inst_dmem_U11879 ( .A1(MEM_stage_inst_dmem_ram_518), .A2(MEM_stage_inst_dmem_n14868), .ZN(MEM_stage_inst_dmem_n14857) );
NAND2_X1 MEM_stage_inst_dmem_U11878 ( .A1(MEM_stage_inst_dmem_n14855), .A2(MEM_stage_inst_dmem_n14854), .ZN(MEM_stage_inst_dmem_n11842) );
NAND2_X1 MEM_stage_inst_dmem_U11877 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n14869), .ZN(MEM_stage_inst_dmem_n14854) );
NAND2_X1 MEM_stage_inst_dmem_U11876 ( .A1(MEM_stage_inst_dmem_ram_519), .A2(MEM_stage_inst_dmem_n14868), .ZN(MEM_stage_inst_dmem_n14855) );
NAND2_X1 MEM_stage_inst_dmem_U11875 ( .A1(MEM_stage_inst_dmem_n14853), .A2(MEM_stage_inst_dmem_n14852), .ZN(MEM_stage_inst_dmem_n11843) );
NAND2_X1 MEM_stage_inst_dmem_U11874 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n14869), .ZN(MEM_stage_inst_dmem_n14852) );
NAND2_X1 MEM_stage_inst_dmem_U11873 ( .A1(MEM_stage_inst_dmem_ram_520), .A2(MEM_stage_inst_dmem_n14868), .ZN(MEM_stage_inst_dmem_n14853) );
NAND2_X1 MEM_stage_inst_dmem_U11872 ( .A1(MEM_stage_inst_dmem_n14851), .A2(MEM_stage_inst_dmem_n14850), .ZN(MEM_stage_inst_dmem_n11844) );
NAND2_X1 MEM_stage_inst_dmem_U11871 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n14869), .ZN(MEM_stage_inst_dmem_n14850) );
NAND2_X1 MEM_stage_inst_dmem_U11870 ( .A1(MEM_stage_inst_dmem_ram_521), .A2(MEM_stage_inst_dmem_n14868), .ZN(MEM_stage_inst_dmem_n14851) );
NAND2_X1 MEM_stage_inst_dmem_U11869 ( .A1(MEM_stage_inst_dmem_n14849), .A2(MEM_stage_inst_dmem_n14848), .ZN(MEM_stage_inst_dmem_n11845) );
NAND2_X1 MEM_stage_inst_dmem_U11868 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n14869), .ZN(MEM_stage_inst_dmem_n14848) );
NAND2_X1 MEM_stage_inst_dmem_U11867 ( .A1(MEM_stage_inst_dmem_ram_522), .A2(MEM_stage_inst_dmem_n14868), .ZN(MEM_stage_inst_dmem_n14849) );
NAND2_X1 MEM_stage_inst_dmem_U11866 ( .A1(MEM_stage_inst_dmem_n14847), .A2(MEM_stage_inst_dmem_n14846), .ZN(MEM_stage_inst_dmem_n11846) );
NAND2_X1 MEM_stage_inst_dmem_U11865 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n14869), .ZN(MEM_stage_inst_dmem_n14846) );
NAND2_X1 MEM_stage_inst_dmem_U11864 ( .A1(MEM_stage_inst_dmem_ram_523), .A2(MEM_stage_inst_dmem_n14868), .ZN(MEM_stage_inst_dmem_n14847) );
NAND2_X1 MEM_stage_inst_dmem_U11863 ( .A1(MEM_stage_inst_dmem_n14845), .A2(MEM_stage_inst_dmem_n14844), .ZN(MEM_stage_inst_dmem_n11847) );
NAND2_X1 MEM_stage_inst_dmem_U11862 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n14869), .ZN(MEM_stage_inst_dmem_n14844) );
NAND2_X1 MEM_stage_inst_dmem_U11861 ( .A1(MEM_stage_inst_dmem_ram_524), .A2(MEM_stage_inst_dmem_n14868), .ZN(MEM_stage_inst_dmem_n14845) );
NAND2_X1 MEM_stage_inst_dmem_U11860 ( .A1(MEM_stage_inst_dmem_n14843), .A2(MEM_stage_inst_dmem_n14842), .ZN(MEM_stage_inst_dmem_n11848) );
NAND2_X1 MEM_stage_inst_dmem_U11859 ( .A1(MEM_stage_inst_dmem_n15116), .A2(MEM_stage_inst_dmem_n14869), .ZN(MEM_stage_inst_dmem_n14842) );
NAND2_X1 MEM_stage_inst_dmem_U11858 ( .A1(MEM_stage_inst_dmem_ram_525), .A2(MEM_stage_inst_dmem_n14868), .ZN(MEM_stage_inst_dmem_n14843) );
NAND2_X1 MEM_stage_inst_dmem_U11857 ( .A1(MEM_stage_inst_dmem_n14841), .A2(MEM_stage_inst_dmem_n14840), .ZN(MEM_stage_inst_dmem_n11849) );
NAND2_X1 MEM_stage_inst_dmem_U11856 ( .A1(MEM_stage_inst_dmem_n15113), .A2(MEM_stage_inst_dmem_n14869), .ZN(MEM_stage_inst_dmem_n14840) );
NAND2_X1 MEM_stage_inst_dmem_U11855 ( .A1(MEM_stage_inst_dmem_ram_526), .A2(MEM_stage_inst_dmem_n14868), .ZN(MEM_stage_inst_dmem_n14841) );
NAND2_X1 MEM_stage_inst_dmem_U11854 ( .A1(MEM_stage_inst_dmem_n14839), .A2(MEM_stage_inst_dmem_n14838), .ZN(MEM_stage_inst_dmem_n11850) );
NAND2_X1 MEM_stage_inst_dmem_U11853 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n14869), .ZN(MEM_stage_inst_dmem_n14838) );
INV_X1 MEM_stage_inst_dmem_U11852 ( .A(MEM_stage_inst_dmem_n14868), .ZN(MEM_stage_inst_dmem_n14869) );
NAND2_X1 MEM_stage_inst_dmem_U11851 ( .A1(MEM_stage_inst_dmem_ram_527), .A2(MEM_stage_inst_dmem_n14868), .ZN(MEM_stage_inst_dmem_n14839) );
NAND2_X1 MEM_stage_inst_dmem_U11850 ( .A1(MEM_stage_inst_dmem_n21465), .A2(MEM_stage_inst_dmem_n14837), .ZN(MEM_stage_inst_dmem_n14868) );
NAND2_X1 MEM_stage_inst_dmem_U11849 ( .A1(MEM_stage_inst_dmem_n14836), .A2(MEM_stage_inst_dmem_n14835), .ZN(MEM_stage_inst_dmem_n11851) );
NAND2_X1 MEM_stage_inst_dmem_U11848 ( .A1(MEM_stage_inst_dmem_n15145), .A2(MEM_stage_inst_dmem_n14834), .ZN(MEM_stage_inst_dmem_n14835) );
NAND2_X1 MEM_stage_inst_dmem_U11847 ( .A1(MEM_stage_inst_dmem_ram_528), .A2(MEM_stage_inst_dmem_n14833), .ZN(MEM_stage_inst_dmem_n14836) );
NAND2_X1 MEM_stage_inst_dmem_U11846 ( .A1(MEM_stage_inst_dmem_n14832), .A2(MEM_stage_inst_dmem_n14831), .ZN(MEM_stage_inst_dmem_n11852) );
NAND2_X1 MEM_stage_inst_dmem_U11845 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n14834), .ZN(MEM_stage_inst_dmem_n14831) );
NAND2_X1 MEM_stage_inst_dmem_U11844 ( .A1(MEM_stage_inst_dmem_ram_529), .A2(MEM_stage_inst_dmem_n14833), .ZN(MEM_stage_inst_dmem_n14832) );
NAND2_X1 MEM_stage_inst_dmem_U11843 ( .A1(MEM_stage_inst_dmem_n14830), .A2(MEM_stage_inst_dmem_n14829), .ZN(MEM_stage_inst_dmem_n11853) );
NAND2_X1 MEM_stage_inst_dmem_U11842 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n14834), .ZN(MEM_stage_inst_dmem_n14829) );
NAND2_X1 MEM_stage_inst_dmem_U11841 ( .A1(MEM_stage_inst_dmem_ram_530), .A2(MEM_stage_inst_dmem_n14833), .ZN(MEM_stage_inst_dmem_n14830) );
NAND2_X1 MEM_stage_inst_dmem_U11840 ( .A1(MEM_stage_inst_dmem_n14828), .A2(MEM_stage_inst_dmem_n14827), .ZN(MEM_stage_inst_dmem_n11854) );
NAND2_X1 MEM_stage_inst_dmem_U11839 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n14834), .ZN(MEM_stage_inst_dmem_n14827) );
NAND2_X1 MEM_stage_inst_dmem_U11838 ( .A1(MEM_stage_inst_dmem_ram_531), .A2(MEM_stage_inst_dmem_n14833), .ZN(MEM_stage_inst_dmem_n14828) );
NAND2_X1 MEM_stage_inst_dmem_U11837 ( .A1(MEM_stage_inst_dmem_n14826), .A2(MEM_stage_inst_dmem_n14825), .ZN(MEM_stage_inst_dmem_n11855) );
NAND2_X1 MEM_stage_inst_dmem_U11836 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n14834), .ZN(MEM_stage_inst_dmem_n14825) );
NAND2_X1 MEM_stage_inst_dmem_U11835 ( .A1(MEM_stage_inst_dmem_ram_532), .A2(MEM_stage_inst_dmem_n14833), .ZN(MEM_stage_inst_dmem_n14826) );
NAND2_X1 MEM_stage_inst_dmem_U11834 ( .A1(MEM_stage_inst_dmem_n14824), .A2(MEM_stage_inst_dmem_n14823), .ZN(MEM_stage_inst_dmem_n11856) );
NAND2_X1 MEM_stage_inst_dmem_U11833 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n14834), .ZN(MEM_stage_inst_dmem_n14823) );
NAND2_X1 MEM_stage_inst_dmem_U11832 ( .A1(MEM_stage_inst_dmem_ram_533), .A2(MEM_stage_inst_dmem_n14833), .ZN(MEM_stage_inst_dmem_n14824) );
NAND2_X1 MEM_stage_inst_dmem_U11831 ( .A1(MEM_stage_inst_dmem_n14822), .A2(MEM_stage_inst_dmem_n14821), .ZN(MEM_stage_inst_dmem_n11857) );
NAND2_X1 MEM_stage_inst_dmem_U11830 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n14834), .ZN(MEM_stage_inst_dmem_n14821) );
NAND2_X1 MEM_stage_inst_dmem_U11829 ( .A1(MEM_stage_inst_dmem_ram_534), .A2(MEM_stage_inst_dmem_n14833), .ZN(MEM_stage_inst_dmem_n14822) );
NAND2_X1 MEM_stage_inst_dmem_U11828 ( .A1(MEM_stage_inst_dmem_n14820), .A2(MEM_stage_inst_dmem_n14819), .ZN(MEM_stage_inst_dmem_n11858) );
NAND2_X1 MEM_stage_inst_dmem_U11827 ( .A1(MEM_stage_inst_dmem_n112), .A2(MEM_stage_inst_dmem_n14834), .ZN(MEM_stage_inst_dmem_n14819) );
NAND2_X1 MEM_stage_inst_dmem_U11826 ( .A1(MEM_stage_inst_dmem_ram_535), .A2(MEM_stage_inst_dmem_n14833), .ZN(MEM_stage_inst_dmem_n14820) );
NAND2_X1 MEM_stage_inst_dmem_U11825 ( .A1(MEM_stage_inst_dmem_n14818), .A2(MEM_stage_inst_dmem_n14817), .ZN(MEM_stage_inst_dmem_n11859) );
NAND2_X1 MEM_stage_inst_dmem_U11824 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n14834), .ZN(MEM_stage_inst_dmem_n14817) );
NAND2_X1 MEM_stage_inst_dmem_U11823 ( .A1(MEM_stage_inst_dmem_ram_536), .A2(MEM_stage_inst_dmem_n14833), .ZN(MEM_stage_inst_dmem_n14818) );
NAND2_X1 MEM_stage_inst_dmem_U11822 ( .A1(MEM_stage_inst_dmem_n14816), .A2(MEM_stage_inst_dmem_n14815), .ZN(MEM_stage_inst_dmem_n11860) );
NAND2_X1 MEM_stage_inst_dmem_U11821 ( .A1(MEM_stage_inst_dmem_n19251), .A2(MEM_stage_inst_dmem_n14834), .ZN(MEM_stage_inst_dmem_n14815) );
NAND2_X1 MEM_stage_inst_dmem_U11820 ( .A1(MEM_stage_inst_dmem_ram_537), .A2(MEM_stage_inst_dmem_n14833), .ZN(MEM_stage_inst_dmem_n14816) );
NAND2_X1 MEM_stage_inst_dmem_U11819 ( .A1(MEM_stage_inst_dmem_n14814), .A2(MEM_stage_inst_dmem_n14813), .ZN(MEM_stage_inst_dmem_n11861) );
NAND2_X1 MEM_stage_inst_dmem_U11818 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n14834), .ZN(MEM_stage_inst_dmem_n14813) );
NAND2_X1 MEM_stage_inst_dmem_U11817 ( .A1(MEM_stage_inst_dmem_ram_538), .A2(MEM_stage_inst_dmem_n14833), .ZN(MEM_stage_inst_dmem_n14814) );
NAND2_X1 MEM_stage_inst_dmem_U11816 ( .A1(MEM_stage_inst_dmem_n14812), .A2(MEM_stage_inst_dmem_n14811), .ZN(MEM_stage_inst_dmem_n11862) );
NAND2_X1 MEM_stage_inst_dmem_U11815 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n14834), .ZN(MEM_stage_inst_dmem_n14811) );
NAND2_X1 MEM_stage_inst_dmem_U11814 ( .A1(MEM_stage_inst_dmem_ram_539), .A2(MEM_stage_inst_dmem_n14833), .ZN(MEM_stage_inst_dmem_n14812) );
NAND2_X1 MEM_stage_inst_dmem_U11813 ( .A1(MEM_stage_inst_dmem_n14810), .A2(MEM_stage_inst_dmem_n14809), .ZN(MEM_stage_inst_dmem_n11863) );
NAND2_X1 MEM_stage_inst_dmem_U11812 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n14834), .ZN(MEM_stage_inst_dmem_n14809) );
NAND2_X1 MEM_stage_inst_dmem_U11811 ( .A1(MEM_stage_inst_dmem_ram_540), .A2(MEM_stage_inst_dmem_n14833), .ZN(MEM_stage_inst_dmem_n14810) );
NAND2_X1 MEM_stage_inst_dmem_U11810 ( .A1(MEM_stage_inst_dmem_n14808), .A2(MEM_stage_inst_dmem_n14807), .ZN(MEM_stage_inst_dmem_n11864) );
NAND2_X1 MEM_stage_inst_dmem_U11809 ( .A1(MEM_stage_inst_dmem_n15116), .A2(MEM_stage_inst_dmem_n14834), .ZN(MEM_stage_inst_dmem_n14807) );
NAND2_X1 MEM_stage_inst_dmem_U11808 ( .A1(MEM_stage_inst_dmem_ram_541), .A2(MEM_stage_inst_dmem_n14833), .ZN(MEM_stage_inst_dmem_n14808) );
NAND2_X1 MEM_stage_inst_dmem_U11807 ( .A1(MEM_stage_inst_dmem_n14806), .A2(MEM_stage_inst_dmem_n14805), .ZN(MEM_stage_inst_dmem_n11865) );
NAND2_X1 MEM_stage_inst_dmem_U11806 ( .A1(MEM_stage_inst_dmem_n15113), .A2(MEM_stage_inst_dmem_n14834), .ZN(MEM_stage_inst_dmem_n14805) );
NAND2_X1 MEM_stage_inst_dmem_U11805 ( .A1(MEM_stage_inst_dmem_ram_542), .A2(MEM_stage_inst_dmem_n14833), .ZN(MEM_stage_inst_dmem_n14806) );
NAND2_X1 MEM_stage_inst_dmem_U11804 ( .A1(MEM_stage_inst_dmem_n14804), .A2(MEM_stage_inst_dmem_n14803), .ZN(MEM_stage_inst_dmem_n11866) );
NAND2_X1 MEM_stage_inst_dmem_U11803 ( .A1(MEM_stage_inst_dmem_n16343), .A2(MEM_stage_inst_dmem_n14834), .ZN(MEM_stage_inst_dmem_n14803) );
INV_X1 MEM_stage_inst_dmem_U11802 ( .A(MEM_stage_inst_dmem_n14833), .ZN(MEM_stage_inst_dmem_n14834) );
NAND2_X1 MEM_stage_inst_dmem_U11801 ( .A1(MEM_stage_inst_dmem_ram_543), .A2(MEM_stage_inst_dmem_n14833), .ZN(MEM_stage_inst_dmem_n14804) );
NAND2_X1 MEM_stage_inst_dmem_U11800 ( .A1(MEM_stage_inst_dmem_n21429), .A2(MEM_stage_inst_dmem_n14837), .ZN(MEM_stage_inst_dmem_n14833) );
NAND2_X1 MEM_stage_inst_dmem_U11799 ( .A1(MEM_stage_inst_dmem_n14802), .A2(MEM_stage_inst_dmem_n14801), .ZN(MEM_stage_inst_dmem_n11867) );
NAND2_X1 MEM_stage_inst_dmem_U11798 ( .A1(MEM_stage_inst_dmem_n15145), .A2(MEM_stage_inst_dmem_n14800), .ZN(MEM_stage_inst_dmem_n14801) );
NAND2_X1 MEM_stage_inst_dmem_U11797 ( .A1(MEM_stage_inst_dmem_ram_544), .A2(MEM_stage_inst_dmem_n14799), .ZN(MEM_stage_inst_dmem_n14802) );
NAND2_X1 MEM_stage_inst_dmem_U11796 ( .A1(MEM_stage_inst_dmem_n14798), .A2(MEM_stage_inst_dmem_n14797), .ZN(MEM_stage_inst_dmem_n11868) );
NAND2_X1 MEM_stage_inst_dmem_U11795 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n14800), .ZN(MEM_stage_inst_dmem_n14797) );
NAND2_X1 MEM_stage_inst_dmem_U11794 ( .A1(MEM_stage_inst_dmem_ram_545), .A2(MEM_stage_inst_dmem_n14799), .ZN(MEM_stage_inst_dmem_n14798) );
NAND2_X1 MEM_stage_inst_dmem_U11793 ( .A1(MEM_stage_inst_dmem_n14796), .A2(MEM_stage_inst_dmem_n14795), .ZN(MEM_stage_inst_dmem_n11869) );
NAND2_X1 MEM_stage_inst_dmem_U11792 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n14800), .ZN(MEM_stage_inst_dmem_n14795) );
NAND2_X1 MEM_stage_inst_dmem_U11791 ( .A1(MEM_stage_inst_dmem_ram_546), .A2(MEM_stage_inst_dmem_n14799), .ZN(MEM_stage_inst_dmem_n14796) );
NAND2_X1 MEM_stage_inst_dmem_U11790 ( .A1(MEM_stage_inst_dmem_n14794), .A2(MEM_stage_inst_dmem_n14793), .ZN(MEM_stage_inst_dmem_n11870) );
NAND2_X1 MEM_stage_inst_dmem_U11789 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n14800), .ZN(MEM_stage_inst_dmem_n14793) );
NAND2_X1 MEM_stage_inst_dmem_U11788 ( .A1(MEM_stage_inst_dmem_ram_547), .A2(MEM_stage_inst_dmem_n14799), .ZN(MEM_stage_inst_dmem_n14794) );
NAND2_X1 MEM_stage_inst_dmem_U11787 ( .A1(MEM_stage_inst_dmem_n14792), .A2(MEM_stage_inst_dmem_n14791), .ZN(MEM_stage_inst_dmem_n11871) );
NAND2_X1 MEM_stage_inst_dmem_U11786 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n14800), .ZN(MEM_stage_inst_dmem_n14791) );
NAND2_X1 MEM_stage_inst_dmem_U11785 ( .A1(MEM_stage_inst_dmem_ram_548), .A2(MEM_stage_inst_dmem_n14799), .ZN(MEM_stage_inst_dmem_n14792) );
NAND2_X1 MEM_stage_inst_dmem_U11784 ( .A1(MEM_stage_inst_dmem_n14790), .A2(MEM_stage_inst_dmem_n14789), .ZN(MEM_stage_inst_dmem_n11872) );
NAND2_X1 MEM_stage_inst_dmem_U11783 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n14800), .ZN(MEM_stage_inst_dmem_n14789) );
NAND2_X1 MEM_stage_inst_dmem_U11782 ( .A1(MEM_stage_inst_dmem_ram_549), .A2(MEM_stage_inst_dmem_n14799), .ZN(MEM_stage_inst_dmem_n14790) );
NAND2_X1 MEM_stage_inst_dmem_U11781 ( .A1(MEM_stage_inst_dmem_n14788), .A2(MEM_stage_inst_dmem_n14787), .ZN(MEM_stage_inst_dmem_n11873) );
NAND2_X1 MEM_stage_inst_dmem_U11780 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n14800), .ZN(MEM_stage_inst_dmem_n14787) );
NAND2_X1 MEM_stage_inst_dmem_U11779 ( .A1(MEM_stage_inst_dmem_ram_550), .A2(MEM_stage_inst_dmem_n14799), .ZN(MEM_stage_inst_dmem_n14788) );
NAND2_X1 MEM_stage_inst_dmem_U11778 ( .A1(MEM_stage_inst_dmem_n14786), .A2(MEM_stage_inst_dmem_n14785), .ZN(MEM_stage_inst_dmem_n11874) );
NAND2_X1 MEM_stage_inst_dmem_U11777 ( .A1(MEM_stage_inst_dmem_n16361), .A2(MEM_stage_inst_dmem_n14800), .ZN(MEM_stage_inst_dmem_n14785) );
NAND2_X1 MEM_stage_inst_dmem_U11776 ( .A1(MEM_stage_inst_dmem_ram_551), .A2(MEM_stage_inst_dmem_n14799), .ZN(MEM_stage_inst_dmem_n14786) );
NAND2_X1 MEM_stage_inst_dmem_U11775 ( .A1(MEM_stage_inst_dmem_n14784), .A2(MEM_stage_inst_dmem_n14783), .ZN(MEM_stage_inst_dmem_n11875) );
NAND2_X1 MEM_stage_inst_dmem_U11774 ( .A1(MEM_stage_inst_dmem_n20527), .A2(MEM_stage_inst_dmem_n14800), .ZN(MEM_stage_inst_dmem_n14783) );
NAND2_X1 MEM_stage_inst_dmem_U11773 ( .A1(MEM_stage_inst_dmem_ram_552), .A2(MEM_stage_inst_dmem_n14799), .ZN(MEM_stage_inst_dmem_n14784) );
NAND2_X1 MEM_stage_inst_dmem_U11772 ( .A1(MEM_stage_inst_dmem_n14782), .A2(MEM_stage_inst_dmem_n14781), .ZN(MEM_stage_inst_dmem_n11876) );
NAND2_X1 MEM_stage_inst_dmem_U11771 ( .A1(MEM_stage_inst_dmem_n19251), .A2(MEM_stage_inst_dmem_n14800), .ZN(MEM_stage_inst_dmem_n14781) );
NAND2_X1 MEM_stage_inst_dmem_U11770 ( .A1(MEM_stage_inst_dmem_ram_553), .A2(MEM_stage_inst_dmem_n14799), .ZN(MEM_stage_inst_dmem_n14782) );
NAND2_X1 MEM_stage_inst_dmem_U11769 ( .A1(MEM_stage_inst_dmem_n14780), .A2(MEM_stage_inst_dmem_n14779), .ZN(MEM_stage_inst_dmem_n11877) );
NAND2_X1 MEM_stage_inst_dmem_U11768 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n14800), .ZN(MEM_stage_inst_dmem_n14779) );
NAND2_X1 MEM_stage_inst_dmem_U11767 ( .A1(MEM_stage_inst_dmem_ram_554), .A2(MEM_stage_inst_dmem_n14799), .ZN(MEM_stage_inst_dmem_n14780) );
NAND2_X1 MEM_stage_inst_dmem_U11766 ( .A1(MEM_stage_inst_dmem_n14778), .A2(MEM_stage_inst_dmem_n14777), .ZN(MEM_stage_inst_dmem_n11878) );
NAND2_X1 MEM_stage_inst_dmem_U11765 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n14800), .ZN(MEM_stage_inst_dmem_n14777) );
NAND2_X1 MEM_stage_inst_dmem_U11764 ( .A1(MEM_stage_inst_dmem_ram_555), .A2(MEM_stage_inst_dmem_n14799), .ZN(MEM_stage_inst_dmem_n14778) );
NAND2_X1 MEM_stage_inst_dmem_U11763 ( .A1(MEM_stage_inst_dmem_n14776), .A2(MEM_stage_inst_dmem_n14775), .ZN(MEM_stage_inst_dmem_n11879) );
NAND2_X1 MEM_stage_inst_dmem_U11762 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n14800), .ZN(MEM_stage_inst_dmem_n14775) );
NAND2_X1 MEM_stage_inst_dmem_U11761 ( .A1(MEM_stage_inst_dmem_ram_556), .A2(MEM_stage_inst_dmem_n14799), .ZN(MEM_stage_inst_dmem_n14776) );
NAND2_X1 MEM_stage_inst_dmem_U11760 ( .A1(MEM_stage_inst_dmem_n14774), .A2(MEM_stage_inst_dmem_n14773), .ZN(MEM_stage_inst_dmem_n11880) );
NAND2_X1 MEM_stage_inst_dmem_U11759 ( .A1(MEM_stage_inst_dmem_n15116), .A2(MEM_stage_inst_dmem_n14800), .ZN(MEM_stage_inst_dmem_n14773) );
NAND2_X1 MEM_stage_inst_dmem_U11758 ( .A1(MEM_stage_inst_dmem_ram_557), .A2(MEM_stage_inst_dmem_n14799), .ZN(MEM_stage_inst_dmem_n14774) );
NAND2_X1 MEM_stage_inst_dmem_U11757 ( .A1(MEM_stage_inst_dmem_n14772), .A2(MEM_stage_inst_dmem_n14771), .ZN(MEM_stage_inst_dmem_n11881) );
NAND2_X1 MEM_stage_inst_dmem_U11756 ( .A1(MEM_stage_inst_dmem_n15113), .A2(MEM_stage_inst_dmem_n14800), .ZN(MEM_stage_inst_dmem_n14771) );
NAND2_X1 MEM_stage_inst_dmem_U11755 ( .A1(MEM_stage_inst_dmem_ram_558), .A2(MEM_stage_inst_dmem_n14799), .ZN(MEM_stage_inst_dmem_n14772) );
NAND2_X1 MEM_stage_inst_dmem_U11754 ( .A1(MEM_stage_inst_dmem_n14770), .A2(MEM_stage_inst_dmem_n14769), .ZN(MEM_stage_inst_dmem_n11882) );
NAND2_X1 MEM_stage_inst_dmem_U11753 ( .A1(MEM_stage_inst_dmem_n14693), .A2(MEM_stage_inst_dmem_n14800), .ZN(MEM_stage_inst_dmem_n14769) );
INV_X1 MEM_stage_inst_dmem_U11752 ( .A(MEM_stage_inst_dmem_n14799), .ZN(MEM_stage_inst_dmem_n14800) );
NAND2_X1 MEM_stage_inst_dmem_U11751 ( .A1(MEM_stage_inst_dmem_ram_559), .A2(MEM_stage_inst_dmem_n14799), .ZN(MEM_stage_inst_dmem_n14770) );
NAND2_X1 MEM_stage_inst_dmem_U11750 ( .A1(MEM_stage_inst_dmem_n21394), .A2(MEM_stage_inst_dmem_n14837), .ZN(MEM_stage_inst_dmem_n14799) );
NAND2_X1 MEM_stage_inst_dmem_U11749 ( .A1(MEM_stage_inst_dmem_n14768), .A2(MEM_stage_inst_dmem_n14767), .ZN(MEM_stage_inst_dmem_n11883) );
NAND2_X1 MEM_stage_inst_dmem_U11748 ( .A1(MEM_stage_inst_dmem_n15145), .A2(MEM_stage_inst_dmem_n14766), .ZN(MEM_stage_inst_dmem_n14767) );
NAND2_X1 MEM_stage_inst_dmem_U11747 ( .A1(MEM_stage_inst_dmem_ram_560), .A2(MEM_stage_inst_dmem_n14765), .ZN(MEM_stage_inst_dmem_n14768) );
NAND2_X1 MEM_stage_inst_dmem_U11746 ( .A1(MEM_stage_inst_dmem_n14764), .A2(MEM_stage_inst_dmem_n14763), .ZN(MEM_stage_inst_dmem_n11884) );
NAND2_X1 MEM_stage_inst_dmem_U11745 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n14766), .ZN(MEM_stage_inst_dmem_n14763) );
NAND2_X1 MEM_stage_inst_dmem_U11744 ( .A1(MEM_stage_inst_dmem_ram_561), .A2(MEM_stage_inst_dmem_n14765), .ZN(MEM_stage_inst_dmem_n14764) );
NAND2_X1 MEM_stage_inst_dmem_U11743 ( .A1(MEM_stage_inst_dmem_n14762), .A2(MEM_stage_inst_dmem_n14761), .ZN(MEM_stage_inst_dmem_n11885) );
NAND2_X1 MEM_stage_inst_dmem_U11742 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n14766), .ZN(MEM_stage_inst_dmem_n14761) );
NAND2_X1 MEM_stage_inst_dmem_U11741 ( .A1(MEM_stage_inst_dmem_ram_562), .A2(MEM_stage_inst_dmem_n14765), .ZN(MEM_stage_inst_dmem_n14762) );
NAND2_X1 MEM_stage_inst_dmem_U11740 ( .A1(MEM_stage_inst_dmem_n14760), .A2(MEM_stage_inst_dmem_n14759), .ZN(MEM_stage_inst_dmem_n11886) );
NAND2_X1 MEM_stage_inst_dmem_U11739 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n14766), .ZN(MEM_stage_inst_dmem_n14759) );
NAND2_X1 MEM_stage_inst_dmem_U11738 ( .A1(MEM_stage_inst_dmem_ram_563), .A2(MEM_stage_inst_dmem_n14765), .ZN(MEM_stage_inst_dmem_n14760) );
NAND2_X1 MEM_stage_inst_dmem_U11737 ( .A1(MEM_stage_inst_dmem_n14758), .A2(MEM_stage_inst_dmem_n14757), .ZN(MEM_stage_inst_dmem_n11887) );
NAND2_X1 MEM_stage_inst_dmem_U11736 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n14766), .ZN(MEM_stage_inst_dmem_n14757) );
NAND2_X1 MEM_stage_inst_dmem_U11735 ( .A1(MEM_stage_inst_dmem_ram_564), .A2(MEM_stage_inst_dmem_n14765), .ZN(MEM_stage_inst_dmem_n14758) );
NAND2_X1 MEM_stage_inst_dmem_U11734 ( .A1(MEM_stage_inst_dmem_n14756), .A2(MEM_stage_inst_dmem_n14755), .ZN(MEM_stage_inst_dmem_n11888) );
NAND2_X1 MEM_stage_inst_dmem_U11733 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n14766), .ZN(MEM_stage_inst_dmem_n14755) );
NAND2_X1 MEM_stage_inst_dmem_U11732 ( .A1(MEM_stage_inst_dmem_ram_565), .A2(MEM_stage_inst_dmem_n14765), .ZN(MEM_stage_inst_dmem_n14756) );
NAND2_X1 MEM_stage_inst_dmem_U11731 ( .A1(MEM_stage_inst_dmem_n14754), .A2(MEM_stage_inst_dmem_n14753), .ZN(MEM_stage_inst_dmem_n11889) );
NAND2_X1 MEM_stage_inst_dmem_U11730 ( .A1(MEM_stage_inst_dmem_n20533), .A2(MEM_stage_inst_dmem_n14766), .ZN(MEM_stage_inst_dmem_n14753) );
NAND2_X1 MEM_stage_inst_dmem_U11729 ( .A1(MEM_stage_inst_dmem_ram_566), .A2(MEM_stage_inst_dmem_n14765), .ZN(MEM_stage_inst_dmem_n14754) );
NAND2_X1 MEM_stage_inst_dmem_U11728 ( .A1(MEM_stage_inst_dmem_n14752), .A2(MEM_stage_inst_dmem_n14751), .ZN(MEM_stage_inst_dmem_n11890) );
NAND2_X1 MEM_stage_inst_dmem_U11727 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n14766), .ZN(MEM_stage_inst_dmem_n14751) );
NAND2_X1 MEM_stage_inst_dmem_U11726 ( .A1(MEM_stage_inst_dmem_ram_567), .A2(MEM_stage_inst_dmem_n14765), .ZN(MEM_stage_inst_dmem_n14752) );
NAND2_X1 MEM_stage_inst_dmem_U11725 ( .A1(MEM_stage_inst_dmem_n14750), .A2(MEM_stage_inst_dmem_n14749), .ZN(MEM_stage_inst_dmem_n11891) );
NAND2_X1 MEM_stage_inst_dmem_U11724 ( .A1(MEM_stage_inst_dmem_n13883), .A2(MEM_stage_inst_dmem_n14766), .ZN(MEM_stage_inst_dmem_n14749) );
NAND2_X1 MEM_stage_inst_dmem_U11723 ( .A1(MEM_stage_inst_dmem_ram_568), .A2(MEM_stage_inst_dmem_n14765), .ZN(MEM_stage_inst_dmem_n14750) );
NAND2_X1 MEM_stage_inst_dmem_U11722 ( .A1(MEM_stage_inst_dmem_n14748), .A2(MEM_stage_inst_dmem_n14747), .ZN(MEM_stage_inst_dmem_n11892) );
NAND2_X1 MEM_stage_inst_dmem_U11721 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n14766), .ZN(MEM_stage_inst_dmem_n14747) );
NAND2_X1 MEM_stage_inst_dmem_U11720 ( .A1(MEM_stage_inst_dmem_ram_569), .A2(MEM_stage_inst_dmem_n14765), .ZN(MEM_stage_inst_dmem_n14748) );
NAND2_X1 MEM_stage_inst_dmem_U11719 ( .A1(MEM_stage_inst_dmem_n14746), .A2(MEM_stage_inst_dmem_n14745), .ZN(MEM_stage_inst_dmem_n11893) );
NAND2_X1 MEM_stage_inst_dmem_U11718 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n14766), .ZN(MEM_stage_inst_dmem_n14745) );
NAND2_X1 MEM_stage_inst_dmem_U11717 ( .A1(MEM_stage_inst_dmem_ram_570), .A2(MEM_stage_inst_dmem_n14765), .ZN(MEM_stage_inst_dmem_n14746) );
NAND2_X1 MEM_stage_inst_dmem_U11716 ( .A1(MEM_stage_inst_dmem_n14744), .A2(MEM_stage_inst_dmem_n14743), .ZN(MEM_stage_inst_dmem_n11894) );
NAND2_X1 MEM_stage_inst_dmem_U11715 ( .A1(MEM_stage_inst_dmem_n20904), .A2(MEM_stage_inst_dmem_n14766), .ZN(MEM_stage_inst_dmem_n14743) );
NAND2_X1 MEM_stage_inst_dmem_U11714 ( .A1(MEM_stage_inst_dmem_ram_571), .A2(MEM_stage_inst_dmem_n14765), .ZN(MEM_stage_inst_dmem_n14744) );
NAND2_X1 MEM_stage_inst_dmem_U11713 ( .A1(MEM_stage_inst_dmem_n14742), .A2(MEM_stage_inst_dmem_n14741), .ZN(MEM_stage_inst_dmem_n11895) );
NAND2_X1 MEM_stage_inst_dmem_U11712 ( .A1(MEM_stage_inst_dmem_n21474), .A2(MEM_stage_inst_dmem_n14766), .ZN(MEM_stage_inst_dmem_n14741) );
NAND2_X1 MEM_stage_inst_dmem_U11711 ( .A1(MEM_stage_inst_dmem_ram_572), .A2(MEM_stage_inst_dmem_n14765), .ZN(MEM_stage_inst_dmem_n14742) );
NAND2_X1 MEM_stage_inst_dmem_U11710 ( .A1(MEM_stage_inst_dmem_n14740), .A2(MEM_stage_inst_dmem_n14739), .ZN(MEM_stage_inst_dmem_n11896) );
NAND2_X1 MEM_stage_inst_dmem_U11709 ( .A1(MEM_stage_inst_dmem_n15116), .A2(MEM_stage_inst_dmem_n14766), .ZN(MEM_stage_inst_dmem_n14739) );
NAND2_X1 MEM_stage_inst_dmem_U11708 ( .A1(MEM_stage_inst_dmem_ram_573), .A2(MEM_stage_inst_dmem_n14765), .ZN(MEM_stage_inst_dmem_n14740) );
NAND2_X1 MEM_stage_inst_dmem_U11707 ( .A1(MEM_stage_inst_dmem_n14738), .A2(MEM_stage_inst_dmem_n14737), .ZN(MEM_stage_inst_dmem_n11897) );
NAND2_X1 MEM_stage_inst_dmem_U11706 ( .A1(MEM_stage_inst_dmem_n15113), .A2(MEM_stage_inst_dmem_n14766), .ZN(MEM_stage_inst_dmem_n14737) );
NAND2_X1 MEM_stage_inst_dmem_U11705 ( .A1(MEM_stage_inst_dmem_ram_574), .A2(MEM_stage_inst_dmem_n14765), .ZN(MEM_stage_inst_dmem_n14738) );
NAND2_X1 MEM_stage_inst_dmem_U11704 ( .A1(MEM_stage_inst_dmem_n14736), .A2(MEM_stage_inst_dmem_n14735), .ZN(MEM_stage_inst_dmem_n11898) );
NAND2_X1 MEM_stage_inst_dmem_U11703 ( .A1(MEM_stage_inst_dmem_n15110), .A2(MEM_stage_inst_dmem_n14766), .ZN(MEM_stage_inst_dmem_n14735) );
INV_X1 MEM_stage_inst_dmem_U11702 ( .A(MEM_stage_inst_dmem_n14765), .ZN(MEM_stage_inst_dmem_n14766) );
NAND2_X1 MEM_stage_inst_dmem_U11701 ( .A1(MEM_stage_inst_dmem_ram_575), .A2(MEM_stage_inst_dmem_n14765), .ZN(MEM_stage_inst_dmem_n14736) );
NAND2_X1 MEM_stage_inst_dmem_U11700 ( .A1(MEM_stage_inst_dmem_n21359), .A2(MEM_stage_inst_dmem_n14837), .ZN(MEM_stage_inst_dmem_n14765) );
NAND2_X1 MEM_stage_inst_dmem_U11699 ( .A1(MEM_stage_inst_dmem_n14734), .A2(MEM_stage_inst_dmem_n14733), .ZN(MEM_stage_inst_dmem_n11899) );
NAND2_X1 MEM_stage_inst_dmem_U11698 ( .A1(MEM_stage_inst_dmem_n14732), .A2(MEM_stage_inst_dmem_n14731), .ZN(MEM_stage_inst_dmem_n14733) );
NAND2_X1 MEM_stage_inst_dmem_U11697 ( .A1(MEM_stage_inst_dmem_ram_576), .A2(MEM_stage_inst_dmem_n14730), .ZN(MEM_stage_inst_dmem_n14734) );
NAND2_X1 MEM_stage_inst_dmem_U11696 ( .A1(MEM_stage_inst_dmem_n14729), .A2(MEM_stage_inst_dmem_n14728), .ZN(MEM_stage_inst_dmem_n11900) );
NAND2_X1 MEM_stage_inst_dmem_U11695 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n14731), .ZN(MEM_stage_inst_dmem_n14728) );
NAND2_X1 MEM_stage_inst_dmem_U11694 ( .A1(MEM_stage_inst_dmem_ram_577), .A2(MEM_stage_inst_dmem_n14730), .ZN(MEM_stage_inst_dmem_n14729) );
NAND2_X1 MEM_stage_inst_dmem_U11693 ( .A1(MEM_stage_inst_dmem_n14727), .A2(MEM_stage_inst_dmem_n14726), .ZN(MEM_stage_inst_dmem_n11901) );
NAND2_X1 MEM_stage_inst_dmem_U11692 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n14731), .ZN(MEM_stage_inst_dmem_n14726) );
NAND2_X1 MEM_stage_inst_dmem_U11691 ( .A1(MEM_stage_inst_dmem_ram_578), .A2(MEM_stage_inst_dmem_n14730), .ZN(MEM_stage_inst_dmem_n14727) );
NAND2_X1 MEM_stage_inst_dmem_U11690 ( .A1(MEM_stage_inst_dmem_n14725), .A2(MEM_stage_inst_dmem_n14724), .ZN(MEM_stage_inst_dmem_n11902) );
NAND2_X1 MEM_stage_inst_dmem_U11689 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n14731), .ZN(MEM_stage_inst_dmem_n14724) );
NAND2_X1 MEM_stage_inst_dmem_U11688 ( .A1(MEM_stage_inst_dmem_ram_579), .A2(MEM_stage_inst_dmem_n14730), .ZN(MEM_stage_inst_dmem_n14725) );
NAND2_X1 MEM_stage_inst_dmem_U11687 ( .A1(MEM_stage_inst_dmem_n14723), .A2(MEM_stage_inst_dmem_n14722), .ZN(MEM_stage_inst_dmem_n11903) );
NAND2_X1 MEM_stage_inst_dmem_U11686 ( .A1(MEM_stage_inst_dmem_n16368), .A2(MEM_stage_inst_dmem_n14731), .ZN(MEM_stage_inst_dmem_n14722) );
NAND2_X1 MEM_stage_inst_dmem_U11685 ( .A1(MEM_stage_inst_dmem_ram_580), .A2(MEM_stage_inst_dmem_n14730), .ZN(MEM_stage_inst_dmem_n14723) );
NAND2_X1 MEM_stage_inst_dmem_U11684 ( .A1(MEM_stage_inst_dmem_n14721), .A2(MEM_stage_inst_dmem_n14720), .ZN(MEM_stage_inst_dmem_n11904) );
NAND2_X1 MEM_stage_inst_dmem_U11683 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n14731), .ZN(MEM_stage_inst_dmem_n14720) );
NAND2_X1 MEM_stage_inst_dmem_U11682 ( .A1(MEM_stage_inst_dmem_ram_581), .A2(MEM_stage_inst_dmem_n14730), .ZN(MEM_stage_inst_dmem_n14721) );
NAND2_X1 MEM_stage_inst_dmem_U11681 ( .A1(MEM_stage_inst_dmem_n14719), .A2(MEM_stage_inst_dmem_n14718), .ZN(MEM_stage_inst_dmem_n11905) );
NAND2_X1 MEM_stage_inst_dmem_U11680 ( .A1(MEM_stage_inst_dmem_n14717), .A2(MEM_stage_inst_dmem_n14731), .ZN(MEM_stage_inst_dmem_n14718) );
NAND2_X1 MEM_stage_inst_dmem_U11679 ( .A1(MEM_stage_inst_dmem_ram_582), .A2(MEM_stage_inst_dmem_n14730), .ZN(MEM_stage_inst_dmem_n14719) );
NAND2_X1 MEM_stage_inst_dmem_U11678 ( .A1(MEM_stage_inst_dmem_n14716), .A2(MEM_stage_inst_dmem_n14715), .ZN(MEM_stage_inst_dmem_n11906) );
NAND2_X1 MEM_stage_inst_dmem_U11677 ( .A1(MEM_stage_inst_dmem_n16777), .A2(MEM_stage_inst_dmem_n14731), .ZN(MEM_stage_inst_dmem_n14715) );
NAND2_X1 MEM_stage_inst_dmem_U11676 ( .A1(MEM_stage_inst_dmem_ram_583), .A2(MEM_stage_inst_dmem_n14730), .ZN(MEM_stage_inst_dmem_n14716) );
NAND2_X1 MEM_stage_inst_dmem_U11675 ( .A1(MEM_stage_inst_dmem_n14713), .A2(MEM_stage_inst_dmem_n14712), .ZN(MEM_stage_inst_dmem_n11907) );
NAND2_X1 MEM_stage_inst_dmem_U11674 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n14731), .ZN(MEM_stage_inst_dmem_n14712) );
NAND2_X1 MEM_stage_inst_dmem_U11673 ( .A1(MEM_stage_inst_dmem_ram_584), .A2(MEM_stage_inst_dmem_n14730), .ZN(MEM_stage_inst_dmem_n14713) );
NAND2_X1 MEM_stage_inst_dmem_U11672 ( .A1(MEM_stage_inst_dmem_n14711), .A2(MEM_stage_inst_dmem_n14710), .ZN(MEM_stage_inst_dmem_n11908) );
NAND2_X1 MEM_stage_inst_dmem_U11671 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n14731), .ZN(MEM_stage_inst_dmem_n14710) );
NAND2_X1 MEM_stage_inst_dmem_U11670 ( .A1(MEM_stage_inst_dmem_ram_585), .A2(MEM_stage_inst_dmem_n14730), .ZN(MEM_stage_inst_dmem_n14711) );
NAND2_X1 MEM_stage_inst_dmem_U11669 ( .A1(MEM_stage_inst_dmem_n14709), .A2(MEM_stage_inst_dmem_n14708), .ZN(MEM_stage_inst_dmem_n11909) );
NAND2_X1 MEM_stage_inst_dmem_U11668 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n14731), .ZN(MEM_stage_inst_dmem_n14708) );
NAND2_X1 MEM_stage_inst_dmem_U11667 ( .A1(MEM_stage_inst_dmem_ram_586), .A2(MEM_stage_inst_dmem_n14730), .ZN(MEM_stage_inst_dmem_n14709) );
NAND2_X1 MEM_stage_inst_dmem_U11666 ( .A1(MEM_stage_inst_dmem_n14707), .A2(MEM_stage_inst_dmem_n14706), .ZN(MEM_stage_inst_dmem_n11910) );
NAND2_X1 MEM_stage_inst_dmem_U11665 ( .A1(MEM_stage_inst_dmem_n20904), .A2(MEM_stage_inst_dmem_n14731), .ZN(MEM_stage_inst_dmem_n14706) );
NAND2_X1 MEM_stage_inst_dmem_U11664 ( .A1(MEM_stage_inst_dmem_ram_587), .A2(MEM_stage_inst_dmem_n14730), .ZN(MEM_stage_inst_dmem_n14707) );
NAND2_X1 MEM_stage_inst_dmem_U11663 ( .A1(MEM_stage_inst_dmem_n14704), .A2(MEM_stage_inst_dmem_n14703), .ZN(MEM_stage_inst_dmem_n11911) );
NAND2_X1 MEM_stage_inst_dmem_U11662 ( .A1(MEM_stage_inst_dmem_n21474), .A2(MEM_stage_inst_dmem_n14731), .ZN(MEM_stage_inst_dmem_n14703) );
NAND2_X1 MEM_stage_inst_dmem_U11661 ( .A1(MEM_stage_inst_dmem_ram_588), .A2(MEM_stage_inst_dmem_n14730), .ZN(MEM_stage_inst_dmem_n14704) );
NAND2_X1 MEM_stage_inst_dmem_U11660 ( .A1(MEM_stage_inst_dmem_n14701), .A2(MEM_stage_inst_dmem_n14700), .ZN(MEM_stage_inst_dmem_n11912) );
NAND2_X1 MEM_stage_inst_dmem_U11659 ( .A1(MEM_stage_inst_dmem_n116), .A2(MEM_stage_inst_dmem_n14731), .ZN(MEM_stage_inst_dmem_n14700) );
NAND2_X1 MEM_stage_inst_dmem_U11658 ( .A1(MEM_stage_inst_dmem_ram_589), .A2(MEM_stage_inst_dmem_n14730), .ZN(MEM_stage_inst_dmem_n14701) );
NAND2_X1 MEM_stage_inst_dmem_U11657 ( .A1(MEM_stage_inst_dmem_n14698), .A2(MEM_stage_inst_dmem_n14697), .ZN(MEM_stage_inst_dmem_n11913) );
NAND2_X1 MEM_stage_inst_dmem_U11656 ( .A1(MEM_stage_inst_dmem_n14696), .A2(MEM_stage_inst_dmem_n14731), .ZN(MEM_stage_inst_dmem_n14697) );
NAND2_X1 MEM_stage_inst_dmem_U11655 ( .A1(MEM_stage_inst_dmem_ram_590), .A2(MEM_stage_inst_dmem_n14730), .ZN(MEM_stage_inst_dmem_n14698) );
NAND2_X1 MEM_stage_inst_dmem_U11654 ( .A1(MEM_stage_inst_dmem_n14695), .A2(MEM_stage_inst_dmem_n14694), .ZN(MEM_stage_inst_dmem_n11914) );
NAND2_X1 MEM_stage_inst_dmem_U11653 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n14731), .ZN(MEM_stage_inst_dmem_n14694) );
INV_X1 MEM_stage_inst_dmem_U11652 ( .A(MEM_stage_inst_dmem_n14730), .ZN(MEM_stage_inst_dmem_n14731) );
NAND2_X1 MEM_stage_inst_dmem_U11651 ( .A1(MEM_stage_inst_dmem_ram_591), .A2(MEM_stage_inst_dmem_n14730), .ZN(MEM_stage_inst_dmem_n14695) );
NAND2_X1 MEM_stage_inst_dmem_U11650 ( .A1(MEM_stage_inst_dmem_n21319), .A2(MEM_stage_inst_dmem_n14837), .ZN(MEM_stage_inst_dmem_n14730) );
NAND2_X1 MEM_stage_inst_dmem_U11649 ( .A1(MEM_stage_inst_dmem_n14692), .A2(MEM_stage_inst_dmem_n14691), .ZN(MEM_stage_inst_dmem_n11915) );
NAND2_X1 MEM_stage_inst_dmem_U11648 ( .A1(MEM_stage_inst_dmem_n14732), .A2(MEM_stage_inst_dmem_n14690), .ZN(MEM_stage_inst_dmem_n14691) );
NAND2_X1 MEM_stage_inst_dmem_U11647 ( .A1(MEM_stage_inst_dmem_ram_592), .A2(MEM_stage_inst_dmem_n14689), .ZN(MEM_stage_inst_dmem_n14692) );
NAND2_X1 MEM_stage_inst_dmem_U11646 ( .A1(MEM_stage_inst_dmem_n14688), .A2(MEM_stage_inst_dmem_n14687), .ZN(MEM_stage_inst_dmem_n11916) );
NAND2_X1 MEM_stage_inst_dmem_U11645 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n14690), .ZN(MEM_stage_inst_dmem_n14687) );
NAND2_X1 MEM_stage_inst_dmem_U11644 ( .A1(MEM_stage_inst_dmem_ram_593), .A2(MEM_stage_inst_dmem_n14689), .ZN(MEM_stage_inst_dmem_n14688) );
NAND2_X1 MEM_stage_inst_dmem_U11643 ( .A1(MEM_stage_inst_dmem_n14686), .A2(MEM_stage_inst_dmem_n14685), .ZN(MEM_stage_inst_dmem_n11917) );
NAND2_X1 MEM_stage_inst_dmem_U11642 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n14690), .ZN(MEM_stage_inst_dmem_n14685) );
NAND2_X1 MEM_stage_inst_dmem_U11641 ( .A1(MEM_stage_inst_dmem_ram_594), .A2(MEM_stage_inst_dmem_n14689), .ZN(MEM_stage_inst_dmem_n14686) );
NAND2_X1 MEM_stage_inst_dmem_U11640 ( .A1(MEM_stage_inst_dmem_n14684), .A2(MEM_stage_inst_dmem_n14683), .ZN(MEM_stage_inst_dmem_n11918) );
NAND2_X1 MEM_stage_inst_dmem_U11639 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n14690), .ZN(MEM_stage_inst_dmem_n14683) );
NAND2_X1 MEM_stage_inst_dmem_U11638 ( .A1(MEM_stage_inst_dmem_ram_595), .A2(MEM_stage_inst_dmem_n14689), .ZN(MEM_stage_inst_dmem_n14684) );
NAND2_X1 MEM_stage_inst_dmem_U11637 ( .A1(MEM_stage_inst_dmem_n14682), .A2(MEM_stage_inst_dmem_n14681), .ZN(MEM_stage_inst_dmem_n11919) );
NAND2_X1 MEM_stage_inst_dmem_U11636 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n14690), .ZN(MEM_stage_inst_dmem_n14681) );
NAND2_X1 MEM_stage_inst_dmem_U11635 ( .A1(MEM_stage_inst_dmem_ram_596), .A2(MEM_stage_inst_dmem_n14689), .ZN(MEM_stage_inst_dmem_n14682) );
NAND2_X1 MEM_stage_inst_dmem_U11634 ( .A1(MEM_stage_inst_dmem_n14680), .A2(MEM_stage_inst_dmem_n14679), .ZN(MEM_stage_inst_dmem_n11920) );
NAND2_X1 MEM_stage_inst_dmem_U11633 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n14690), .ZN(MEM_stage_inst_dmem_n14679) );
NAND2_X1 MEM_stage_inst_dmem_U11632 ( .A1(MEM_stage_inst_dmem_ram_597), .A2(MEM_stage_inst_dmem_n14689), .ZN(MEM_stage_inst_dmem_n14680) );
NAND2_X1 MEM_stage_inst_dmem_U11631 ( .A1(MEM_stage_inst_dmem_n14678), .A2(MEM_stage_inst_dmem_n14677), .ZN(MEM_stage_inst_dmem_n11921) );
NAND2_X1 MEM_stage_inst_dmem_U11630 ( .A1(MEM_stage_inst_dmem_n14717), .A2(MEM_stage_inst_dmem_n14690), .ZN(MEM_stage_inst_dmem_n14677) );
NAND2_X1 MEM_stage_inst_dmem_U11629 ( .A1(MEM_stage_inst_dmem_ram_598), .A2(MEM_stage_inst_dmem_n14689), .ZN(MEM_stage_inst_dmem_n14678) );
NAND2_X1 MEM_stage_inst_dmem_U11628 ( .A1(MEM_stage_inst_dmem_n14676), .A2(MEM_stage_inst_dmem_n14675), .ZN(MEM_stage_inst_dmem_n11922) );
NAND2_X1 MEM_stage_inst_dmem_U11627 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n14690), .ZN(MEM_stage_inst_dmem_n14675) );
NAND2_X1 MEM_stage_inst_dmem_U11626 ( .A1(MEM_stage_inst_dmem_ram_599), .A2(MEM_stage_inst_dmem_n14689), .ZN(MEM_stage_inst_dmem_n14676) );
NAND2_X1 MEM_stage_inst_dmem_U11625 ( .A1(MEM_stage_inst_dmem_n14674), .A2(MEM_stage_inst_dmem_n14673), .ZN(MEM_stage_inst_dmem_n11923) );
NAND2_X1 MEM_stage_inst_dmem_U11624 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n14690), .ZN(MEM_stage_inst_dmem_n14673) );
NAND2_X1 MEM_stage_inst_dmem_U11623 ( .A1(MEM_stage_inst_dmem_ram_600), .A2(MEM_stage_inst_dmem_n14689), .ZN(MEM_stage_inst_dmem_n14674) );
NAND2_X1 MEM_stage_inst_dmem_U11622 ( .A1(MEM_stage_inst_dmem_n14672), .A2(MEM_stage_inst_dmem_n14671), .ZN(MEM_stage_inst_dmem_n11924) );
NAND2_X1 MEM_stage_inst_dmem_U11621 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n14690), .ZN(MEM_stage_inst_dmem_n14671) );
NAND2_X1 MEM_stage_inst_dmem_U11620 ( .A1(MEM_stage_inst_dmem_ram_601), .A2(MEM_stage_inst_dmem_n14689), .ZN(MEM_stage_inst_dmem_n14672) );
NAND2_X1 MEM_stage_inst_dmem_U11619 ( .A1(MEM_stage_inst_dmem_n14670), .A2(MEM_stage_inst_dmem_n14669), .ZN(MEM_stage_inst_dmem_n11925) );
NAND2_X1 MEM_stage_inst_dmem_U11618 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n14690), .ZN(MEM_stage_inst_dmem_n14669) );
NAND2_X1 MEM_stage_inst_dmem_U11617 ( .A1(MEM_stage_inst_dmem_ram_602), .A2(MEM_stage_inst_dmem_n14689), .ZN(MEM_stage_inst_dmem_n14670) );
NAND2_X1 MEM_stage_inst_dmem_U11616 ( .A1(MEM_stage_inst_dmem_n14668), .A2(MEM_stage_inst_dmem_n14667), .ZN(MEM_stage_inst_dmem_n11926) );
NAND2_X1 MEM_stage_inst_dmem_U11615 ( .A1(MEM_stage_inst_dmem_n14705), .A2(MEM_stage_inst_dmem_n14690), .ZN(MEM_stage_inst_dmem_n14667) );
NAND2_X1 MEM_stage_inst_dmem_U11614 ( .A1(MEM_stage_inst_dmem_ram_603), .A2(MEM_stage_inst_dmem_n14689), .ZN(MEM_stage_inst_dmem_n14668) );
NAND2_X1 MEM_stage_inst_dmem_U11613 ( .A1(MEM_stage_inst_dmem_n14666), .A2(MEM_stage_inst_dmem_n14665), .ZN(MEM_stage_inst_dmem_n11927) );
NAND2_X1 MEM_stage_inst_dmem_U11612 ( .A1(MEM_stage_inst_dmem_n14702), .A2(MEM_stage_inst_dmem_n14690), .ZN(MEM_stage_inst_dmem_n14665) );
NAND2_X1 MEM_stage_inst_dmem_U11611 ( .A1(MEM_stage_inst_dmem_ram_604), .A2(MEM_stage_inst_dmem_n14689), .ZN(MEM_stage_inst_dmem_n14666) );
NAND2_X1 MEM_stage_inst_dmem_U11610 ( .A1(MEM_stage_inst_dmem_n14664), .A2(MEM_stage_inst_dmem_n14663), .ZN(MEM_stage_inst_dmem_n11928) );
NAND2_X1 MEM_stage_inst_dmem_U11609 ( .A1(MEM_stage_inst_dmem_n20512), .A2(MEM_stage_inst_dmem_n14690), .ZN(MEM_stage_inst_dmem_n14663) );
NAND2_X1 MEM_stage_inst_dmem_U11608 ( .A1(MEM_stage_inst_dmem_ram_605), .A2(MEM_stage_inst_dmem_n14689), .ZN(MEM_stage_inst_dmem_n14664) );
NAND2_X1 MEM_stage_inst_dmem_U11607 ( .A1(MEM_stage_inst_dmem_n14662), .A2(MEM_stage_inst_dmem_n14661), .ZN(MEM_stage_inst_dmem_n11929) );
NAND2_X1 MEM_stage_inst_dmem_U11606 ( .A1(MEM_stage_inst_dmem_n14696), .A2(MEM_stage_inst_dmem_n14690), .ZN(MEM_stage_inst_dmem_n14661) );
NAND2_X1 MEM_stage_inst_dmem_U11605 ( .A1(MEM_stage_inst_dmem_ram_606), .A2(MEM_stage_inst_dmem_n14689), .ZN(MEM_stage_inst_dmem_n14662) );
NAND2_X1 MEM_stage_inst_dmem_U11604 ( .A1(MEM_stage_inst_dmem_n14660), .A2(MEM_stage_inst_dmem_n14659), .ZN(MEM_stage_inst_dmem_n11930) );
NAND2_X1 MEM_stage_inst_dmem_U11603 ( .A1(MEM_stage_inst_dmem_n16343), .A2(MEM_stage_inst_dmem_n14690), .ZN(MEM_stage_inst_dmem_n14659) );
NAND2_X1 MEM_stage_inst_dmem_U11602 ( .A1(MEM_stage_inst_dmem_ram_607), .A2(MEM_stage_inst_dmem_n14689), .ZN(MEM_stage_inst_dmem_n14660) );
NAND2_X1 MEM_stage_inst_dmem_U11601 ( .A1(MEM_stage_inst_dmem_n21284), .A2(MEM_stage_inst_dmem_n14837), .ZN(MEM_stage_inst_dmem_n14689) );
NAND2_X1 MEM_stage_inst_dmem_U11600 ( .A1(MEM_stage_inst_dmem_n14658), .A2(MEM_stage_inst_dmem_n14657), .ZN(MEM_stage_inst_dmem_n11931) );
NAND2_X1 MEM_stage_inst_dmem_U11599 ( .A1(MEM_stage_inst_dmem_n14732), .A2(MEM_stage_inst_dmem_n14656), .ZN(MEM_stage_inst_dmem_n14657) );
NAND2_X1 MEM_stage_inst_dmem_U11598 ( .A1(MEM_stage_inst_dmem_ram_608), .A2(MEM_stage_inst_dmem_n14655), .ZN(MEM_stage_inst_dmem_n14658) );
NAND2_X1 MEM_stage_inst_dmem_U11597 ( .A1(MEM_stage_inst_dmem_n14654), .A2(MEM_stage_inst_dmem_n14653), .ZN(MEM_stage_inst_dmem_n11932) );
NAND2_X1 MEM_stage_inst_dmem_U11596 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n14656), .ZN(MEM_stage_inst_dmem_n14653) );
NAND2_X1 MEM_stage_inst_dmem_U11595 ( .A1(MEM_stage_inst_dmem_ram_609), .A2(MEM_stage_inst_dmem_n14655), .ZN(MEM_stage_inst_dmem_n14654) );
NAND2_X1 MEM_stage_inst_dmem_U11594 ( .A1(MEM_stage_inst_dmem_n14652), .A2(MEM_stage_inst_dmem_n14651), .ZN(MEM_stage_inst_dmem_n11933) );
NAND2_X1 MEM_stage_inst_dmem_U11593 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n14656), .ZN(MEM_stage_inst_dmem_n14651) );
NAND2_X1 MEM_stage_inst_dmem_U11592 ( .A1(MEM_stage_inst_dmem_ram_610), .A2(MEM_stage_inst_dmem_n14655), .ZN(MEM_stage_inst_dmem_n14652) );
NAND2_X1 MEM_stage_inst_dmem_U11591 ( .A1(MEM_stage_inst_dmem_n14650), .A2(MEM_stage_inst_dmem_n14649), .ZN(MEM_stage_inst_dmem_n11934) );
NAND2_X1 MEM_stage_inst_dmem_U11590 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n14656), .ZN(MEM_stage_inst_dmem_n14649) );
NAND2_X1 MEM_stage_inst_dmem_U11589 ( .A1(MEM_stage_inst_dmem_ram_611), .A2(MEM_stage_inst_dmem_n14655), .ZN(MEM_stage_inst_dmem_n14650) );
NAND2_X1 MEM_stage_inst_dmem_U11588 ( .A1(MEM_stage_inst_dmem_n14648), .A2(MEM_stage_inst_dmem_n14647), .ZN(MEM_stage_inst_dmem_n11935) );
NAND2_X1 MEM_stage_inst_dmem_U11587 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n14656), .ZN(MEM_stage_inst_dmem_n14647) );
NAND2_X1 MEM_stage_inst_dmem_U11586 ( .A1(MEM_stage_inst_dmem_ram_612), .A2(MEM_stage_inst_dmem_n14655), .ZN(MEM_stage_inst_dmem_n14648) );
NAND2_X1 MEM_stage_inst_dmem_U11585 ( .A1(MEM_stage_inst_dmem_n14646), .A2(MEM_stage_inst_dmem_n14645), .ZN(MEM_stage_inst_dmem_n11936) );
NAND2_X1 MEM_stage_inst_dmem_U11584 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n14656), .ZN(MEM_stage_inst_dmem_n14645) );
NAND2_X1 MEM_stage_inst_dmem_U11583 ( .A1(MEM_stage_inst_dmem_ram_613), .A2(MEM_stage_inst_dmem_n14655), .ZN(MEM_stage_inst_dmem_n14646) );
NAND2_X1 MEM_stage_inst_dmem_U11582 ( .A1(MEM_stage_inst_dmem_n14644), .A2(MEM_stage_inst_dmem_n14643), .ZN(MEM_stage_inst_dmem_n11937) );
NAND2_X1 MEM_stage_inst_dmem_U11581 ( .A1(MEM_stage_inst_dmem_n14717), .A2(MEM_stage_inst_dmem_n14656), .ZN(MEM_stage_inst_dmem_n14643) );
NAND2_X1 MEM_stage_inst_dmem_U11580 ( .A1(MEM_stage_inst_dmem_ram_614), .A2(MEM_stage_inst_dmem_n14655), .ZN(MEM_stage_inst_dmem_n14644) );
NAND2_X1 MEM_stage_inst_dmem_U11579 ( .A1(MEM_stage_inst_dmem_n14642), .A2(MEM_stage_inst_dmem_n14641), .ZN(MEM_stage_inst_dmem_n11938) );
NAND2_X1 MEM_stage_inst_dmem_U11578 ( .A1(MEM_stage_inst_dmem_n16361), .A2(MEM_stage_inst_dmem_n14656), .ZN(MEM_stage_inst_dmem_n14641) );
NAND2_X1 MEM_stage_inst_dmem_U11577 ( .A1(MEM_stage_inst_dmem_ram_615), .A2(MEM_stage_inst_dmem_n14655), .ZN(MEM_stage_inst_dmem_n14642) );
NAND2_X1 MEM_stage_inst_dmem_U11576 ( .A1(MEM_stage_inst_dmem_n14640), .A2(MEM_stage_inst_dmem_n14639), .ZN(MEM_stage_inst_dmem_n11939) );
NAND2_X1 MEM_stage_inst_dmem_U11575 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n14656), .ZN(MEM_stage_inst_dmem_n14639) );
NAND2_X1 MEM_stage_inst_dmem_U11574 ( .A1(MEM_stage_inst_dmem_ram_616), .A2(MEM_stage_inst_dmem_n14655), .ZN(MEM_stage_inst_dmem_n14640) );
NAND2_X1 MEM_stage_inst_dmem_U11573 ( .A1(MEM_stage_inst_dmem_n14638), .A2(MEM_stage_inst_dmem_n14637), .ZN(MEM_stage_inst_dmem_n11940) );
NAND2_X1 MEM_stage_inst_dmem_U11572 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n14656), .ZN(MEM_stage_inst_dmem_n14637) );
NAND2_X1 MEM_stage_inst_dmem_U11571 ( .A1(MEM_stage_inst_dmem_ram_617), .A2(MEM_stage_inst_dmem_n14655), .ZN(MEM_stage_inst_dmem_n14638) );
NAND2_X1 MEM_stage_inst_dmem_U11570 ( .A1(MEM_stage_inst_dmem_n14636), .A2(MEM_stage_inst_dmem_n14635), .ZN(MEM_stage_inst_dmem_n11941) );
NAND2_X1 MEM_stage_inst_dmem_U11569 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n14656), .ZN(MEM_stage_inst_dmem_n14635) );
NAND2_X1 MEM_stage_inst_dmem_U11568 ( .A1(MEM_stage_inst_dmem_ram_618), .A2(MEM_stage_inst_dmem_n14655), .ZN(MEM_stage_inst_dmem_n14636) );
NAND2_X1 MEM_stage_inst_dmem_U11567 ( .A1(MEM_stage_inst_dmem_n14634), .A2(MEM_stage_inst_dmem_n14633), .ZN(MEM_stage_inst_dmem_n11942) );
NAND2_X1 MEM_stage_inst_dmem_U11566 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n14656), .ZN(MEM_stage_inst_dmem_n14633) );
NAND2_X1 MEM_stage_inst_dmem_U11565 ( .A1(MEM_stage_inst_dmem_ram_619), .A2(MEM_stage_inst_dmem_n14655), .ZN(MEM_stage_inst_dmem_n14634) );
NAND2_X1 MEM_stage_inst_dmem_U11564 ( .A1(MEM_stage_inst_dmem_n14632), .A2(MEM_stage_inst_dmem_n14631), .ZN(MEM_stage_inst_dmem_n11943) );
NAND2_X1 MEM_stage_inst_dmem_U11563 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n14656), .ZN(MEM_stage_inst_dmem_n14631) );
NAND2_X1 MEM_stage_inst_dmem_U11562 ( .A1(MEM_stage_inst_dmem_ram_620), .A2(MEM_stage_inst_dmem_n14655), .ZN(MEM_stage_inst_dmem_n14632) );
NAND2_X1 MEM_stage_inst_dmem_U11561 ( .A1(MEM_stage_inst_dmem_n14630), .A2(MEM_stage_inst_dmem_n14629), .ZN(MEM_stage_inst_dmem_n11944) );
NAND2_X1 MEM_stage_inst_dmem_U11560 ( .A1(MEM_stage_inst_dmem_n116), .A2(MEM_stage_inst_dmem_n14656), .ZN(MEM_stage_inst_dmem_n14629) );
NAND2_X1 MEM_stage_inst_dmem_U11559 ( .A1(MEM_stage_inst_dmem_ram_621), .A2(MEM_stage_inst_dmem_n14655), .ZN(MEM_stage_inst_dmem_n14630) );
NAND2_X1 MEM_stage_inst_dmem_U11558 ( .A1(MEM_stage_inst_dmem_n14628), .A2(MEM_stage_inst_dmem_n14627), .ZN(MEM_stage_inst_dmem_n11945) );
NAND2_X1 MEM_stage_inst_dmem_U11557 ( .A1(MEM_stage_inst_dmem_n14696), .A2(MEM_stage_inst_dmem_n14656), .ZN(MEM_stage_inst_dmem_n14627) );
NAND2_X1 MEM_stage_inst_dmem_U11556 ( .A1(MEM_stage_inst_dmem_ram_622), .A2(MEM_stage_inst_dmem_n14655), .ZN(MEM_stage_inst_dmem_n14628) );
NAND2_X1 MEM_stage_inst_dmem_U11555 ( .A1(MEM_stage_inst_dmem_n14626), .A2(MEM_stage_inst_dmem_n14625), .ZN(MEM_stage_inst_dmem_n11946) );
NAND2_X1 MEM_stage_inst_dmem_U11554 ( .A1(MEM_stage_inst_dmem_n14693), .A2(MEM_stage_inst_dmem_n14656), .ZN(MEM_stage_inst_dmem_n14625) );
INV_X1 MEM_stage_inst_dmem_U11553 ( .A(MEM_stage_inst_dmem_n14655), .ZN(MEM_stage_inst_dmem_n14656) );
NAND2_X1 MEM_stage_inst_dmem_U11552 ( .A1(MEM_stage_inst_dmem_ram_623), .A2(MEM_stage_inst_dmem_n14655), .ZN(MEM_stage_inst_dmem_n14626) );
NAND2_X1 MEM_stage_inst_dmem_U11551 ( .A1(MEM_stage_inst_dmem_n21249), .A2(MEM_stage_inst_dmem_n14837), .ZN(MEM_stage_inst_dmem_n14655) );
NAND2_X1 MEM_stage_inst_dmem_U11550 ( .A1(MEM_stage_inst_dmem_n14624), .A2(MEM_stage_inst_dmem_n14623), .ZN(MEM_stage_inst_dmem_n11947) );
NAND2_X1 MEM_stage_inst_dmem_U11549 ( .A1(MEM_stage_inst_dmem_n14732), .A2(MEM_stage_inst_dmem_n14622), .ZN(MEM_stage_inst_dmem_n14623) );
NAND2_X1 MEM_stage_inst_dmem_U11548 ( .A1(MEM_stage_inst_dmem_ram_624), .A2(MEM_stage_inst_dmem_n14621), .ZN(MEM_stage_inst_dmem_n14624) );
NAND2_X1 MEM_stage_inst_dmem_U11547 ( .A1(MEM_stage_inst_dmem_n14620), .A2(MEM_stage_inst_dmem_n14619), .ZN(MEM_stage_inst_dmem_n11948) );
NAND2_X1 MEM_stage_inst_dmem_U11546 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n14622), .ZN(MEM_stage_inst_dmem_n14619) );
NAND2_X1 MEM_stage_inst_dmem_U11545 ( .A1(MEM_stage_inst_dmem_ram_625), .A2(MEM_stage_inst_dmem_n14621), .ZN(MEM_stage_inst_dmem_n14620) );
NAND2_X1 MEM_stage_inst_dmem_U11544 ( .A1(MEM_stage_inst_dmem_n14618), .A2(MEM_stage_inst_dmem_n14617), .ZN(MEM_stage_inst_dmem_n11949) );
NAND2_X1 MEM_stage_inst_dmem_U11543 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n14622), .ZN(MEM_stage_inst_dmem_n14617) );
NAND2_X1 MEM_stage_inst_dmem_U11542 ( .A1(MEM_stage_inst_dmem_ram_626), .A2(MEM_stage_inst_dmem_n14621), .ZN(MEM_stage_inst_dmem_n14618) );
NAND2_X1 MEM_stage_inst_dmem_U11541 ( .A1(MEM_stage_inst_dmem_n14616), .A2(MEM_stage_inst_dmem_n14615), .ZN(MEM_stage_inst_dmem_n11950) );
NAND2_X1 MEM_stage_inst_dmem_U11540 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n14622), .ZN(MEM_stage_inst_dmem_n14615) );
NAND2_X1 MEM_stage_inst_dmem_U11539 ( .A1(MEM_stage_inst_dmem_ram_627), .A2(MEM_stage_inst_dmem_n14621), .ZN(MEM_stage_inst_dmem_n14616) );
NAND2_X1 MEM_stage_inst_dmem_U11538 ( .A1(MEM_stage_inst_dmem_n14614), .A2(MEM_stage_inst_dmem_n14613), .ZN(MEM_stage_inst_dmem_n11951) );
NAND2_X1 MEM_stage_inst_dmem_U11537 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n14622), .ZN(MEM_stage_inst_dmem_n14613) );
NAND2_X1 MEM_stage_inst_dmem_U11536 ( .A1(MEM_stage_inst_dmem_ram_628), .A2(MEM_stage_inst_dmem_n14621), .ZN(MEM_stage_inst_dmem_n14614) );
NAND2_X1 MEM_stage_inst_dmem_U11535 ( .A1(MEM_stage_inst_dmem_n14612), .A2(MEM_stage_inst_dmem_n14611), .ZN(MEM_stage_inst_dmem_n11952) );
NAND2_X1 MEM_stage_inst_dmem_U11534 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n14622), .ZN(MEM_stage_inst_dmem_n14611) );
NAND2_X1 MEM_stage_inst_dmem_U11533 ( .A1(MEM_stage_inst_dmem_ram_629), .A2(MEM_stage_inst_dmem_n14621), .ZN(MEM_stage_inst_dmem_n14612) );
NAND2_X1 MEM_stage_inst_dmem_U11532 ( .A1(MEM_stage_inst_dmem_n14610), .A2(MEM_stage_inst_dmem_n14609), .ZN(MEM_stage_inst_dmem_n11953) );
NAND2_X1 MEM_stage_inst_dmem_U11531 ( .A1(MEM_stage_inst_dmem_n14717), .A2(MEM_stage_inst_dmem_n14622), .ZN(MEM_stage_inst_dmem_n14609) );
NAND2_X1 MEM_stage_inst_dmem_U11530 ( .A1(MEM_stage_inst_dmem_ram_630), .A2(MEM_stage_inst_dmem_n14621), .ZN(MEM_stage_inst_dmem_n14610) );
NAND2_X1 MEM_stage_inst_dmem_U11529 ( .A1(MEM_stage_inst_dmem_n14608), .A2(MEM_stage_inst_dmem_n14607), .ZN(MEM_stage_inst_dmem_n11954) );
NAND2_X1 MEM_stage_inst_dmem_U11528 ( .A1(MEM_stage_inst_dmem_n20530), .A2(MEM_stage_inst_dmem_n14622), .ZN(MEM_stage_inst_dmem_n14607) );
NAND2_X1 MEM_stage_inst_dmem_U11527 ( .A1(MEM_stage_inst_dmem_ram_631), .A2(MEM_stage_inst_dmem_n14621), .ZN(MEM_stage_inst_dmem_n14608) );
NAND2_X1 MEM_stage_inst_dmem_U11526 ( .A1(MEM_stage_inst_dmem_n14606), .A2(MEM_stage_inst_dmem_n14605), .ZN(MEM_stage_inst_dmem_n11955) );
NAND2_X1 MEM_stage_inst_dmem_U11525 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n14622), .ZN(MEM_stage_inst_dmem_n14605) );
NAND2_X1 MEM_stage_inst_dmem_U11524 ( .A1(MEM_stage_inst_dmem_ram_632), .A2(MEM_stage_inst_dmem_n14621), .ZN(MEM_stage_inst_dmem_n14606) );
NAND2_X1 MEM_stage_inst_dmem_U11523 ( .A1(MEM_stage_inst_dmem_n14604), .A2(MEM_stage_inst_dmem_n14603), .ZN(MEM_stage_inst_dmem_n11956) );
NAND2_X1 MEM_stage_inst_dmem_U11522 ( .A1(MEM_stage_inst_dmem_n20524), .A2(MEM_stage_inst_dmem_n14622), .ZN(MEM_stage_inst_dmem_n14603) );
NAND2_X1 MEM_stage_inst_dmem_U11521 ( .A1(MEM_stage_inst_dmem_ram_633), .A2(MEM_stage_inst_dmem_n14621), .ZN(MEM_stage_inst_dmem_n14604) );
NAND2_X1 MEM_stage_inst_dmem_U11520 ( .A1(MEM_stage_inst_dmem_n14602), .A2(MEM_stage_inst_dmem_n14601), .ZN(MEM_stage_inst_dmem_n11957) );
NAND2_X1 MEM_stage_inst_dmem_U11519 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n14622), .ZN(MEM_stage_inst_dmem_n14601) );
NAND2_X1 MEM_stage_inst_dmem_U11518 ( .A1(MEM_stage_inst_dmem_ram_634), .A2(MEM_stage_inst_dmem_n14621), .ZN(MEM_stage_inst_dmem_n14602) );
NAND2_X1 MEM_stage_inst_dmem_U11517 ( .A1(MEM_stage_inst_dmem_n14600), .A2(MEM_stage_inst_dmem_n14599), .ZN(MEM_stage_inst_dmem_n11958) );
NAND2_X1 MEM_stage_inst_dmem_U11516 ( .A1(MEM_stage_inst_dmem_n20904), .A2(MEM_stage_inst_dmem_n14622), .ZN(MEM_stage_inst_dmem_n14599) );
NAND2_X1 MEM_stage_inst_dmem_U11515 ( .A1(MEM_stage_inst_dmem_ram_635), .A2(MEM_stage_inst_dmem_n14621), .ZN(MEM_stage_inst_dmem_n14600) );
NAND2_X1 MEM_stage_inst_dmem_U11514 ( .A1(MEM_stage_inst_dmem_n14598), .A2(MEM_stage_inst_dmem_n14597), .ZN(MEM_stage_inst_dmem_n11959) );
NAND2_X1 MEM_stage_inst_dmem_U11513 ( .A1(MEM_stage_inst_dmem_n21474), .A2(MEM_stage_inst_dmem_n14622), .ZN(MEM_stage_inst_dmem_n14597) );
NAND2_X1 MEM_stage_inst_dmem_U11512 ( .A1(MEM_stage_inst_dmem_ram_636), .A2(MEM_stage_inst_dmem_n14621), .ZN(MEM_stage_inst_dmem_n14598) );
NAND2_X1 MEM_stage_inst_dmem_U11511 ( .A1(MEM_stage_inst_dmem_n14596), .A2(MEM_stage_inst_dmem_n14595), .ZN(MEM_stage_inst_dmem_n11960) );
NAND2_X1 MEM_stage_inst_dmem_U11510 ( .A1(MEM_stage_inst_dmem_n116), .A2(MEM_stage_inst_dmem_n14622), .ZN(MEM_stage_inst_dmem_n14595) );
NAND2_X1 MEM_stage_inst_dmem_U11509 ( .A1(MEM_stage_inst_dmem_ram_637), .A2(MEM_stage_inst_dmem_n14621), .ZN(MEM_stage_inst_dmem_n14596) );
NAND2_X1 MEM_stage_inst_dmem_U11508 ( .A1(MEM_stage_inst_dmem_n14594), .A2(MEM_stage_inst_dmem_n14593), .ZN(MEM_stage_inst_dmem_n11961) );
NAND2_X1 MEM_stage_inst_dmem_U11507 ( .A1(MEM_stage_inst_dmem_n14696), .A2(MEM_stage_inst_dmem_n14622), .ZN(MEM_stage_inst_dmem_n14593) );
NAND2_X1 MEM_stage_inst_dmem_U11506 ( .A1(MEM_stage_inst_dmem_ram_638), .A2(MEM_stage_inst_dmem_n14621), .ZN(MEM_stage_inst_dmem_n14594) );
NAND2_X1 MEM_stage_inst_dmem_U11505 ( .A1(MEM_stage_inst_dmem_n14592), .A2(MEM_stage_inst_dmem_n14591), .ZN(MEM_stage_inst_dmem_n11962) );
NAND2_X1 MEM_stage_inst_dmem_U11504 ( .A1(MEM_stage_inst_dmem_n15110), .A2(MEM_stage_inst_dmem_n14622), .ZN(MEM_stage_inst_dmem_n14591) );
INV_X1 MEM_stage_inst_dmem_U11503 ( .A(MEM_stage_inst_dmem_n14621), .ZN(MEM_stage_inst_dmem_n14622) );
NAND2_X1 MEM_stage_inst_dmem_U11502 ( .A1(MEM_stage_inst_dmem_ram_639), .A2(MEM_stage_inst_dmem_n14621), .ZN(MEM_stage_inst_dmem_n14592) );
NAND2_X1 MEM_stage_inst_dmem_U11501 ( .A1(MEM_stage_inst_dmem_n21214), .A2(MEM_stage_inst_dmem_n14837), .ZN(MEM_stage_inst_dmem_n14621) );
NAND2_X1 MEM_stage_inst_dmem_U11500 ( .A1(MEM_stage_inst_dmem_n14590), .A2(MEM_stage_inst_dmem_n14589), .ZN(MEM_stage_inst_dmem_n11963) );
NAND2_X1 MEM_stage_inst_dmem_U11499 ( .A1(MEM_stage_inst_dmem_n14732), .A2(MEM_stage_inst_dmem_n14588), .ZN(MEM_stage_inst_dmem_n14589) );
NAND2_X1 MEM_stage_inst_dmem_U11498 ( .A1(MEM_stage_inst_dmem_ram_640), .A2(MEM_stage_inst_dmem_n14587), .ZN(MEM_stage_inst_dmem_n14590) );
NAND2_X1 MEM_stage_inst_dmem_U11497 ( .A1(MEM_stage_inst_dmem_n14586), .A2(MEM_stage_inst_dmem_n14585), .ZN(MEM_stage_inst_dmem_n11964) );
NAND2_X1 MEM_stage_inst_dmem_U11496 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n14588), .ZN(MEM_stage_inst_dmem_n14585) );
NAND2_X1 MEM_stage_inst_dmem_U11495 ( .A1(MEM_stage_inst_dmem_ram_641), .A2(MEM_stage_inst_dmem_n14587), .ZN(MEM_stage_inst_dmem_n14586) );
NAND2_X1 MEM_stage_inst_dmem_U11494 ( .A1(MEM_stage_inst_dmem_n14584), .A2(MEM_stage_inst_dmem_n14583), .ZN(MEM_stage_inst_dmem_n11965) );
NAND2_X1 MEM_stage_inst_dmem_U11493 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n14588), .ZN(MEM_stage_inst_dmem_n14583) );
NAND2_X1 MEM_stage_inst_dmem_U11492 ( .A1(MEM_stage_inst_dmem_ram_642), .A2(MEM_stage_inst_dmem_n14587), .ZN(MEM_stage_inst_dmem_n14584) );
NAND2_X1 MEM_stage_inst_dmem_U11491 ( .A1(MEM_stage_inst_dmem_n14582), .A2(MEM_stage_inst_dmem_n14581), .ZN(MEM_stage_inst_dmem_n11966) );
NAND2_X1 MEM_stage_inst_dmem_U11490 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n14588), .ZN(MEM_stage_inst_dmem_n14581) );
NAND2_X1 MEM_stage_inst_dmem_U11489 ( .A1(MEM_stage_inst_dmem_ram_643), .A2(MEM_stage_inst_dmem_n14587), .ZN(MEM_stage_inst_dmem_n14582) );
NAND2_X1 MEM_stage_inst_dmem_U11488 ( .A1(MEM_stage_inst_dmem_n14580), .A2(MEM_stage_inst_dmem_n14579), .ZN(MEM_stage_inst_dmem_n11967) );
NAND2_X1 MEM_stage_inst_dmem_U11487 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n14588), .ZN(MEM_stage_inst_dmem_n14579) );
NAND2_X1 MEM_stage_inst_dmem_U11486 ( .A1(MEM_stage_inst_dmem_ram_644), .A2(MEM_stage_inst_dmem_n14587), .ZN(MEM_stage_inst_dmem_n14580) );
NAND2_X1 MEM_stage_inst_dmem_U11485 ( .A1(MEM_stage_inst_dmem_n14578), .A2(MEM_stage_inst_dmem_n14577), .ZN(MEM_stage_inst_dmem_n11968) );
NAND2_X1 MEM_stage_inst_dmem_U11484 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n14588), .ZN(MEM_stage_inst_dmem_n14577) );
NAND2_X1 MEM_stage_inst_dmem_U11483 ( .A1(MEM_stage_inst_dmem_ram_645), .A2(MEM_stage_inst_dmem_n14587), .ZN(MEM_stage_inst_dmem_n14578) );
NAND2_X1 MEM_stage_inst_dmem_U11482 ( .A1(MEM_stage_inst_dmem_n14576), .A2(MEM_stage_inst_dmem_n14575), .ZN(MEM_stage_inst_dmem_n11969) );
NAND2_X1 MEM_stage_inst_dmem_U11481 ( .A1(MEM_stage_inst_dmem_n14717), .A2(MEM_stage_inst_dmem_n14588), .ZN(MEM_stage_inst_dmem_n14575) );
NAND2_X1 MEM_stage_inst_dmem_U11480 ( .A1(MEM_stage_inst_dmem_ram_646), .A2(MEM_stage_inst_dmem_n14587), .ZN(MEM_stage_inst_dmem_n14576) );
NAND2_X1 MEM_stage_inst_dmem_U11479 ( .A1(MEM_stage_inst_dmem_n14574), .A2(MEM_stage_inst_dmem_n14573), .ZN(MEM_stage_inst_dmem_n11970) );
NAND2_X1 MEM_stage_inst_dmem_U11478 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n14588), .ZN(MEM_stage_inst_dmem_n14573) );
NAND2_X1 MEM_stage_inst_dmem_U11477 ( .A1(MEM_stage_inst_dmem_ram_647), .A2(MEM_stage_inst_dmem_n14587), .ZN(MEM_stage_inst_dmem_n14574) );
NAND2_X1 MEM_stage_inst_dmem_U11476 ( .A1(MEM_stage_inst_dmem_n14572), .A2(MEM_stage_inst_dmem_n14571), .ZN(MEM_stage_inst_dmem_n11971) );
NAND2_X1 MEM_stage_inst_dmem_U11475 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n14588), .ZN(MEM_stage_inst_dmem_n14571) );
NAND2_X1 MEM_stage_inst_dmem_U11474 ( .A1(MEM_stage_inst_dmem_ram_648), .A2(MEM_stage_inst_dmem_n14587), .ZN(MEM_stage_inst_dmem_n14572) );
NAND2_X1 MEM_stage_inst_dmem_U11473 ( .A1(MEM_stage_inst_dmem_n14570), .A2(MEM_stage_inst_dmem_n14569), .ZN(MEM_stage_inst_dmem_n11972) );
NAND2_X1 MEM_stage_inst_dmem_U11472 ( .A1(MEM_stage_inst_dmem_n96), .A2(MEM_stage_inst_dmem_n14588), .ZN(MEM_stage_inst_dmem_n14569) );
NAND2_X1 MEM_stage_inst_dmem_U11471 ( .A1(MEM_stage_inst_dmem_ram_649), .A2(MEM_stage_inst_dmem_n14587), .ZN(MEM_stage_inst_dmem_n14570) );
NAND2_X1 MEM_stage_inst_dmem_U11470 ( .A1(MEM_stage_inst_dmem_n14568), .A2(MEM_stage_inst_dmem_n14567), .ZN(MEM_stage_inst_dmem_n11973) );
NAND2_X1 MEM_stage_inst_dmem_U11469 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n14588), .ZN(MEM_stage_inst_dmem_n14567) );
NAND2_X1 MEM_stage_inst_dmem_U11468 ( .A1(MEM_stage_inst_dmem_ram_650), .A2(MEM_stage_inst_dmem_n14587), .ZN(MEM_stage_inst_dmem_n14568) );
NAND2_X1 MEM_stage_inst_dmem_U11467 ( .A1(MEM_stage_inst_dmem_n14566), .A2(MEM_stage_inst_dmem_n14565), .ZN(MEM_stage_inst_dmem_n11974) );
NAND2_X1 MEM_stage_inst_dmem_U11466 ( .A1(MEM_stage_inst_dmem_n14705), .A2(MEM_stage_inst_dmem_n14588), .ZN(MEM_stage_inst_dmem_n14565) );
NAND2_X1 MEM_stage_inst_dmem_U11465 ( .A1(MEM_stage_inst_dmem_ram_651), .A2(MEM_stage_inst_dmem_n14587), .ZN(MEM_stage_inst_dmem_n14566) );
NAND2_X1 MEM_stage_inst_dmem_U11464 ( .A1(MEM_stage_inst_dmem_n14564), .A2(MEM_stage_inst_dmem_n14563), .ZN(MEM_stage_inst_dmem_n11975) );
NAND2_X1 MEM_stage_inst_dmem_U11463 ( .A1(MEM_stage_inst_dmem_n14702), .A2(MEM_stage_inst_dmem_n14588), .ZN(MEM_stage_inst_dmem_n14563) );
NAND2_X1 MEM_stage_inst_dmem_U11462 ( .A1(MEM_stage_inst_dmem_ram_652), .A2(MEM_stage_inst_dmem_n14587), .ZN(MEM_stage_inst_dmem_n14564) );
NAND2_X1 MEM_stage_inst_dmem_U11461 ( .A1(MEM_stage_inst_dmem_n14562), .A2(MEM_stage_inst_dmem_n14561), .ZN(MEM_stage_inst_dmem_n11976) );
NAND2_X1 MEM_stage_inst_dmem_U11460 ( .A1(MEM_stage_inst_dmem_n116), .A2(MEM_stage_inst_dmem_n14588), .ZN(MEM_stage_inst_dmem_n14561) );
NAND2_X1 MEM_stage_inst_dmem_U11459 ( .A1(MEM_stage_inst_dmem_ram_653), .A2(MEM_stage_inst_dmem_n14587), .ZN(MEM_stage_inst_dmem_n14562) );
NAND2_X1 MEM_stage_inst_dmem_U11458 ( .A1(MEM_stage_inst_dmem_n14560), .A2(MEM_stage_inst_dmem_n14559), .ZN(MEM_stage_inst_dmem_n11977) );
NAND2_X1 MEM_stage_inst_dmem_U11457 ( .A1(MEM_stage_inst_dmem_n14696), .A2(MEM_stage_inst_dmem_n14588), .ZN(MEM_stage_inst_dmem_n14559) );
NAND2_X1 MEM_stage_inst_dmem_U11456 ( .A1(MEM_stage_inst_dmem_ram_654), .A2(MEM_stage_inst_dmem_n14587), .ZN(MEM_stage_inst_dmem_n14560) );
NAND2_X1 MEM_stage_inst_dmem_U11455 ( .A1(MEM_stage_inst_dmem_n14558), .A2(MEM_stage_inst_dmem_n14557), .ZN(MEM_stage_inst_dmem_n11978) );
NAND2_X1 MEM_stage_inst_dmem_U11454 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n14588), .ZN(MEM_stage_inst_dmem_n14557) );
INV_X1 MEM_stage_inst_dmem_U11453 ( .A(MEM_stage_inst_dmem_n14587), .ZN(MEM_stage_inst_dmem_n14588) );
NAND2_X1 MEM_stage_inst_dmem_U11452 ( .A1(MEM_stage_inst_dmem_ram_655), .A2(MEM_stage_inst_dmem_n14587), .ZN(MEM_stage_inst_dmem_n14558) );
NAND2_X1 MEM_stage_inst_dmem_U11451 ( .A1(MEM_stage_inst_dmem_n21179), .A2(MEM_stage_inst_dmem_n14837), .ZN(MEM_stage_inst_dmem_n14587) );
NAND2_X1 MEM_stage_inst_dmem_U11450 ( .A1(MEM_stage_inst_dmem_n14556), .A2(MEM_stage_inst_dmem_n14555), .ZN(MEM_stage_inst_dmem_n11979) );
NAND2_X1 MEM_stage_inst_dmem_U11449 ( .A1(MEM_stage_inst_dmem_n14732), .A2(MEM_stage_inst_dmem_n14554), .ZN(MEM_stage_inst_dmem_n14555) );
NAND2_X1 MEM_stage_inst_dmem_U11448 ( .A1(MEM_stage_inst_dmem_ram_656), .A2(MEM_stage_inst_dmem_n14553), .ZN(MEM_stage_inst_dmem_n14556) );
NAND2_X1 MEM_stage_inst_dmem_U11447 ( .A1(MEM_stage_inst_dmem_n14552), .A2(MEM_stage_inst_dmem_n14551), .ZN(MEM_stage_inst_dmem_n11980) );
NAND2_X1 MEM_stage_inst_dmem_U11446 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n14554), .ZN(MEM_stage_inst_dmem_n14551) );
NAND2_X1 MEM_stage_inst_dmem_U11445 ( .A1(MEM_stage_inst_dmem_ram_657), .A2(MEM_stage_inst_dmem_n14553), .ZN(MEM_stage_inst_dmem_n14552) );
NAND2_X1 MEM_stage_inst_dmem_U11444 ( .A1(MEM_stage_inst_dmem_n14550), .A2(MEM_stage_inst_dmem_n14549), .ZN(MEM_stage_inst_dmem_n11981) );
NAND2_X1 MEM_stage_inst_dmem_U11443 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n14554), .ZN(MEM_stage_inst_dmem_n14549) );
NAND2_X1 MEM_stage_inst_dmem_U11442 ( .A1(MEM_stage_inst_dmem_ram_658), .A2(MEM_stage_inst_dmem_n14553), .ZN(MEM_stage_inst_dmem_n14550) );
NAND2_X1 MEM_stage_inst_dmem_U11441 ( .A1(MEM_stage_inst_dmem_n14548), .A2(MEM_stage_inst_dmem_n14547), .ZN(MEM_stage_inst_dmem_n11982) );
NAND2_X1 MEM_stage_inst_dmem_U11440 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n14554), .ZN(MEM_stage_inst_dmem_n14547) );
NAND2_X1 MEM_stage_inst_dmem_U11439 ( .A1(MEM_stage_inst_dmem_ram_659), .A2(MEM_stage_inst_dmem_n14553), .ZN(MEM_stage_inst_dmem_n14548) );
NAND2_X1 MEM_stage_inst_dmem_U11438 ( .A1(MEM_stage_inst_dmem_n14546), .A2(MEM_stage_inst_dmem_n14545), .ZN(MEM_stage_inst_dmem_n11983) );
NAND2_X1 MEM_stage_inst_dmem_U11437 ( .A1(MEM_stage_inst_dmem_n16368), .A2(MEM_stage_inst_dmem_n14554), .ZN(MEM_stage_inst_dmem_n14545) );
NAND2_X1 MEM_stage_inst_dmem_U11436 ( .A1(MEM_stage_inst_dmem_ram_660), .A2(MEM_stage_inst_dmem_n14553), .ZN(MEM_stage_inst_dmem_n14546) );
NAND2_X1 MEM_stage_inst_dmem_U11435 ( .A1(MEM_stage_inst_dmem_n14544), .A2(MEM_stage_inst_dmem_n14543), .ZN(MEM_stage_inst_dmem_n11984) );
NAND2_X1 MEM_stage_inst_dmem_U11434 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n14554), .ZN(MEM_stage_inst_dmem_n14543) );
NAND2_X1 MEM_stage_inst_dmem_U11433 ( .A1(MEM_stage_inst_dmem_ram_661), .A2(MEM_stage_inst_dmem_n14553), .ZN(MEM_stage_inst_dmem_n14544) );
NAND2_X1 MEM_stage_inst_dmem_U11432 ( .A1(MEM_stage_inst_dmem_n14542), .A2(MEM_stage_inst_dmem_n14541), .ZN(MEM_stage_inst_dmem_n11985) );
NAND2_X1 MEM_stage_inst_dmem_U11431 ( .A1(MEM_stage_inst_dmem_n14717), .A2(MEM_stage_inst_dmem_n14554), .ZN(MEM_stage_inst_dmem_n14541) );
NAND2_X1 MEM_stage_inst_dmem_U11430 ( .A1(MEM_stage_inst_dmem_ram_662), .A2(MEM_stage_inst_dmem_n14553), .ZN(MEM_stage_inst_dmem_n14542) );
NAND2_X1 MEM_stage_inst_dmem_U11429 ( .A1(MEM_stage_inst_dmem_n14540), .A2(MEM_stage_inst_dmem_n14539), .ZN(MEM_stage_inst_dmem_n11986) );
NAND2_X1 MEM_stage_inst_dmem_U11428 ( .A1(MEM_stage_inst_dmem_n16361), .A2(MEM_stage_inst_dmem_n14554), .ZN(MEM_stage_inst_dmem_n14539) );
NAND2_X1 MEM_stage_inst_dmem_U11427 ( .A1(MEM_stage_inst_dmem_ram_663), .A2(MEM_stage_inst_dmem_n14553), .ZN(MEM_stage_inst_dmem_n14540) );
NAND2_X1 MEM_stage_inst_dmem_U11426 ( .A1(MEM_stage_inst_dmem_n14538), .A2(MEM_stage_inst_dmem_n14537), .ZN(MEM_stage_inst_dmem_n11987) );
NAND2_X1 MEM_stage_inst_dmem_U11425 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n14554), .ZN(MEM_stage_inst_dmem_n14537) );
NAND2_X1 MEM_stage_inst_dmem_U11424 ( .A1(MEM_stage_inst_dmem_ram_664), .A2(MEM_stage_inst_dmem_n14553), .ZN(MEM_stage_inst_dmem_n14538) );
NAND2_X1 MEM_stage_inst_dmem_U11423 ( .A1(MEM_stage_inst_dmem_n14536), .A2(MEM_stage_inst_dmem_n14535), .ZN(MEM_stage_inst_dmem_n11988) );
NAND2_X1 MEM_stage_inst_dmem_U11422 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n14554), .ZN(MEM_stage_inst_dmem_n14535) );
NAND2_X1 MEM_stage_inst_dmem_U11421 ( .A1(MEM_stage_inst_dmem_ram_665), .A2(MEM_stage_inst_dmem_n14553), .ZN(MEM_stage_inst_dmem_n14536) );
NAND2_X1 MEM_stage_inst_dmem_U11420 ( .A1(MEM_stage_inst_dmem_n14534), .A2(MEM_stage_inst_dmem_n14533), .ZN(MEM_stage_inst_dmem_n11989) );
NAND2_X1 MEM_stage_inst_dmem_U11419 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n14554), .ZN(MEM_stage_inst_dmem_n14533) );
NAND2_X1 MEM_stage_inst_dmem_U11418 ( .A1(MEM_stage_inst_dmem_ram_666), .A2(MEM_stage_inst_dmem_n14553), .ZN(MEM_stage_inst_dmem_n14534) );
NAND2_X1 MEM_stage_inst_dmem_U11417 ( .A1(MEM_stage_inst_dmem_n14532), .A2(MEM_stage_inst_dmem_n14531), .ZN(MEM_stage_inst_dmem_n11990) );
NAND2_X1 MEM_stage_inst_dmem_U11416 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n14554), .ZN(MEM_stage_inst_dmem_n14531) );
NAND2_X1 MEM_stage_inst_dmem_U11415 ( .A1(MEM_stage_inst_dmem_ram_667), .A2(MEM_stage_inst_dmem_n14553), .ZN(MEM_stage_inst_dmem_n14532) );
NAND2_X1 MEM_stage_inst_dmem_U11414 ( .A1(MEM_stage_inst_dmem_n14530), .A2(MEM_stage_inst_dmem_n14529), .ZN(MEM_stage_inst_dmem_n11991) );
NAND2_X1 MEM_stage_inst_dmem_U11413 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n14554), .ZN(MEM_stage_inst_dmem_n14529) );
NAND2_X1 MEM_stage_inst_dmem_U11412 ( .A1(MEM_stage_inst_dmem_ram_668), .A2(MEM_stage_inst_dmem_n14553), .ZN(MEM_stage_inst_dmem_n14530) );
NAND2_X1 MEM_stage_inst_dmem_U11411 ( .A1(MEM_stage_inst_dmem_n14528), .A2(MEM_stage_inst_dmem_n14527), .ZN(MEM_stage_inst_dmem_n11992) );
NAND2_X1 MEM_stage_inst_dmem_U11410 ( .A1(MEM_stage_inst_dmem_n116), .A2(MEM_stage_inst_dmem_n14554), .ZN(MEM_stage_inst_dmem_n14527) );
NAND2_X1 MEM_stage_inst_dmem_U11409 ( .A1(MEM_stage_inst_dmem_ram_669), .A2(MEM_stage_inst_dmem_n14553), .ZN(MEM_stage_inst_dmem_n14528) );
NAND2_X1 MEM_stage_inst_dmem_U11408 ( .A1(MEM_stage_inst_dmem_n14526), .A2(MEM_stage_inst_dmem_n14525), .ZN(MEM_stage_inst_dmem_n11993) );
NAND2_X1 MEM_stage_inst_dmem_U11407 ( .A1(MEM_stage_inst_dmem_n14696), .A2(MEM_stage_inst_dmem_n14554), .ZN(MEM_stage_inst_dmem_n14525) );
NAND2_X1 MEM_stage_inst_dmem_U11406 ( .A1(MEM_stage_inst_dmem_ram_670), .A2(MEM_stage_inst_dmem_n14553), .ZN(MEM_stage_inst_dmem_n14526) );
NAND2_X1 MEM_stage_inst_dmem_U11405 ( .A1(MEM_stage_inst_dmem_n14524), .A2(MEM_stage_inst_dmem_n14523), .ZN(MEM_stage_inst_dmem_n11994) );
NAND2_X1 MEM_stage_inst_dmem_U11404 ( .A1(MEM_stage_inst_dmem_n16343), .A2(MEM_stage_inst_dmem_n14554), .ZN(MEM_stage_inst_dmem_n14523) );
INV_X1 MEM_stage_inst_dmem_U11403 ( .A(MEM_stage_inst_dmem_n14553), .ZN(MEM_stage_inst_dmem_n14554) );
NAND2_X1 MEM_stage_inst_dmem_U11402 ( .A1(MEM_stage_inst_dmem_ram_671), .A2(MEM_stage_inst_dmem_n14553), .ZN(MEM_stage_inst_dmem_n14524) );
NAND2_X1 MEM_stage_inst_dmem_U11401 ( .A1(MEM_stage_inst_dmem_n21144), .A2(MEM_stage_inst_dmem_n14837), .ZN(MEM_stage_inst_dmem_n14553) );
NAND2_X1 MEM_stage_inst_dmem_U11400 ( .A1(MEM_stage_inst_dmem_n14522), .A2(MEM_stage_inst_dmem_n14521), .ZN(MEM_stage_inst_dmem_n11995) );
NAND2_X1 MEM_stage_inst_dmem_U11399 ( .A1(MEM_stage_inst_dmem_n14732), .A2(MEM_stage_inst_dmem_n14520), .ZN(MEM_stage_inst_dmem_n14521) );
NAND2_X1 MEM_stage_inst_dmem_U11398 ( .A1(MEM_stage_inst_dmem_ram_672), .A2(MEM_stage_inst_dmem_n14519), .ZN(MEM_stage_inst_dmem_n14522) );
NAND2_X1 MEM_stage_inst_dmem_U11397 ( .A1(MEM_stage_inst_dmem_n14518), .A2(MEM_stage_inst_dmem_n14517), .ZN(MEM_stage_inst_dmem_n11996) );
NAND2_X1 MEM_stage_inst_dmem_U11396 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n14520), .ZN(MEM_stage_inst_dmem_n14517) );
NAND2_X1 MEM_stage_inst_dmem_U11395 ( .A1(MEM_stage_inst_dmem_ram_673), .A2(MEM_stage_inst_dmem_n14519), .ZN(MEM_stage_inst_dmem_n14518) );
NAND2_X1 MEM_stage_inst_dmem_U11394 ( .A1(MEM_stage_inst_dmem_n14516), .A2(MEM_stage_inst_dmem_n14515), .ZN(MEM_stage_inst_dmem_n11997) );
NAND2_X1 MEM_stage_inst_dmem_U11393 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n14520), .ZN(MEM_stage_inst_dmem_n14515) );
NAND2_X1 MEM_stage_inst_dmem_U11392 ( .A1(MEM_stage_inst_dmem_ram_674), .A2(MEM_stage_inst_dmem_n14519), .ZN(MEM_stage_inst_dmem_n14516) );
NAND2_X1 MEM_stage_inst_dmem_U11391 ( .A1(MEM_stage_inst_dmem_n14514), .A2(MEM_stage_inst_dmem_n14513), .ZN(MEM_stage_inst_dmem_n11998) );
NAND2_X1 MEM_stage_inst_dmem_U11390 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n14520), .ZN(MEM_stage_inst_dmem_n14513) );
NAND2_X1 MEM_stage_inst_dmem_U11389 ( .A1(MEM_stage_inst_dmem_ram_675), .A2(MEM_stage_inst_dmem_n14519), .ZN(MEM_stage_inst_dmem_n14514) );
NAND2_X1 MEM_stage_inst_dmem_U11388 ( .A1(MEM_stage_inst_dmem_n14512), .A2(MEM_stage_inst_dmem_n14511), .ZN(MEM_stage_inst_dmem_n11999) );
NAND2_X1 MEM_stage_inst_dmem_U11387 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n14520), .ZN(MEM_stage_inst_dmem_n14511) );
NAND2_X1 MEM_stage_inst_dmem_U11386 ( .A1(MEM_stage_inst_dmem_ram_676), .A2(MEM_stage_inst_dmem_n14519), .ZN(MEM_stage_inst_dmem_n14512) );
NAND2_X1 MEM_stage_inst_dmem_U11385 ( .A1(MEM_stage_inst_dmem_n14510), .A2(MEM_stage_inst_dmem_n14509), .ZN(MEM_stage_inst_dmem_n12000) );
NAND2_X1 MEM_stage_inst_dmem_U11384 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n14520), .ZN(MEM_stage_inst_dmem_n14509) );
NAND2_X1 MEM_stage_inst_dmem_U11383 ( .A1(MEM_stage_inst_dmem_ram_677), .A2(MEM_stage_inst_dmem_n14519), .ZN(MEM_stage_inst_dmem_n14510) );
NAND2_X1 MEM_stage_inst_dmem_U11382 ( .A1(MEM_stage_inst_dmem_n14508), .A2(MEM_stage_inst_dmem_n14507), .ZN(MEM_stage_inst_dmem_n12001) );
NAND2_X1 MEM_stage_inst_dmem_U11381 ( .A1(MEM_stage_inst_dmem_n14717), .A2(MEM_stage_inst_dmem_n14520), .ZN(MEM_stage_inst_dmem_n14507) );
NAND2_X1 MEM_stage_inst_dmem_U11380 ( .A1(MEM_stage_inst_dmem_ram_678), .A2(MEM_stage_inst_dmem_n14519), .ZN(MEM_stage_inst_dmem_n14508) );
NAND2_X1 MEM_stage_inst_dmem_U11379 ( .A1(MEM_stage_inst_dmem_n14506), .A2(MEM_stage_inst_dmem_n14505), .ZN(MEM_stage_inst_dmem_n12002) );
NAND2_X1 MEM_stage_inst_dmem_U11378 ( .A1(MEM_stage_inst_dmem_n112), .A2(MEM_stage_inst_dmem_n14520), .ZN(MEM_stage_inst_dmem_n14505) );
NAND2_X1 MEM_stage_inst_dmem_U11377 ( .A1(MEM_stage_inst_dmem_ram_679), .A2(MEM_stage_inst_dmem_n14519), .ZN(MEM_stage_inst_dmem_n14506) );
NAND2_X1 MEM_stage_inst_dmem_U11376 ( .A1(MEM_stage_inst_dmem_n14504), .A2(MEM_stage_inst_dmem_n14503), .ZN(MEM_stage_inst_dmem_n12003) );
NAND2_X1 MEM_stage_inst_dmem_U11375 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n14520), .ZN(MEM_stage_inst_dmem_n14503) );
NAND2_X1 MEM_stage_inst_dmem_U11374 ( .A1(MEM_stage_inst_dmem_ram_680), .A2(MEM_stage_inst_dmem_n14519), .ZN(MEM_stage_inst_dmem_n14504) );
NAND2_X1 MEM_stage_inst_dmem_U11373 ( .A1(MEM_stage_inst_dmem_n14502), .A2(MEM_stage_inst_dmem_n14501), .ZN(MEM_stage_inst_dmem_n12004) );
NAND2_X1 MEM_stage_inst_dmem_U11372 ( .A1(MEM_stage_inst_dmem_n16772), .A2(MEM_stage_inst_dmem_n14520), .ZN(MEM_stage_inst_dmem_n14501) );
NAND2_X1 MEM_stage_inst_dmem_U11371 ( .A1(MEM_stage_inst_dmem_ram_681), .A2(MEM_stage_inst_dmem_n14519), .ZN(MEM_stage_inst_dmem_n14502) );
NAND2_X1 MEM_stage_inst_dmem_U11370 ( .A1(MEM_stage_inst_dmem_n14500), .A2(MEM_stage_inst_dmem_n14499), .ZN(MEM_stage_inst_dmem_n12005) );
NAND2_X1 MEM_stage_inst_dmem_U11369 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n14520), .ZN(MEM_stage_inst_dmem_n14499) );
NAND2_X1 MEM_stage_inst_dmem_U11368 ( .A1(MEM_stage_inst_dmem_ram_682), .A2(MEM_stage_inst_dmem_n14519), .ZN(MEM_stage_inst_dmem_n14500) );
NAND2_X1 MEM_stage_inst_dmem_U11367 ( .A1(MEM_stage_inst_dmem_n14498), .A2(MEM_stage_inst_dmem_n14497), .ZN(MEM_stage_inst_dmem_n12006) );
NAND2_X1 MEM_stage_inst_dmem_U11366 ( .A1(MEM_stage_inst_dmem_n20904), .A2(MEM_stage_inst_dmem_n14520), .ZN(MEM_stage_inst_dmem_n14497) );
NAND2_X1 MEM_stage_inst_dmem_U11365 ( .A1(MEM_stage_inst_dmem_ram_683), .A2(MEM_stage_inst_dmem_n14519), .ZN(MEM_stage_inst_dmem_n14498) );
NAND2_X1 MEM_stage_inst_dmem_U11364 ( .A1(MEM_stage_inst_dmem_n14496), .A2(MEM_stage_inst_dmem_n14495), .ZN(MEM_stage_inst_dmem_n12007) );
NAND2_X1 MEM_stage_inst_dmem_U11363 ( .A1(MEM_stage_inst_dmem_n21474), .A2(MEM_stage_inst_dmem_n14520), .ZN(MEM_stage_inst_dmem_n14495) );
NAND2_X1 MEM_stage_inst_dmem_U11362 ( .A1(MEM_stage_inst_dmem_ram_684), .A2(MEM_stage_inst_dmem_n14519), .ZN(MEM_stage_inst_dmem_n14496) );
NAND2_X1 MEM_stage_inst_dmem_U11361 ( .A1(MEM_stage_inst_dmem_n14494), .A2(MEM_stage_inst_dmem_n14493), .ZN(MEM_stage_inst_dmem_n12008) );
NAND2_X1 MEM_stage_inst_dmem_U11360 ( .A1(MEM_stage_inst_dmem_n116), .A2(MEM_stage_inst_dmem_n14520), .ZN(MEM_stage_inst_dmem_n14493) );
NAND2_X1 MEM_stage_inst_dmem_U11359 ( .A1(MEM_stage_inst_dmem_ram_685), .A2(MEM_stage_inst_dmem_n14519), .ZN(MEM_stage_inst_dmem_n14494) );
NAND2_X1 MEM_stage_inst_dmem_U11358 ( .A1(MEM_stage_inst_dmem_n14492), .A2(MEM_stage_inst_dmem_n14491), .ZN(MEM_stage_inst_dmem_n12009) );
NAND2_X1 MEM_stage_inst_dmem_U11357 ( .A1(MEM_stage_inst_dmem_n14696), .A2(MEM_stage_inst_dmem_n14520), .ZN(MEM_stage_inst_dmem_n14491) );
NAND2_X1 MEM_stage_inst_dmem_U11356 ( .A1(MEM_stage_inst_dmem_ram_686), .A2(MEM_stage_inst_dmem_n14519), .ZN(MEM_stage_inst_dmem_n14492) );
NAND2_X1 MEM_stage_inst_dmem_U11355 ( .A1(MEM_stage_inst_dmem_n14490), .A2(MEM_stage_inst_dmem_n14489), .ZN(MEM_stage_inst_dmem_n12010) );
NAND2_X1 MEM_stage_inst_dmem_U11354 ( .A1(MEM_stage_inst_dmem_n14693), .A2(MEM_stage_inst_dmem_n14520), .ZN(MEM_stage_inst_dmem_n14489) );
INV_X1 MEM_stage_inst_dmem_U11353 ( .A(MEM_stage_inst_dmem_n14519), .ZN(MEM_stage_inst_dmem_n14520) );
NAND2_X1 MEM_stage_inst_dmem_U11352 ( .A1(MEM_stage_inst_dmem_ram_687), .A2(MEM_stage_inst_dmem_n14519), .ZN(MEM_stage_inst_dmem_n14490) );
NAND2_X1 MEM_stage_inst_dmem_U11351 ( .A1(MEM_stage_inst_dmem_n21109), .A2(MEM_stage_inst_dmem_n14837), .ZN(MEM_stage_inst_dmem_n14519) );
NAND2_X1 MEM_stage_inst_dmem_U11350 ( .A1(MEM_stage_inst_dmem_n14488), .A2(MEM_stage_inst_dmem_n14487), .ZN(MEM_stage_inst_dmem_n12011) );
NAND2_X1 MEM_stage_inst_dmem_U11349 ( .A1(MEM_stage_inst_dmem_n14732), .A2(MEM_stage_inst_dmem_n14486), .ZN(MEM_stage_inst_dmem_n14487) );
NAND2_X1 MEM_stage_inst_dmem_U11348 ( .A1(MEM_stage_inst_dmem_ram_688), .A2(MEM_stage_inst_dmem_n14485), .ZN(MEM_stage_inst_dmem_n14488) );
NAND2_X1 MEM_stage_inst_dmem_U11347 ( .A1(MEM_stage_inst_dmem_n14484), .A2(MEM_stage_inst_dmem_n14483), .ZN(MEM_stage_inst_dmem_n12012) );
NAND2_X1 MEM_stage_inst_dmem_U11346 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n14486), .ZN(MEM_stage_inst_dmem_n14483) );
NAND2_X1 MEM_stage_inst_dmem_U11345 ( .A1(MEM_stage_inst_dmem_ram_689), .A2(MEM_stage_inst_dmem_n14485), .ZN(MEM_stage_inst_dmem_n14484) );
NAND2_X1 MEM_stage_inst_dmem_U11344 ( .A1(MEM_stage_inst_dmem_n14482), .A2(MEM_stage_inst_dmem_n14481), .ZN(MEM_stage_inst_dmem_n12013) );
NAND2_X1 MEM_stage_inst_dmem_U11343 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n14486), .ZN(MEM_stage_inst_dmem_n14481) );
NAND2_X1 MEM_stage_inst_dmem_U11342 ( .A1(MEM_stage_inst_dmem_ram_690), .A2(MEM_stage_inst_dmem_n14485), .ZN(MEM_stage_inst_dmem_n14482) );
NAND2_X1 MEM_stage_inst_dmem_U11341 ( .A1(MEM_stage_inst_dmem_n14480), .A2(MEM_stage_inst_dmem_n14479), .ZN(MEM_stage_inst_dmem_n12014) );
NAND2_X1 MEM_stage_inst_dmem_U11340 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n14486), .ZN(MEM_stage_inst_dmem_n14479) );
NAND2_X1 MEM_stage_inst_dmem_U11339 ( .A1(MEM_stage_inst_dmem_ram_691), .A2(MEM_stage_inst_dmem_n14485), .ZN(MEM_stage_inst_dmem_n14480) );
NAND2_X1 MEM_stage_inst_dmem_U11338 ( .A1(MEM_stage_inst_dmem_n14478), .A2(MEM_stage_inst_dmem_n14477), .ZN(MEM_stage_inst_dmem_n12015) );
NAND2_X1 MEM_stage_inst_dmem_U11337 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n14486), .ZN(MEM_stage_inst_dmem_n14477) );
NAND2_X1 MEM_stage_inst_dmem_U11336 ( .A1(MEM_stage_inst_dmem_ram_692), .A2(MEM_stage_inst_dmem_n14485), .ZN(MEM_stage_inst_dmem_n14478) );
NAND2_X1 MEM_stage_inst_dmem_U11335 ( .A1(MEM_stage_inst_dmem_n14476), .A2(MEM_stage_inst_dmem_n14475), .ZN(MEM_stage_inst_dmem_n12016) );
NAND2_X1 MEM_stage_inst_dmem_U11334 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n14486), .ZN(MEM_stage_inst_dmem_n14475) );
NAND2_X1 MEM_stage_inst_dmem_U11333 ( .A1(MEM_stage_inst_dmem_ram_693), .A2(MEM_stage_inst_dmem_n14485), .ZN(MEM_stage_inst_dmem_n14476) );
NAND2_X1 MEM_stage_inst_dmem_U11332 ( .A1(MEM_stage_inst_dmem_n14474), .A2(MEM_stage_inst_dmem_n14473), .ZN(MEM_stage_inst_dmem_n12017) );
NAND2_X1 MEM_stage_inst_dmem_U11331 ( .A1(MEM_stage_inst_dmem_n14717), .A2(MEM_stage_inst_dmem_n14486), .ZN(MEM_stage_inst_dmem_n14473) );
NAND2_X1 MEM_stage_inst_dmem_U11330 ( .A1(MEM_stage_inst_dmem_ram_694), .A2(MEM_stage_inst_dmem_n14485), .ZN(MEM_stage_inst_dmem_n14474) );
NAND2_X1 MEM_stage_inst_dmem_U11329 ( .A1(MEM_stage_inst_dmem_n14472), .A2(MEM_stage_inst_dmem_n14471), .ZN(MEM_stage_inst_dmem_n12018) );
NAND2_X1 MEM_stage_inst_dmem_U11328 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n14486), .ZN(MEM_stage_inst_dmem_n14471) );
NAND2_X1 MEM_stage_inst_dmem_U11327 ( .A1(MEM_stage_inst_dmem_ram_695), .A2(MEM_stage_inst_dmem_n14485), .ZN(MEM_stage_inst_dmem_n14472) );
NAND2_X1 MEM_stage_inst_dmem_U11326 ( .A1(MEM_stage_inst_dmem_n14470), .A2(MEM_stage_inst_dmem_n14469), .ZN(MEM_stage_inst_dmem_n12019) );
NAND2_X1 MEM_stage_inst_dmem_U11325 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n14486), .ZN(MEM_stage_inst_dmem_n14469) );
NAND2_X1 MEM_stage_inst_dmem_U11324 ( .A1(MEM_stage_inst_dmem_ram_696), .A2(MEM_stage_inst_dmem_n14485), .ZN(MEM_stage_inst_dmem_n14470) );
NAND2_X1 MEM_stage_inst_dmem_U11323 ( .A1(MEM_stage_inst_dmem_n14468), .A2(MEM_stage_inst_dmem_n14467), .ZN(MEM_stage_inst_dmem_n12020) );
NAND2_X1 MEM_stage_inst_dmem_U11322 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n14486), .ZN(MEM_stage_inst_dmem_n14467) );
NAND2_X1 MEM_stage_inst_dmem_U11321 ( .A1(MEM_stage_inst_dmem_ram_697), .A2(MEM_stage_inst_dmem_n14485), .ZN(MEM_stage_inst_dmem_n14468) );
NAND2_X1 MEM_stage_inst_dmem_U11320 ( .A1(MEM_stage_inst_dmem_n14466), .A2(MEM_stage_inst_dmem_n14465), .ZN(MEM_stage_inst_dmem_n12021) );
NAND2_X1 MEM_stage_inst_dmem_U11319 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n14486), .ZN(MEM_stage_inst_dmem_n14465) );
NAND2_X1 MEM_stage_inst_dmem_U11318 ( .A1(MEM_stage_inst_dmem_ram_698), .A2(MEM_stage_inst_dmem_n14485), .ZN(MEM_stage_inst_dmem_n14466) );
NAND2_X1 MEM_stage_inst_dmem_U11317 ( .A1(MEM_stage_inst_dmem_n14464), .A2(MEM_stage_inst_dmem_n14463), .ZN(MEM_stage_inst_dmem_n12022) );
NAND2_X1 MEM_stage_inst_dmem_U11316 ( .A1(MEM_stage_inst_dmem_n14705), .A2(MEM_stage_inst_dmem_n14486), .ZN(MEM_stage_inst_dmem_n14463) );
NAND2_X1 MEM_stage_inst_dmem_U11315 ( .A1(MEM_stage_inst_dmem_ram_699), .A2(MEM_stage_inst_dmem_n14485), .ZN(MEM_stage_inst_dmem_n14464) );
NAND2_X1 MEM_stage_inst_dmem_U11314 ( .A1(MEM_stage_inst_dmem_n14462), .A2(MEM_stage_inst_dmem_n14461), .ZN(MEM_stage_inst_dmem_n12023) );
NAND2_X1 MEM_stage_inst_dmem_U11313 ( .A1(MEM_stage_inst_dmem_n14702), .A2(MEM_stage_inst_dmem_n14486), .ZN(MEM_stage_inst_dmem_n14461) );
NAND2_X1 MEM_stage_inst_dmem_U11312 ( .A1(MEM_stage_inst_dmem_ram_700), .A2(MEM_stage_inst_dmem_n14485), .ZN(MEM_stage_inst_dmem_n14462) );
NAND2_X1 MEM_stage_inst_dmem_U11311 ( .A1(MEM_stage_inst_dmem_n14460), .A2(MEM_stage_inst_dmem_n14459), .ZN(MEM_stage_inst_dmem_n12024) );
NAND2_X1 MEM_stage_inst_dmem_U11310 ( .A1(MEM_stage_inst_dmem_n116), .A2(MEM_stage_inst_dmem_n14486), .ZN(MEM_stage_inst_dmem_n14459) );
NAND2_X1 MEM_stage_inst_dmem_U11309 ( .A1(MEM_stage_inst_dmem_ram_701), .A2(MEM_stage_inst_dmem_n14485), .ZN(MEM_stage_inst_dmem_n14460) );
NAND2_X1 MEM_stage_inst_dmem_U11308 ( .A1(MEM_stage_inst_dmem_n14458), .A2(MEM_stage_inst_dmem_n14457), .ZN(MEM_stage_inst_dmem_n12025) );
NAND2_X1 MEM_stage_inst_dmem_U11307 ( .A1(MEM_stage_inst_dmem_n14696), .A2(MEM_stage_inst_dmem_n14486), .ZN(MEM_stage_inst_dmem_n14457) );
NAND2_X1 MEM_stage_inst_dmem_U11306 ( .A1(MEM_stage_inst_dmem_ram_702), .A2(MEM_stage_inst_dmem_n14485), .ZN(MEM_stage_inst_dmem_n14458) );
NAND2_X1 MEM_stage_inst_dmem_U11305 ( .A1(MEM_stage_inst_dmem_n14456), .A2(MEM_stage_inst_dmem_n14455), .ZN(MEM_stage_inst_dmem_n12026) );
NAND2_X1 MEM_stage_inst_dmem_U11304 ( .A1(MEM_stage_inst_dmem_n15110), .A2(MEM_stage_inst_dmem_n14486), .ZN(MEM_stage_inst_dmem_n14455) );
INV_X1 MEM_stage_inst_dmem_U11303 ( .A(MEM_stage_inst_dmem_n14485), .ZN(MEM_stage_inst_dmem_n14486) );
NAND2_X1 MEM_stage_inst_dmem_U11302 ( .A1(MEM_stage_inst_dmem_ram_703), .A2(MEM_stage_inst_dmem_n14485), .ZN(MEM_stage_inst_dmem_n14456) );
NAND2_X1 MEM_stage_inst_dmem_U11301 ( .A1(MEM_stage_inst_dmem_n21074), .A2(MEM_stage_inst_dmem_n14837), .ZN(MEM_stage_inst_dmem_n14485) );
NAND2_X1 MEM_stage_inst_dmem_U11300 ( .A1(MEM_stage_inst_dmem_n14454), .A2(MEM_stage_inst_dmem_n14453), .ZN(MEM_stage_inst_dmem_n12027) );
NAND2_X1 MEM_stage_inst_dmem_U11299 ( .A1(MEM_stage_inst_dmem_n14732), .A2(MEM_stage_inst_dmem_n14452), .ZN(MEM_stage_inst_dmem_n14453) );
NAND2_X1 MEM_stage_inst_dmem_U11298 ( .A1(MEM_stage_inst_dmem_ram_704), .A2(MEM_stage_inst_dmem_n14451), .ZN(MEM_stage_inst_dmem_n14454) );
NAND2_X1 MEM_stage_inst_dmem_U11297 ( .A1(MEM_stage_inst_dmem_n14450), .A2(MEM_stage_inst_dmem_n14449), .ZN(MEM_stage_inst_dmem_n12028) );
NAND2_X1 MEM_stage_inst_dmem_U11296 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n14452), .ZN(MEM_stage_inst_dmem_n14449) );
NAND2_X1 MEM_stage_inst_dmem_U11295 ( .A1(MEM_stage_inst_dmem_ram_705), .A2(MEM_stage_inst_dmem_n14451), .ZN(MEM_stage_inst_dmem_n14450) );
NAND2_X1 MEM_stage_inst_dmem_U11294 ( .A1(MEM_stage_inst_dmem_n14448), .A2(MEM_stage_inst_dmem_n14447), .ZN(MEM_stage_inst_dmem_n12029) );
NAND2_X1 MEM_stage_inst_dmem_U11293 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n14452), .ZN(MEM_stage_inst_dmem_n14447) );
NAND2_X1 MEM_stage_inst_dmem_U11292 ( .A1(MEM_stage_inst_dmem_ram_706), .A2(MEM_stage_inst_dmem_n14451), .ZN(MEM_stage_inst_dmem_n14448) );
NAND2_X1 MEM_stage_inst_dmem_U11291 ( .A1(MEM_stage_inst_dmem_n14446), .A2(MEM_stage_inst_dmem_n14445), .ZN(MEM_stage_inst_dmem_n12030) );
NAND2_X1 MEM_stage_inst_dmem_U11290 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n14452), .ZN(MEM_stage_inst_dmem_n14445) );
NAND2_X1 MEM_stage_inst_dmem_U11289 ( .A1(MEM_stage_inst_dmem_ram_707), .A2(MEM_stage_inst_dmem_n14451), .ZN(MEM_stage_inst_dmem_n14446) );
NAND2_X1 MEM_stage_inst_dmem_U11288 ( .A1(MEM_stage_inst_dmem_n14444), .A2(MEM_stage_inst_dmem_n14443), .ZN(MEM_stage_inst_dmem_n12031) );
NAND2_X1 MEM_stage_inst_dmem_U11287 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n14452), .ZN(MEM_stage_inst_dmem_n14443) );
NAND2_X1 MEM_stage_inst_dmem_U11286 ( .A1(MEM_stage_inst_dmem_ram_708), .A2(MEM_stage_inst_dmem_n14451), .ZN(MEM_stage_inst_dmem_n14444) );
NAND2_X1 MEM_stage_inst_dmem_U11285 ( .A1(MEM_stage_inst_dmem_n14442), .A2(MEM_stage_inst_dmem_n14441), .ZN(MEM_stage_inst_dmem_n12032) );
NAND2_X1 MEM_stage_inst_dmem_U11284 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n14452), .ZN(MEM_stage_inst_dmem_n14441) );
NAND2_X1 MEM_stage_inst_dmem_U11283 ( .A1(MEM_stage_inst_dmem_ram_709), .A2(MEM_stage_inst_dmem_n14451), .ZN(MEM_stage_inst_dmem_n14442) );
NAND2_X1 MEM_stage_inst_dmem_U11282 ( .A1(MEM_stage_inst_dmem_n14440), .A2(MEM_stage_inst_dmem_n14439), .ZN(MEM_stage_inst_dmem_n12033) );
NAND2_X1 MEM_stage_inst_dmem_U11281 ( .A1(MEM_stage_inst_dmem_n14717), .A2(MEM_stage_inst_dmem_n14452), .ZN(MEM_stage_inst_dmem_n14439) );
NAND2_X1 MEM_stage_inst_dmem_U11280 ( .A1(MEM_stage_inst_dmem_ram_710), .A2(MEM_stage_inst_dmem_n14451), .ZN(MEM_stage_inst_dmem_n14440) );
NAND2_X1 MEM_stage_inst_dmem_U11279 ( .A1(MEM_stage_inst_dmem_n14438), .A2(MEM_stage_inst_dmem_n14437), .ZN(MEM_stage_inst_dmem_n12034) );
NAND2_X1 MEM_stage_inst_dmem_U11278 ( .A1(MEM_stage_inst_dmem_n16361), .A2(MEM_stage_inst_dmem_n14452), .ZN(MEM_stage_inst_dmem_n14437) );
NAND2_X1 MEM_stage_inst_dmem_U11277 ( .A1(MEM_stage_inst_dmem_ram_711), .A2(MEM_stage_inst_dmem_n14451), .ZN(MEM_stage_inst_dmem_n14438) );
NAND2_X1 MEM_stage_inst_dmem_U11276 ( .A1(MEM_stage_inst_dmem_n14436), .A2(MEM_stage_inst_dmem_n14435), .ZN(MEM_stage_inst_dmem_n12035) );
NAND2_X1 MEM_stage_inst_dmem_U11275 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n14452), .ZN(MEM_stage_inst_dmem_n14435) );
NAND2_X1 MEM_stage_inst_dmem_U11274 ( .A1(MEM_stage_inst_dmem_ram_712), .A2(MEM_stage_inst_dmem_n14451), .ZN(MEM_stage_inst_dmem_n14436) );
NAND2_X1 MEM_stage_inst_dmem_U11273 ( .A1(MEM_stage_inst_dmem_n14434), .A2(MEM_stage_inst_dmem_n14433), .ZN(MEM_stage_inst_dmem_n12036) );
NAND2_X1 MEM_stage_inst_dmem_U11272 ( .A1(MEM_stage_inst_dmem_n19251), .A2(MEM_stage_inst_dmem_n14452), .ZN(MEM_stage_inst_dmem_n14433) );
NAND2_X1 MEM_stage_inst_dmem_U11271 ( .A1(MEM_stage_inst_dmem_ram_713), .A2(MEM_stage_inst_dmem_n14451), .ZN(MEM_stage_inst_dmem_n14434) );
NAND2_X1 MEM_stage_inst_dmem_U11270 ( .A1(MEM_stage_inst_dmem_n14432), .A2(MEM_stage_inst_dmem_n14431), .ZN(MEM_stage_inst_dmem_n12037) );
NAND2_X1 MEM_stage_inst_dmem_U11269 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n14452), .ZN(MEM_stage_inst_dmem_n14431) );
NAND2_X1 MEM_stage_inst_dmem_U11268 ( .A1(MEM_stage_inst_dmem_ram_714), .A2(MEM_stage_inst_dmem_n14451), .ZN(MEM_stage_inst_dmem_n14432) );
NAND2_X1 MEM_stage_inst_dmem_U11267 ( .A1(MEM_stage_inst_dmem_n14430), .A2(MEM_stage_inst_dmem_n14429), .ZN(MEM_stage_inst_dmem_n12038) );
NAND2_X1 MEM_stage_inst_dmem_U11266 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n14452), .ZN(MEM_stage_inst_dmem_n14429) );
NAND2_X1 MEM_stage_inst_dmem_U11265 ( .A1(MEM_stage_inst_dmem_ram_715), .A2(MEM_stage_inst_dmem_n14451), .ZN(MEM_stage_inst_dmem_n14430) );
NAND2_X1 MEM_stage_inst_dmem_U11264 ( .A1(MEM_stage_inst_dmem_n14428), .A2(MEM_stage_inst_dmem_n14427), .ZN(MEM_stage_inst_dmem_n12039) );
NAND2_X1 MEM_stage_inst_dmem_U11263 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n14452), .ZN(MEM_stage_inst_dmem_n14427) );
NAND2_X1 MEM_stage_inst_dmem_U11262 ( .A1(MEM_stage_inst_dmem_ram_716), .A2(MEM_stage_inst_dmem_n14451), .ZN(MEM_stage_inst_dmem_n14428) );
NAND2_X1 MEM_stage_inst_dmem_U11261 ( .A1(MEM_stage_inst_dmem_n14426), .A2(MEM_stage_inst_dmem_n14425), .ZN(MEM_stage_inst_dmem_n12040) );
NAND2_X1 MEM_stage_inst_dmem_U11260 ( .A1(MEM_stage_inst_dmem_n116), .A2(MEM_stage_inst_dmem_n14452), .ZN(MEM_stage_inst_dmem_n14425) );
NAND2_X1 MEM_stage_inst_dmem_U11259 ( .A1(MEM_stage_inst_dmem_ram_717), .A2(MEM_stage_inst_dmem_n14451), .ZN(MEM_stage_inst_dmem_n14426) );
NAND2_X1 MEM_stage_inst_dmem_U11258 ( .A1(MEM_stage_inst_dmem_n14424), .A2(MEM_stage_inst_dmem_n14423), .ZN(MEM_stage_inst_dmem_n12041) );
NAND2_X1 MEM_stage_inst_dmem_U11257 ( .A1(MEM_stage_inst_dmem_n14696), .A2(MEM_stage_inst_dmem_n14452), .ZN(MEM_stage_inst_dmem_n14423) );
NAND2_X1 MEM_stage_inst_dmem_U11256 ( .A1(MEM_stage_inst_dmem_ram_718), .A2(MEM_stage_inst_dmem_n14451), .ZN(MEM_stage_inst_dmem_n14424) );
NAND2_X1 MEM_stage_inst_dmem_U11255 ( .A1(MEM_stage_inst_dmem_n14422), .A2(MEM_stage_inst_dmem_n14421), .ZN(MEM_stage_inst_dmem_n12042) );
NAND2_X1 MEM_stage_inst_dmem_U11254 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n14452), .ZN(MEM_stage_inst_dmem_n14421) );
NAND2_X1 MEM_stage_inst_dmem_U11253 ( .A1(MEM_stage_inst_dmem_ram_719), .A2(MEM_stage_inst_dmem_n14451), .ZN(MEM_stage_inst_dmem_n14422) );
NAND2_X1 MEM_stage_inst_dmem_U11252 ( .A1(MEM_stage_inst_dmem_n21039), .A2(MEM_stage_inst_dmem_n14837), .ZN(MEM_stage_inst_dmem_n14451) );
NAND2_X1 MEM_stage_inst_dmem_U11251 ( .A1(MEM_stage_inst_dmem_n14420), .A2(MEM_stage_inst_dmem_n14419), .ZN(MEM_stage_inst_dmem_n12043) );
NAND2_X1 MEM_stage_inst_dmem_U11250 ( .A1(MEM_stage_inst_dmem_n14732), .A2(MEM_stage_inst_dmem_n14418), .ZN(MEM_stage_inst_dmem_n14419) );
NAND2_X1 MEM_stage_inst_dmem_U11249 ( .A1(MEM_stage_inst_dmem_ram_720), .A2(MEM_stage_inst_dmem_n14417), .ZN(MEM_stage_inst_dmem_n14420) );
NAND2_X1 MEM_stage_inst_dmem_U11248 ( .A1(MEM_stage_inst_dmem_n14416), .A2(MEM_stage_inst_dmem_n14415), .ZN(MEM_stage_inst_dmem_n12044) );
NAND2_X1 MEM_stage_inst_dmem_U11247 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n14418), .ZN(MEM_stage_inst_dmem_n14415) );
NAND2_X1 MEM_stage_inst_dmem_U11246 ( .A1(MEM_stage_inst_dmem_ram_721), .A2(MEM_stage_inst_dmem_n14417), .ZN(MEM_stage_inst_dmem_n14416) );
NAND2_X1 MEM_stage_inst_dmem_U11245 ( .A1(MEM_stage_inst_dmem_n14414), .A2(MEM_stage_inst_dmem_n14413), .ZN(MEM_stage_inst_dmem_n12045) );
NAND2_X1 MEM_stage_inst_dmem_U11244 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n14418), .ZN(MEM_stage_inst_dmem_n14413) );
NAND2_X1 MEM_stage_inst_dmem_U11243 ( .A1(MEM_stage_inst_dmem_ram_722), .A2(MEM_stage_inst_dmem_n14417), .ZN(MEM_stage_inst_dmem_n14414) );
NAND2_X1 MEM_stage_inst_dmem_U11242 ( .A1(MEM_stage_inst_dmem_n14412), .A2(MEM_stage_inst_dmem_n14411), .ZN(MEM_stage_inst_dmem_n12046) );
NAND2_X1 MEM_stage_inst_dmem_U11241 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n14418), .ZN(MEM_stage_inst_dmem_n14411) );
NAND2_X1 MEM_stage_inst_dmem_U11240 ( .A1(MEM_stage_inst_dmem_ram_723), .A2(MEM_stage_inst_dmem_n14417), .ZN(MEM_stage_inst_dmem_n14412) );
NAND2_X1 MEM_stage_inst_dmem_U11239 ( .A1(MEM_stage_inst_dmem_n14410), .A2(MEM_stage_inst_dmem_n14409), .ZN(MEM_stage_inst_dmem_n12047) );
NAND2_X1 MEM_stage_inst_dmem_U11238 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n14418), .ZN(MEM_stage_inst_dmem_n14409) );
NAND2_X1 MEM_stage_inst_dmem_U11237 ( .A1(MEM_stage_inst_dmem_ram_724), .A2(MEM_stage_inst_dmem_n14417), .ZN(MEM_stage_inst_dmem_n14410) );
NAND2_X1 MEM_stage_inst_dmem_U11236 ( .A1(MEM_stage_inst_dmem_n14408), .A2(MEM_stage_inst_dmem_n14407), .ZN(MEM_stage_inst_dmem_n12048) );
NAND2_X1 MEM_stage_inst_dmem_U11235 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n14418), .ZN(MEM_stage_inst_dmem_n14407) );
NAND2_X1 MEM_stage_inst_dmem_U11234 ( .A1(MEM_stage_inst_dmem_ram_725), .A2(MEM_stage_inst_dmem_n14417), .ZN(MEM_stage_inst_dmem_n14408) );
NAND2_X1 MEM_stage_inst_dmem_U11233 ( .A1(MEM_stage_inst_dmem_n14406), .A2(MEM_stage_inst_dmem_n14405), .ZN(MEM_stage_inst_dmem_n12049) );
NAND2_X1 MEM_stage_inst_dmem_U11232 ( .A1(MEM_stage_inst_dmem_n14717), .A2(MEM_stage_inst_dmem_n14418), .ZN(MEM_stage_inst_dmem_n14405) );
NAND2_X1 MEM_stage_inst_dmem_U11231 ( .A1(MEM_stage_inst_dmem_ram_726), .A2(MEM_stage_inst_dmem_n14417), .ZN(MEM_stage_inst_dmem_n14406) );
NAND2_X1 MEM_stage_inst_dmem_U11230 ( .A1(MEM_stage_inst_dmem_n14404), .A2(MEM_stage_inst_dmem_n14403), .ZN(MEM_stage_inst_dmem_n12050) );
NAND2_X1 MEM_stage_inst_dmem_U11229 ( .A1(MEM_stage_inst_dmem_n16777), .A2(MEM_stage_inst_dmem_n14418), .ZN(MEM_stage_inst_dmem_n14403) );
NAND2_X1 MEM_stage_inst_dmem_U11228 ( .A1(MEM_stage_inst_dmem_ram_727), .A2(MEM_stage_inst_dmem_n14417), .ZN(MEM_stage_inst_dmem_n14404) );
NAND2_X1 MEM_stage_inst_dmem_U11227 ( .A1(MEM_stage_inst_dmem_n14402), .A2(MEM_stage_inst_dmem_n14401), .ZN(MEM_stage_inst_dmem_n12051) );
NAND2_X1 MEM_stage_inst_dmem_U11226 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n14418), .ZN(MEM_stage_inst_dmem_n14401) );
NAND2_X1 MEM_stage_inst_dmem_U11225 ( .A1(MEM_stage_inst_dmem_ram_728), .A2(MEM_stage_inst_dmem_n14417), .ZN(MEM_stage_inst_dmem_n14402) );
NAND2_X1 MEM_stage_inst_dmem_U11224 ( .A1(MEM_stage_inst_dmem_n14400), .A2(MEM_stage_inst_dmem_n14399), .ZN(MEM_stage_inst_dmem_n12052) );
NAND2_X1 MEM_stage_inst_dmem_U11223 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n14418), .ZN(MEM_stage_inst_dmem_n14399) );
NAND2_X1 MEM_stage_inst_dmem_U11222 ( .A1(MEM_stage_inst_dmem_ram_729), .A2(MEM_stage_inst_dmem_n14417), .ZN(MEM_stage_inst_dmem_n14400) );
NAND2_X1 MEM_stage_inst_dmem_U11221 ( .A1(MEM_stage_inst_dmem_n14398), .A2(MEM_stage_inst_dmem_n14397), .ZN(MEM_stage_inst_dmem_n12053) );
NAND2_X1 MEM_stage_inst_dmem_U11220 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n14418), .ZN(MEM_stage_inst_dmem_n14397) );
NAND2_X1 MEM_stage_inst_dmem_U11219 ( .A1(MEM_stage_inst_dmem_ram_730), .A2(MEM_stage_inst_dmem_n14417), .ZN(MEM_stage_inst_dmem_n14398) );
NAND2_X1 MEM_stage_inst_dmem_U11218 ( .A1(MEM_stage_inst_dmem_n14396), .A2(MEM_stage_inst_dmem_n14395), .ZN(MEM_stage_inst_dmem_n12054) );
NAND2_X1 MEM_stage_inst_dmem_U11217 ( .A1(MEM_stage_inst_dmem_n20904), .A2(MEM_stage_inst_dmem_n14418), .ZN(MEM_stage_inst_dmem_n14395) );
NAND2_X1 MEM_stage_inst_dmem_U11216 ( .A1(MEM_stage_inst_dmem_ram_731), .A2(MEM_stage_inst_dmem_n14417), .ZN(MEM_stage_inst_dmem_n14396) );
NAND2_X1 MEM_stage_inst_dmem_U11215 ( .A1(MEM_stage_inst_dmem_n14394), .A2(MEM_stage_inst_dmem_n14393), .ZN(MEM_stage_inst_dmem_n12055) );
NAND2_X1 MEM_stage_inst_dmem_U11214 ( .A1(MEM_stage_inst_dmem_n21474), .A2(MEM_stage_inst_dmem_n14418), .ZN(MEM_stage_inst_dmem_n14393) );
NAND2_X1 MEM_stage_inst_dmem_U11213 ( .A1(MEM_stage_inst_dmem_ram_732), .A2(MEM_stage_inst_dmem_n14417), .ZN(MEM_stage_inst_dmem_n14394) );
NAND2_X1 MEM_stage_inst_dmem_U11212 ( .A1(MEM_stage_inst_dmem_n14392), .A2(MEM_stage_inst_dmem_n14391), .ZN(MEM_stage_inst_dmem_n12056) );
NAND2_X1 MEM_stage_inst_dmem_U11211 ( .A1(MEM_stage_inst_dmem_n116), .A2(MEM_stage_inst_dmem_n14418), .ZN(MEM_stage_inst_dmem_n14391) );
NAND2_X1 MEM_stage_inst_dmem_U11210 ( .A1(MEM_stage_inst_dmem_ram_733), .A2(MEM_stage_inst_dmem_n14417), .ZN(MEM_stage_inst_dmem_n14392) );
NAND2_X1 MEM_stage_inst_dmem_U11209 ( .A1(MEM_stage_inst_dmem_n14390), .A2(MEM_stage_inst_dmem_n14389), .ZN(MEM_stage_inst_dmem_n12057) );
NAND2_X1 MEM_stage_inst_dmem_U11208 ( .A1(MEM_stage_inst_dmem_n14696), .A2(MEM_stage_inst_dmem_n14418), .ZN(MEM_stage_inst_dmem_n14389) );
NAND2_X1 MEM_stage_inst_dmem_U11207 ( .A1(MEM_stage_inst_dmem_ram_734), .A2(MEM_stage_inst_dmem_n14417), .ZN(MEM_stage_inst_dmem_n14390) );
NAND2_X1 MEM_stage_inst_dmem_U11206 ( .A1(MEM_stage_inst_dmem_n14388), .A2(MEM_stage_inst_dmem_n14387), .ZN(MEM_stage_inst_dmem_n12058) );
NAND2_X1 MEM_stage_inst_dmem_U11205 ( .A1(MEM_stage_inst_dmem_n16343), .A2(MEM_stage_inst_dmem_n14418), .ZN(MEM_stage_inst_dmem_n14387) );
INV_X1 MEM_stage_inst_dmem_U11204 ( .A(MEM_stage_inst_dmem_n14417), .ZN(MEM_stage_inst_dmem_n14418) );
NAND2_X1 MEM_stage_inst_dmem_U11203 ( .A1(MEM_stage_inst_dmem_ram_735), .A2(MEM_stage_inst_dmem_n14417), .ZN(MEM_stage_inst_dmem_n14388) );
NAND2_X1 MEM_stage_inst_dmem_U11202 ( .A1(MEM_stage_inst_dmem_n21004), .A2(MEM_stage_inst_dmem_n14837), .ZN(MEM_stage_inst_dmem_n14417) );
NAND2_X1 MEM_stage_inst_dmem_U11201 ( .A1(MEM_stage_inst_dmem_n14386), .A2(MEM_stage_inst_dmem_n14385), .ZN(MEM_stage_inst_dmem_n12059) );
NAND2_X1 MEM_stage_inst_dmem_U11200 ( .A1(MEM_stage_inst_dmem_n14732), .A2(MEM_stage_inst_dmem_n14384), .ZN(MEM_stage_inst_dmem_n14385) );
NAND2_X1 MEM_stage_inst_dmem_U11199 ( .A1(MEM_stage_inst_dmem_ram_736), .A2(MEM_stage_inst_dmem_n14383), .ZN(MEM_stage_inst_dmem_n14386) );
NAND2_X1 MEM_stage_inst_dmem_U11198 ( .A1(MEM_stage_inst_dmem_n14382), .A2(MEM_stage_inst_dmem_n14381), .ZN(MEM_stage_inst_dmem_n12060) );
NAND2_X1 MEM_stage_inst_dmem_U11197 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n14384), .ZN(MEM_stage_inst_dmem_n14381) );
NAND2_X1 MEM_stage_inst_dmem_U11196 ( .A1(MEM_stage_inst_dmem_ram_737), .A2(MEM_stage_inst_dmem_n14383), .ZN(MEM_stage_inst_dmem_n14382) );
NAND2_X1 MEM_stage_inst_dmem_U11195 ( .A1(MEM_stage_inst_dmem_n14380), .A2(MEM_stage_inst_dmem_n14379), .ZN(MEM_stage_inst_dmem_n12061) );
NAND2_X1 MEM_stage_inst_dmem_U11194 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n14384), .ZN(MEM_stage_inst_dmem_n14379) );
NAND2_X1 MEM_stage_inst_dmem_U11193 ( .A1(MEM_stage_inst_dmem_ram_738), .A2(MEM_stage_inst_dmem_n14383), .ZN(MEM_stage_inst_dmem_n14380) );
NAND2_X1 MEM_stage_inst_dmem_U11192 ( .A1(MEM_stage_inst_dmem_n14378), .A2(MEM_stage_inst_dmem_n14377), .ZN(MEM_stage_inst_dmem_n12062) );
NAND2_X1 MEM_stage_inst_dmem_U11191 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n14384), .ZN(MEM_stage_inst_dmem_n14377) );
NAND2_X1 MEM_stage_inst_dmem_U11190 ( .A1(MEM_stage_inst_dmem_ram_739), .A2(MEM_stage_inst_dmem_n14383), .ZN(MEM_stage_inst_dmem_n14378) );
NAND2_X1 MEM_stage_inst_dmem_U11189 ( .A1(MEM_stage_inst_dmem_n14376), .A2(MEM_stage_inst_dmem_n14375), .ZN(MEM_stage_inst_dmem_n12063) );
NAND2_X1 MEM_stage_inst_dmem_U11188 ( .A1(MEM_stage_inst_dmem_n16368), .A2(MEM_stage_inst_dmem_n14384), .ZN(MEM_stage_inst_dmem_n14375) );
NAND2_X1 MEM_stage_inst_dmem_U11187 ( .A1(MEM_stage_inst_dmem_ram_740), .A2(MEM_stage_inst_dmem_n14383), .ZN(MEM_stage_inst_dmem_n14376) );
NAND2_X1 MEM_stage_inst_dmem_U11186 ( .A1(MEM_stage_inst_dmem_n14374), .A2(MEM_stage_inst_dmem_n14373), .ZN(MEM_stage_inst_dmem_n12064) );
NAND2_X1 MEM_stage_inst_dmem_U11185 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n14384), .ZN(MEM_stage_inst_dmem_n14373) );
NAND2_X1 MEM_stage_inst_dmem_U11184 ( .A1(MEM_stage_inst_dmem_ram_741), .A2(MEM_stage_inst_dmem_n14383), .ZN(MEM_stage_inst_dmem_n14374) );
NAND2_X1 MEM_stage_inst_dmem_U11183 ( .A1(MEM_stage_inst_dmem_n14372), .A2(MEM_stage_inst_dmem_n14371), .ZN(MEM_stage_inst_dmem_n12065) );
NAND2_X1 MEM_stage_inst_dmem_U11182 ( .A1(MEM_stage_inst_dmem_n14717), .A2(MEM_stage_inst_dmem_n14384), .ZN(MEM_stage_inst_dmem_n14371) );
NAND2_X1 MEM_stage_inst_dmem_U11181 ( .A1(MEM_stage_inst_dmem_ram_742), .A2(MEM_stage_inst_dmem_n14383), .ZN(MEM_stage_inst_dmem_n14372) );
NAND2_X1 MEM_stage_inst_dmem_U11180 ( .A1(MEM_stage_inst_dmem_n14370), .A2(MEM_stage_inst_dmem_n14369), .ZN(MEM_stage_inst_dmem_n12066) );
NAND2_X1 MEM_stage_inst_dmem_U11179 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n14384), .ZN(MEM_stage_inst_dmem_n14369) );
NAND2_X1 MEM_stage_inst_dmem_U11178 ( .A1(MEM_stage_inst_dmem_ram_743), .A2(MEM_stage_inst_dmem_n14383), .ZN(MEM_stage_inst_dmem_n14370) );
NAND2_X1 MEM_stage_inst_dmem_U11177 ( .A1(MEM_stage_inst_dmem_n14368), .A2(MEM_stage_inst_dmem_n14367), .ZN(MEM_stage_inst_dmem_n12067) );
NAND2_X1 MEM_stage_inst_dmem_U11176 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n14384), .ZN(MEM_stage_inst_dmem_n14367) );
NAND2_X1 MEM_stage_inst_dmem_U11175 ( .A1(MEM_stage_inst_dmem_ram_744), .A2(MEM_stage_inst_dmem_n14383), .ZN(MEM_stage_inst_dmem_n14368) );
NAND2_X1 MEM_stage_inst_dmem_U11174 ( .A1(MEM_stage_inst_dmem_n14366), .A2(MEM_stage_inst_dmem_n14365), .ZN(MEM_stage_inst_dmem_n12068) );
NAND2_X1 MEM_stage_inst_dmem_U11173 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n14384), .ZN(MEM_stage_inst_dmem_n14365) );
NAND2_X1 MEM_stage_inst_dmem_U11172 ( .A1(MEM_stage_inst_dmem_ram_745), .A2(MEM_stage_inst_dmem_n14383), .ZN(MEM_stage_inst_dmem_n14366) );
NAND2_X1 MEM_stage_inst_dmem_U11171 ( .A1(MEM_stage_inst_dmem_n14364), .A2(MEM_stage_inst_dmem_n14363), .ZN(MEM_stage_inst_dmem_n12069) );
NAND2_X1 MEM_stage_inst_dmem_U11170 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n14384), .ZN(MEM_stage_inst_dmem_n14363) );
NAND2_X1 MEM_stage_inst_dmem_U11169 ( .A1(MEM_stage_inst_dmem_ram_746), .A2(MEM_stage_inst_dmem_n14383), .ZN(MEM_stage_inst_dmem_n14364) );
NAND2_X1 MEM_stage_inst_dmem_U11168 ( .A1(MEM_stage_inst_dmem_n14362), .A2(MEM_stage_inst_dmem_n14361), .ZN(MEM_stage_inst_dmem_n12070) );
NAND2_X1 MEM_stage_inst_dmem_U11167 ( .A1(MEM_stage_inst_dmem_n14705), .A2(MEM_stage_inst_dmem_n14384), .ZN(MEM_stage_inst_dmem_n14361) );
NAND2_X1 MEM_stage_inst_dmem_U11166 ( .A1(MEM_stage_inst_dmem_ram_747), .A2(MEM_stage_inst_dmem_n14383), .ZN(MEM_stage_inst_dmem_n14362) );
NAND2_X1 MEM_stage_inst_dmem_U11165 ( .A1(MEM_stage_inst_dmem_n14360), .A2(MEM_stage_inst_dmem_n14359), .ZN(MEM_stage_inst_dmem_n12071) );
NAND2_X1 MEM_stage_inst_dmem_U11164 ( .A1(MEM_stage_inst_dmem_n14702), .A2(MEM_stage_inst_dmem_n14384), .ZN(MEM_stage_inst_dmem_n14359) );
NAND2_X1 MEM_stage_inst_dmem_U11163 ( .A1(MEM_stage_inst_dmem_ram_748), .A2(MEM_stage_inst_dmem_n14383), .ZN(MEM_stage_inst_dmem_n14360) );
NAND2_X1 MEM_stage_inst_dmem_U11162 ( .A1(MEM_stage_inst_dmem_n14358), .A2(MEM_stage_inst_dmem_n14357), .ZN(MEM_stage_inst_dmem_n12072) );
NAND2_X1 MEM_stage_inst_dmem_U11161 ( .A1(MEM_stage_inst_dmem_n116), .A2(MEM_stage_inst_dmem_n14384), .ZN(MEM_stage_inst_dmem_n14357) );
NAND2_X1 MEM_stage_inst_dmem_U11160 ( .A1(MEM_stage_inst_dmem_ram_749), .A2(MEM_stage_inst_dmem_n14383), .ZN(MEM_stage_inst_dmem_n14358) );
NAND2_X1 MEM_stage_inst_dmem_U11159 ( .A1(MEM_stage_inst_dmem_n14356), .A2(MEM_stage_inst_dmem_n14355), .ZN(MEM_stage_inst_dmem_n12073) );
NAND2_X1 MEM_stage_inst_dmem_U11158 ( .A1(MEM_stage_inst_dmem_n14696), .A2(MEM_stage_inst_dmem_n14384), .ZN(MEM_stage_inst_dmem_n14355) );
NAND2_X1 MEM_stage_inst_dmem_U11157 ( .A1(MEM_stage_inst_dmem_ram_750), .A2(MEM_stage_inst_dmem_n14383), .ZN(MEM_stage_inst_dmem_n14356) );
NAND2_X1 MEM_stage_inst_dmem_U11156 ( .A1(MEM_stage_inst_dmem_n14354), .A2(MEM_stage_inst_dmem_n14353), .ZN(MEM_stage_inst_dmem_n12074) );
NAND2_X1 MEM_stage_inst_dmem_U11155 ( .A1(MEM_stage_inst_dmem_n14693), .A2(MEM_stage_inst_dmem_n14384), .ZN(MEM_stage_inst_dmem_n14353) );
INV_X1 MEM_stage_inst_dmem_U11154 ( .A(MEM_stage_inst_dmem_n14383), .ZN(MEM_stage_inst_dmem_n14384) );
NAND2_X1 MEM_stage_inst_dmem_U11153 ( .A1(MEM_stage_inst_dmem_ram_751), .A2(MEM_stage_inst_dmem_n14383), .ZN(MEM_stage_inst_dmem_n14354) );
NAND2_X1 MEM_stage_inst_dmem_U11152 ( .A1(MEM_stage_inst_dmem_n20969), .A2(MEM_stage_inst_dmem_n14837), .ZN(MEM_stage_inst_dmem_n14383) );
NAND2_X1 MEM_stage_inst_dmem_U11151 ( .A1(MEM_stage_inst_dmem_n14352), .A2(MEM_stage_inst_dmem_n14351), .ZN(MEM_stage_inst_dmem_n12075) );
NAND2_X1 MEM_stage_inst_dmem_U11150 ( .A1(MEM_stage_inst_dmem_n14732), .A2(MEM_stage_inst_dmem_n14350), .ZN(MEM_stage_inst_dmem_n14351) );
BUF_X1 MEM_stage_inst_dmem_U11149 ( .A(EX_pipeline_reg_out_5), .Z(MEM_stage_inst_dmem_n20551) );
NAND2_X1 MEM_stage_inst_dmem_U11148 ( .A1(MEM_stage_inst_dmem_ram_752), .A2(MEM_stage_inst_dmem_n14349), .ZN(MEM_stage_inst_dmem_n14352) );
NAND2_X1 MEM_stage_inst_dmem_U11147 ( .A1(MEM_stage_inst_dmem_n14348), .A2(MEM_stage_inst_dmem_n14347), .ZN(MEM_stage_inst_dmem_n12076) );
NAND2_X1 MEM_stage_inst_dmem_U11146 ( .A1(MEM_stage_inst_dmem_n20547), .A2(MEM_stage_inst_dmem_n14350), .ZN(MEM_stage_inst_dmem_n14347) );
BUF_X1 MEM_stage_inst_dmem_U11145 ( .A(EX_pipeline_reg_out_6), .Z(MEM_stage_inst_dmem_n20547) );
NAND2_X1 MEM_stage_inst_dmem_U11144 ( .A1(MEM_stage_inst_dmem_ram_753), .A2(MEM_stage_inst_dmem_n14349), .ZN(MEM_stage_inst_dmem_n14348) );
NAND2_X1 MEM_stage_inst_dmem_U11143 ( .A1(MEM_stage_inst_dmem_n14346), .A2(MEM_stage_inst_dmem_n14345), .ZN(MEM_stage_inst_dmem_n12077) );
NAND2_X1 MEM_stage_inst_dmem_U11142 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n14350), .ZN(MEM_stage_inst_dmem_n14345) );
BUF_X1 MEM_stage_inst_dmem_U11141 ( .A(EX_pipeline_reg_out_7), .Z(MEM_stage_inst_dmem_n20544) );
NAND2_X1 MEM_stage_inst_dmem_U11140 ( .A1(MEM_stage_inst_dmem_ram_754), .A2(MEM_stage_inst_dmem_n14349), .ZN(MEM_stage_inst_dmem_n14346) );
NAND2_X1 MEM_stage_inst_dmem_U11139 ( .A1(MEM_stage_inst_dmem_n14344), .A2(MEM_stage_inst_dmem_n14343), .ZN(MEM_stage_inst_dmem_n12078) );
NAND2_X1 MEM_stage_inst_dmem_U11138 ( .A1(MEM_stage_inst_dmem_n20541), .A2(MEM_stage_inst_dmem_n14350), .ZN(MEM_stage_inst_dmem_n14343) );
NAND2_X1 MEM_stage_inst_dmem_U11137 ( .A1(MEM_stage_inst_dmem_ram_755), .A2(MEM_stage_inst_dmem_n14349), .ZN(MEM_stage_inst_dmem_n14344) );
NAND2_X1 MEM_stage_inst_dmem_U11136 ( .A1(MEM_stage_inst_dmem_n14342), .A2(MEM_stage_inst_dmem_n14341), .ZN(MEM_stage_inst_dmem_n12079) );
NAND2_X1 MEM_stage_inst_dmem_U11135 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n14350), .ZN(MEM_stage_inst_dmem_n14341) );
NAND2_X1 MEM_stage_inst_dmem_U11134 ( .A1(MEM_stage_inst_dmem_ram_756), .A2(MEM_stage_inst_dmem_n14349), .ZN(MEM_stage_inst_dmem_n14342) );
NAND2_X1 MEM_stage_inst_dmem_U11133 ( .A1(MEM_stage_inst_dmem_n14340), .A2(MEM_stage_inst_dmem_n14339), .ZN(MEM_stage_inst_dmem_n12080) );
NAND2_X1 MEM_stage_inst_dmem_U11132 ( .A1(MEM_stage_inst_dmem_n20536), .A2(MEM_stage_inst_dmem_n14350), .ZN(MEM_stage_inst_dmem_n14339) );
NAND2_X1 MEM_stage_inst_dmem_U11131 ( .A1(MEM_stage_inst_dmem_ram_757), .A2(MEM_stage_inst_dmem_n14349), .ZN(MEM_stage_inst_dmem_n14340) );
NAND2_X1 MEM_stage_inst_dmem_U11130 ( .A1(MEM_stage_inst_dmem_n14338), .A2(MEM_stage_inst_dmem_n14337), .ZN(MEM_stage_inst_dmem_n12081) );
NAND2_X1 MEM_stage_inst_dmem_U11129 ( .A1(MEM_stage_inst_dmem_n14717), .A2(MEM_stage_inst_dmem_n14350), .ZN(MEM_stage_inst_dmem_n14337) );
NAND2_X1 MEM_stage_inst_dmem_U11128 ( .A1(MEM_stage_inst_dmem_ram_758), .A2(MEM_stage_inst_dmem_n14349), .ZN(MEM_stage_inst_dmem_n14338) );
NAND2_X1 MEM_stage_inst_dmem_U11127 ( .A1(MEM_stage_inst_dmem_n14336), .A2(MEM_stage_inst_dmem_n14335), .ZN(MEM_stage_inst_dmem_n12082) );
NAND2_X1 MEM_stage_inst_dmem_U11126 ( .A1(MEM_stage_inst_dmem_n16361), .A2(MEM_stage_inst_dmem_n14350), .ZN(MEM_stage_inst_dmem_n14335) );
BUF_X1 MEM_stage_inst_dmem_U11125 ( .A(EX_pipeline_reg_out_12), .Z(MEM_stage_inst_dmem_n20530) );
NAND2_X1 MEM_stage_inst_dmem_U11124 ( .A1(MEM_stage_inst_dmem_ram_759), .A2(MEM_stage_inst_dmem_n14349), .ZN(MEM_stage_inst_dmem_n14336) );
NAND2_X1 MEM_stage_inst_dmem_U11123 ( .A1(MEM_stage_inst_dmem_n14334), .A2(MEM_stage_inst_dmem_n14333), .ZN(MEM_stage_inst_dmem_n12083) );
NAND2_X1 MEM_stage_inst_dmem_U11122 ( .A1(MEM_stage_inst_dmem_n104), .A2(MEM_stage_inst_dmem_n14350), .ZN(MEM_stage_inst_dmem_n14333) );
BUF_X1 MEM_stage_inst_dmem_U11121 ( .A(EX_pipeline_reg_out_13), .Z(MEM_stage_inst_dmem_n20527) );
NAND2_X1 MEM_stage_inst_dmem_U11120 ( .A1(MEM_stage_inst_dmem_ram_760), .A2(MEM_stage_inst_dmem_n14349), .ZN(MEM_stage_inst_dmem_n14334) );
NAND2_X1 MEM_stage_inst_dmem_U11119 ( .A1(MEM_stage_inst_dmem_n14332), .A2(MEM_stage_inst_dmem_n14331), .ZN(MEM_stage_inst_dmem_n12084) );
NAND2_X1 MEM_stage_inst_dmem_U11118 ( .A1(EX_pipeline_reg_out_14), .A2(MEM_stage_inst_dmem_n14350), .ZN(MEM_stage_inst_dmem_n14331) );
BUF_X1 MEM_stage_inst_dmem_U11117 ( .A(EX_pipeline_reg_out_14), .Z(MEM_stage_inst_dmem_n20524) );
NAND2_X1 MEM_stage_inst_dmem_U11116 ( .A1(MEM_stage_inst_dmem_ram_761), .A2(MEM_stage_inst_dmem_n14349), .ZN(MEM_stage_inst_dmem_n14332) );
NAND2_X1 MEM_stage_inst_dmem_U11115 ( .A1(MEM_stage_inst_dmem_n14330), .A2(MEM_stage_inst_dmem_n14329), .ZN(MEM_stage_inst_dmem_n12085) );
NAND2_X1 MEM_stage_inst_dmem_U11114 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n14350), .ZN(MEM_stage_inst_dmem_n14329) );
BUF_X1 MEM_stage_inst_dmem_U11113 ( .A(EX_pipeline_reg_out_15), .Z(MEM_stage_inst_dmem_n20521) );
NAND2_X1 MEM_stage_inst_dmem_U11112 ( .A1(MEM_stage_inst_dmem_ram_762), .A2(MEM_stage_inst_dmem_n14349), .ZN(MEM_stage_inst_dmem_n14330) );
NAND2_X1 MEM_stage_inst_dmem_U11111 ( .A1(MEM_stage_inst_dmem_n14328), .A2(MEM_stage_inst_dmem_n14327), .ZN(MEM_stage_inst_dmem_n12086) );
NAND2_X1 MEM_stage_inst_dmem_U11110 ( .A1(MEM_stage_inst_dmem_n103), .A2(MEM_stage_inst_dmem_n14350), .ZN(MEM_stage_inst_dmem_n14327) );
BUF_X1 MEM_stage_inst_dmem_U11109 ( .A(EX_pipeline_reg_out_16), .Z(MEM_stage_inst_dmem_n20518) );
NAND2_X1 MEM_stage_inst_dmem_U11108 ( .A1(MEM_stage_inst_dmem_ram_763), .A2(MEM_stage_inst_dmem_n14349), .ZN(MEM_stage_inst_dmem_n14328) );
NAND2_X1 MEM_stage_inst_dmem_U11107 ( .A1(MEM_stage_inst_dmem_n14326), .A2(MEM_stage_inst_dmem_n14325), .ZN(MEM_stage_inst_dmem_n12087) );
NAND2_X1 MEM_stage_inst_dmem_U11106 ( .A1(MEM_stage_inst_dmem_n105), .A2(MEM_stage_inst_dmem_n14350), .ZN(MEM_stage_inst_dmem_n14325) );
BUF_X1 MEM_stage_inst_dmem_U11105 ( .A(EX_pipeline_reg_out_17), .Z(MEM_stage_inst_dmem_n20515) );
NAND2_X1 MEM_stage_inst_dmem_U11104 ( .A1(MEM_stage_inst_dmem_ram_764), .A2(MEM_stage_inst_dmem_n14349), .ZN(MEM_stage_inst_dmem_n14326) );
NAND2_X1 MEM_stage_inst_dmem_U11103 ( .A1(MEM_stage_inst_dmem_n14324), .A2(MEM_stage_inst_dmem_n14323), .ZN(MEM_stage_inst_dmem_n12088) );
NAND2_X1 MEM_stage_inst_dmem_U11102 ( .A1(MEM_stage_inst_dmem_n116), .A2(MEM_stage_inst_dmem_n14350), .ZN(MEM_stage_inst_dmem_n14323) );
BUF_X1 MEM_stage_inst_dmem_U11101 ( .A(EX_pipeline_reg_out_18), .Z(MEM_stage_inst_dmem_n20512) );
NAND2_X1 MEM_stage_inst_dmem_U11100 ( .A1(MEM_stage_inst_dmem_ram_765), .A2(MEM_stage_inst_dmem_n14349), .ZN(MEM_stage_inst_dmem_n14324) );
NAND2_X1 MEM_stage_inst_dmem_U11099 ( .A1(MEM_stage_inst_dmem_n14322), .A2(MEM_stage_inst_dmem_n14321), .ZN(MEM_stage_inst_dmem_n12089) );
NAND2_X1 MEM_stage_inst_dmem_U11098 ( .A1(MEM_stage_inst_dmem_n14696), .A2(MEM_stage_inst_dmem_n14350), .ZN(MEM_stage_inst_dmem_n14321) );
BUF_X1 MEM_stage_inst_dmem_U11097 ( .A(EX_pipeline_reg_out_19), .Z(MEM_stage_inst_dmem_n20509) );
NAND2_X1 MEM_stage_inst_dmem_U11096 ( .A1(MEM_stage_inst_dmem_ram_766), .A2(MEM_stage_inst_dmem_n14349), .ZN(MEM_stage_inst_dmem_n14322) );
NAND2_X1 MEM_stage_inst_dmem_U11095 ( .A1(MEM_stage_inst_dmem_n14320), .A2(MEM_stage_inst_dmem_n14319), .ZN(MEM_stage_inst_dmem_n12090) );
NAND2_X1 MEM_stage_inst_dmem_U11094 ( .A1(MEM_stage_inst_dmem_n15110), .A2(MEM_stage_inst_dmem_n14350), .ZN(MEM_stage_inst_dmem_n14319) );
INV_X1 MEM_stage_inst_dmem_U11093 ( .A(MEM_stage_inst_dmem_n14349), .ZN(MEM_stage_inst_dmem_n14350) );
BUF_X1 MEM_stage_inst_dmem_U11092 ( .A(EX_pipeline_reg_out_20), .Z(MEM_stage_inst_dmem_n20506) );
NAND2_X1 MEM_stage_inst_dmem_U11091 ( .A1(MEM_stage_inst_dmem_ram_767), .A2(MEM_stage_inst_dmem_n14349), .ZN(MEM_stage_inst_dmem_n14320) );
NAND2_X1 MEM_stage_inst_dmem_U11090 ( .A1(MEM_stage_inst_dmem_n20934), .A2(MEM_stage_inst_dmem_n14837), .ZN(MEM_stage_inst_dmem_n14349) );
NOR2_X2 MEM_stage_inst_dmem_U11089 ( .A1(MEM_stage_inst_dmem_n16519), .A2(MEM_stage_inst_dmem_n18718), .ZN(MEM_stage_inst_dmem_n14837) );
NAND2_X1 MEM_stage_inst_dmem_U11088 ( .A1(MEM_stage_inst_dmem_n14318), .A2(MEM_stage_inst_dmem_n14317), .ZN(MEM_stage_inst_dmem_n12091) );
NAND2_X1 MEM_stage_inst_dmem_U11087 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n14316), .ZN(MEM_stage_inst_dmem_n14317) );
NAND2_X1 MEM_stage_inst_dmem_U11086 ( .A1(MEM_stage_inst_dmem_ram_768), .A2(MEM_stage_inst_dmem_n14315), .ZN(MEM_stage_inst_dmem_n14318) );
NAND2_X1 MEM_stage_inst_dmem_U11085 ( .A1(MEM_stage_inst_dmem_n14314), .A2(MEM_stage_inst_dmem_n14313), .ZN(MEM_stage_inst_dmem_n12092) );
NAND2_X1 MEM_stage_inst_dmem_U11084 ( .A1(EX_pipeline_reg_out_6), .A2(MEM_stage_inst_dmem_n14316), .ZN(MEM_stage_inst_dmem_n14313) );
NAND2_X1 MEM_stage_inst_dmem_U11083 ( .A1(MEM_stage_inst_dmem_ram_769), .A2(MEM_stage_inst_dmem_n14315), .ZN(MEM_stage_inst_dmem_n14314) );
NAND2_X1 MEM_stage_inst_dmem_U11082 ( .A1(MEM_stage_inst_dmem_n14312), .A2(MEM_stage_inst_dmem_n14311), .ZN(MEM_stage_inst_dmem_n12093) );
NAND2_X1 MEM_stage_inst_dmem_U11081 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n14316), .ZN(MEM_stage_inst_dmem_n14311) );
NAND2_X1 MEM_stage_inst_dmem_U11080 ( .A1(MEM_stage_inst_dmem_ram_770), .A2(MEM_stage_inst_dmem_n14315), .ZN(MEM_stage_inst_dmem_n14312) );
NAND2_X1 MEM_stage_inst_dmem_U11079 ( .A1(MEM_stage_inst_dmem_n14310), .A2(MEM_stage_inst_dmem_n14309), .ZN(MEM_stage_inst_dmem_n12094) );
NAND2_X1 MEM_stage_inst_dmem_U11078 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n14316), .ZN(MEM_stage_inst_dmem_n14309) );
NAND2_X1 MEM_stage_inst_dmem_U11077 ( .A1(MEM_stage_inst_dmem_ram_771), .A2(MEM_stage_inst_dmem_n14315), .ZN(MEM_stage_inst_dmem_n14310) );
NAND2_X1 MEM_stage_inst_dmem_U11076 ( .A1(MEM_stage_inst_dmem_n14308), .A2(MEM_stage_inst_dmem_n14307), .ZN(MEM_stage_inst_dmem_n12095) );
NAND2_X1 MEM_stage_inst_dmem_U11075 ( .A1(EX_pipeline_reg_out_9), .A2(MEM_stage_inst_dmem_n14316), .ZN(MEM_stage_inst_dmem_n14307) );
NAND2_X1 MEM_stage_inst_dmem_U11074 ( .A1(MEM_stage_inst_dmem_ram_772), .A2(MEM_stage_inst_dmem_n14315), .ZN(MEM_stage_inst_dmem_n14308) );
NAND2_X1 MEM_stage_inst_dmem_U11073 ( .A1(MEM_stage_inst_dmem_n14306), .A2(MEM_stage_inst_dmem_n14305), .ZN(MEM_stage_inst_dmem_n12096) );
NAND2_X1 MEM_stage_inst_dmem_U11072 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n14316), .ZN(MEM_stage_inst_dmem_n14305) );
NAND2_X1 MEM_stage_inst_dmem_U11071 ( .A1(MEM_stage_inst_dmem_ram_773), .A2(MEM_stage_inst_dmem_n14315), .ZN(MEM_stage_inst_dmem_n14306) );
NAND2_X1 MEM_stage_inst_dmem_U11070 ( .A1(MEM_stage_inst_dmem_n14304), .A2(MEM_stage_inst_dmem_n14303), .ZN(MEM_stage_inst_dmem_n12097) );
NAND2_X1 MEM_stage_inst_dmem_U11069 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n14316), .ZN(MEM_stage_inst_dmem_n14303) );
NAND2_X1 MEM_stage_inst_dmem_U11068 ( .A1(MEM_stage_inst_dmem_ram_774), .A2(MEM_stage_inst_dmem_n14315), .ZN(MEM_stage_inst_dmem_n14304) );
NAND2_X1 MEM_stage_inst_dmem_U11067 ( .A1(MEM_stage_inst_dmem_n14302), .A2(MEM_stage_inst_dmem_n14301), .ZN(MEM_stage_inst_dmem_n12098) );
NAND2_X1 MEM_stage_inst_dmem_U11066 ( .A1(MEM_stage_inst_dmem_n17), .A2(MEM_stage_inst_dmem_n14316), .ZN(MEM_stage_inst_dmem_n14301) );
NAND2_X1 MEM_stage_inst_dmem_U11065 ( .A1(MEM_stage_inst_dmem_ram_775), .A2(MEM_stage_inst_dmem_n14315), .ZN(MEM_stage_inst_dmem_n14302) );
NAND2_X1 MEM_stage_inst_dmem_U11064 ( .A1(MEM_stage_inst_dmem_n14300), .A2(MEM_stage_inst_dmem_n14299), .ZN(MEM_stage_inst_dmem_n12099) );
NAND2_X1 MEM_stage_inst_dmem_U11063 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n14316), .ZN(MEM_stage_inst_dmem_n14299) );
NAND2_X1 MEM_stage_inst_dmem_U11062 ( .A1(MEM_stage_inst_dmem_ram_776), .A2(MEM_stage_inst_dmem_n14315), .ZN(MEM_stage_inst_dmem_n14300) );
NAND2_X1 MEM_stage_inst_dmem_U11061 ( .A1(MEM_stage_inst_dmem_n14298), .A2(MEM_stage_inst_dmem_n14297), .ZN(MEM_stage_inst_dmem_n12100) );
NAND2_X1 MEM_stage_inst_dmem_U11060 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n14316), .ZN(MEM_stage_inst_dmem_n14297) );
NAND2_X1 MEM_stage_inst_dmem_U11059 ( .A1(MEM_stage_inst_dmem_ram_777), .A2(MEM_stage_inst_dmem_n14315), .ZN(MEM_stage_inst_dmem_n14298) );
NAND2_X1 MEM_stage_inst_dmem_U11058 ( .A1(MEM_stage_inst_dmem_n14296), .A2(MEM_stage_inst_dmem_n14295), .ZN(MEM_stage_inst_dmem_n12101) );
NAND2_X1 MEM_stage_inst_dmem_U11057 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n14316), .ZN(MEM_stage_inst_dmem_n14295) );
NAND2_X1 MEM_stage_inst_dmem_U11056 ( .A1(MEM_stage_inst_dmem_ram_778), .A2(MEM_stage_inst_dmem_n14315), .ZN(MEM_stage_inst_dmem_n14296) );
NAND2_X1 MEM_stage_inst_dmem_U11055 ( .A1(MEM_stage_inst_dmem_n14294), .A2(MEM_stage_inst_dmem_n14293), .ZN(MEM_stage_inst_dmem_n12102) );
NAND2_X1 MEM_stage_inst_dmem_U11054 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n14316), .ZN(MEM_stage_inst_dmem_n14293) );
NAND2_X1 MEM_stage_inst_dmem_U11053 ( .A1(MEM_stage_inst_dmem_ram_779), .A2(MEM_stage_inst_dmem_n14315), .ZN(MEM_stage_inst_dmem_n14294) );
NAND2_X1 MEM_stage_inst_dmem_U11052 ( .A1(MEM_stage_inst_dmem_n14292), .A2(MEM_stage_inst_dmem_n14291), .ZN(MEM_stage_inst_dmem_n12103) );
NAND2_X1 MEM_stage_inst_dmem_U11051 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n14316), .ZN(MEM_stage_inst_dmem_n14291) );
NAND2_X1 MEM_stage_inst_dmem_U11050 ( .A1(MEM_stage_inst_dmem_ram_780), .A2(MEM_stage_inst_dmem_n14315), .ZN(MEM_stage_inst_dmem_n14292) );
NAND2_X1 MEM_stage_inst_dmem_U11049 ( .A1(MEM_stage_inst_dmem_n14290), .A2(MEM_stage_inst_dmem_n14289), .ZN(MEM_stage_inst_dmem_n12104) );
NAND2_X1 MEM_stage_inst_dmem_U11048 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n14316), .ZN(MEM_stage_inst_dmem_n14289) );
NAND2_X1 MEM_stage_inst_dmem_U11047 ( .A1(MEM_stage_inst_dmem_ram_781), .A2(MEM_stage_inst_dmem_n14315), .ZN(MEM_stage_inst_dmem_n14290) );
NAND2_X1 MEM_stage_inst_dmem_U11046 ( .A1(MEM_stage_inst_dmem_n14288), .A2(MEM_stage_inst_dmem_n14287), .ZN(MEM_stage_inst_dmem_n12105) );
NAND2_X1 MEM_stage_inst_dmem_U11045 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n14316), .ZN(MEM_stage_inst_dmem_n14287) );
NAND2_X1 MEM_stage_inst_dmem_U11044 ( .A1(MEM_stage_inst_dmem_ram_782), .A2(MEM_stage_inst_dmem_n14315), .ZN(MEM_stage_inst_dmem_n14288) );
NAND2_X1 MEM_stage_inst_dmem_U11043 ( .A1(MEM_stage_inst_dmem_n14286), .A2(MEM_stage_inst_dmem_n14285), .ZN(MEM_stage_inst_dmem_n12106) );
NAND2_X1 MEM_stage_inst_dmem_U11042 ( .A1(MEM_stage_inst_dmem_n15110), .A2(MEM_stage_inst_dmem_n14316), .ZN(MEM_stage_inst_dmem_n14285) );
INV_X1 MEM_stage_inst_dmem_U11041 ( .A(MEM_stage_inst_dmem_n14315), .ZN(MEM_stage_inst_dmem_n14316) );
NAND2_X1 MEM_stage_inst_dmem_U11040 ( .A1(MEM_stage_inst_dmem_ram_783), .A2(MEM_stage_inst_dmem_n14315), .ZN(MEM_stage_inst_dmem_n14286) );
NAND2_X1 MEM_stage_inst_dmem_U11039 ( .A1(MEM_stage_inst_dmem_n21465), .A2(MEM_stage_inst_dmem_n14284), .ZN(MEM_stage_inst_dmem_n14315) );
NAND2_X1 MEM_stage_inst_dmem_U11038 ( .A1(MEM_stage_inst_dmem_n14283), .A2(MEM_stage_inst_dmem_n14282), .ZN(MEM_stage_inst_dmem_n12107) );
NAND2_X1 MEM_stage_inst_dmem_U11037 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n14281), .ZN(MEM_stage_inst_dmem_n14282) );
NAND2_X1 MEM_stage_inst_dmem_U11036 ( .A1(MEM_stage_inst_dmem_ram_784), .A2(MEM_stage_inst_dmem_n14280), .ZN(MEM_stage_inst_dmem_n14283) );
NAND2_X1 MEM_stage_inst_dmem_U11035 ( .A1(MEM_stage_inst_dmem_n14279), .A2(MEM_stage_inst_dmem_n14278), .ZN(MEM_stage_inst_dmem_n12108) );
NAND2_X1 MEM_stage_inst_dmem_U11034 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n14281), .ZN(MEM_stage_inst_dmem_n14278) );
NAND2_X1 MEM_stage_inst_dmem_U11033 ( .A1(MEM_stage_inst_dmem_ram_785), .A2(MEM_stage_inst_dmem_n14280), .ZN(MEM_stage_inst_dmem_n14279) );
NAND2_X1 MEM_stage_inst_dmem_U11032 ( .A1(MEM_stage_inst_dmem_n14277), .A2(MEM_stage_inst_dmem_n14276), .ZN(MEM_stage_inst_dmem_n12109) );
NAND2_X1 MEM_stage_inst_dmem_U11031 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n14281), .ZN(MEM_stage_inst_dmem_n14276) );
NAND2_X1 MEM_stage_inst_dmem_U11030 ( .A1(MEM_stage_inst_dmem_ram_786), .A2(MEM_stage_inst_dmem_n14280), .ZN(MEM_stage_inst_dmem_n14277) );
NAND2_X1 MEM_stage_inst_dmem_U11029 ( .A1(MEM_stage_inst_dmem_n14275), .A2(MEM_stage_inst_dmem_n14274), .ZN(MEM_stage_inst_dmem_n12110) );
NAND2_X1 MEM_stage_inst_dmem_U11028 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n14281), .ZN(MEM_stage_inst_dmem_n14274) );
NAND2_X1 MEM_stage_inst_dmem_U11027 ( .A1(MEM_stage_inst_dmem_ram_787), .A2(MEM_stage_inst_dmem_n14280), .ZN(MEM_stage_inst_dmem_n14275) );
NAND2_X1 MEM_stage_inst_dmem_U11026 ( .A1(MEM_stage_inst_dmem_n14273), .A2(MEM_stage_inst_dmem_n14272), .ZN(MEM_stage_inst_dmem_n12111) );
NAND2_X1 MEM_stage_inst_dmem_U11025 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n14281), .ZN(MEM_stage_inst_dmem_n14272) );
NAND2_X1 MEM_stage_inst_dmem_U11024 ( .A1(MEM_stage_inst_dmem_ram_788), .A2(MEM_stage_inst_dmem_n14280), .ZN(MEM_stage_inst_dmem_n14273) );
NAND2_X1 MEM_stage_inst_dmem_U11023 ( .A1(MEM_stage_inst_dmem_n14271), .A2(MEM_stage_inst_dmem_n14270), .ZN(MEM_stage_inst_dmem_n12112) );
NAND2_X1 MEM_stage_inst_dmem_U11022 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n14281), .ZN(MEM_stage_inst_dmem_n14270) );
NAND2_X1 MEM_stage_inst_dmem_U11021 ( .A1(MEM_stage_inst_dmem_ram_789), .A2(MEM_stage_inst_dmem_n14280), .ZN(MEM_stage_inst_dmem_n14271) );
NAND2_X1 MEM_stage_inst_dmem_U11020 ( .A1(MEM_stage_inst_dmem_n14269), .A2(MEM_stage_inst_dmem_n14268), .ZN(MEM_stage_inst_dmem_n12113) );
NAND2_X1 MEM_stage_inst_dmem_U11019 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n14281), .ZN(MEM_stage_inst_dmem_n14268) );
NAND2_X1 MEM_stage_inst_dmem_U11018 ( .A1(MEM_stage_inst_dmem_ram_790), .A2(MEM_stage_inst_dmem_n14280), .ZN(MEM_stage_inst_dmem_n14269) );
NAND2_X1 MEM_stage_inst_dmem_U11017 ( .A1(MEM_stage_inst_dmem_n14267), .A2(MEM_stage_inst_dmem_n14266), .ZN(MEM_stage_inst_dmem_n12114) );
NAND2_X1 MEM_stage_inst_dmem_U11016 ( .A1(MEM_stage_inst_dmem_n18), .A2(MEM_stage_inst_dmem_n14281), .ZN(MEM_stage_inst_dmem_n14266) );
NAND2_X1 MEM_stage_inst_dmem_U11015 ( .A1(MEM_stage_inst_dmem_ram_791), .A2(MEM_stage_inst_dmem_n14280), .ZN(MEM_stage_inst_dmem_n14267) );
NAND2_X1 MEM_stage_inst_dmem_U11014 ( .A1(MEM_stage_inst_dmem_n14265), .A2(MEM_stage_inst_dmem_n14264), .ZN(MEM_stage_inst_dmem_n12115) );
NAND2_X1 MEM_stage_inst_dmem_U11013 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n14281), .ZN(MEM_stage_inst_dmem_n14264) );
NAND2_X1 MEM_stage_inst_dmem_U11012 ( .A1(MEM_stage_inst_dmem_ram_792), .A2(MEM_stage_inst_dmem_n14280), .ZN(MEM_stage_inst_dmem_n14265) );
NAND2_X1 MEM_stage_inst_dmem_U11011 ( .A1(MEM_stage_inst_dmem_n14263), .A2(MEM_stage_inst_dmem_n14262), .ZN(MEM_stage_inst_dmem_n12116) );
NAND2_X1 MEM_stage_inst_dmem_U11010 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n14281), .ZN(MEM_stage_inst_dmem_n14262) );
NAND2_X1 MEM_stage_inst_dmem_U11009 ( .A1(MEM_stage_inst_dmem_ram_793), .A2(MEM_stage_inst_dmem_n14280), .ZN(MEM_stage_inst_dmem_n14263) );
NAND2_X1 MEM_stage_inst_dmem_U11008 ( .A1(MEM_stage_inst_dmem_n14261), .A2(MEM_stage_inst_dmem_n14260), .ZN(MEM_stage_inst_dmem_n12117) );
NAND2_X1 MEM_stage_inst_dmem_U11007 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n14281), .ZN(MEM_stage_inst_dmem_n14260) );
NAND2_X1 MEM_stage_inst_dmem_U11006 ( .A1(MEM_stage_inst_dmem_ram_794), .A2(MEM_stage_inst_dmem_n14280), .ZN(MEM_stage_inst_dmem_n14261) );
NAND2_X1 MEM_stage_inst_dmem_U11005 ( .A1(MEM_stage_inst_dmem_n14259), .A2(MEM_stage_inst_dmem_n14258), .ZN(MEM_stage_inst_dmem_n12118) );
NAND2_X1 MEM_stage_inst_dmem_U11004 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n14281), .ZN(MEM_stage_inst_dmem_n14258) );
NAND2_X1 MEM_stage_inst_dmem_U11003 ( .A1(MEM_stage_inst_dmem_ram_795), .A2(MEM_stage_inst_dmem_n14280), .ZN(MEM_stage_inst_dmem_n14259) );
NAND2_X1 MEM_stage_inst_dmem_U11002 ( .A1(MEM_stage_inst_dmem_n14257), .A2(MEM_stage_inst_dmem_n14256), .ZN(MEM_stage_inst_dmem_n12119) );
NAND2_X1 MEM_stage_inst_dmem_U11001 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n14281), .ZN(MEM_stage_inst_dmem_n14256) );
NAND2_X1 MEM_stage_inst_dmem_U11000 ( .A1(MEM_stage_inst_dmem_ram_796), .A2(MEM_stage_inst_dmem_n14280), .ZN(MEM_stage_inst_dmem_n14257) );
NAND2_X1 MEM_stage_inst_dmem_U10999 ( .A1(MEM_stage_inst_dmem_n14255), .A2(MEM_stage_inst_dmem_n14254), .ZN(MEM_stage_inst_dmem_n12120) );
NAND2_X1 MEM_stage_inst_dmem_U10998 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n14281), .ZN(MEM_stage_inst_dmem_n14254) );
NAND2_X1 MEM_stage_inst_dmem_U10997 ( .A1(MEM_stage_inst_dmem_ram_797), .A2(MEM_stage_inst_dmem_n14280), .ZN(MEM_stage_inst_dmem_n14255) );
NAND2_X1 MEM_stage_inst_dmem_U10996 ( .A1(MEM_stage_inst_dmem_n14253), .A2(MEM_stage_inst_dmem_n14252), .ZN(MEM_stage_inst_dmem_n12121) );
NAND2_X1 MEM_stage_inst_dmem_U10995 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n14281), .ZN(MEM_stage_inst_dmem_n14252) );
NAND2_X1 MEM_stage_inst_dmem_U10994 ( .A1(MEM_stage_inst_dmem_ram_798), .A2(MEM_stage_inst_dmem_n14280), .ZN(MEM_stage_inst_dmem_n14253) );
NAND2_X1 MEM_stage_inst_dmem_U10993 ( .A1(MEM_stage_inst_dmem_n14251), .A2(MEM_stage_inst_dmem_n14250), .ZN(MEM_stage_inst_dmem_n12122) );
NAND2_X1 MEM_stage_inst_dmem_U10992 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n14281), .ZN(MEM_stage_inst_dmem_n14250) );
INV_X1 MEM_stage_inst_dmem_U10991 ( .A(MEM_stage_inst_dmem_n14280), .ZN(MEM_stage_inst_dmem_n14281) );
NAND2_X1 MEM_stage_inst_dmem_U10990 ( .A1(MEM_stage_inst_dmem_ram_799), .A2(MEM_stage_inst_dmem_n14280), .ZN(MEM_stage_inst_dmem_n14251) );
NAND2_X1 MEM_stage_inst_dmem_U10989 ( .A1(MEM_stage_inst_dmem_n21429), .A2(MEM_stage_inst_dmem_n14284), .ZN(MEM_stage_inst_dmem_n14280) );
NAND2_X1 MEM_stage_inst_dmem_U10988 ( .A1(MEM_stage_inst_dmem_n14249), .A2(MEM_stage_inst_dmem_n14248), .ZN(MEM_stage_inst_dmem_n12123) );
NAND2_X1 MEM_stage_inst_dmem_U10987 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n14247), .ZN(MEM_stage_inst_dmem_n14248) );
NAND2_X1 MEM_stage_inst_dmem_U10986 ( .A1(MEM_stage_inst_dmem_ram_800), .A2(MEM_stage_inst_dmem_n14246), .ZN(MEM_stage_inst_dmem_n14249) );
NAND2_X1 MEM_stage_inst_dmem_U10985 ( .A1(MEM_stage_inst_dmem_n14245), .A2(MEM_stage_inst_dmem_n14244), .ZN(MEM_stage_inst_dmem_n12124) );
NAND2_X1 MEM_stage_inst_dmem_U10984 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n14247), .ZN(MEM_stage_inst_dmem_n14244) );
NAND2_X1 MEM_stage_inst_dmem_U10983 ( .A1(MEM_stage_inst_dmem_ram_801), .A2(MEM_stage_inst_dmem_n14246), .ZN(MEM_stage_inst_dmem_n14245) );
NAND2_X1 MEM_stage_inst_dmem_U10982 ( .A1(MEM_stage_inst_dmem_n14243), .A2(MEM_stage_inst_dmem_n14242), .ZN(MEM_stage_inst_dmem_n12125) );
NAND2_X1 MEM_stage_inst_dmem_U10981 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n14247), .ZN(MEM_stage_inst_dmem_n14242) );
NAND2_X1 MEM_stage_inst_dmem_U10980 ( .A1(MEM_stage_inst_dmem_ram_802), .A2(MEM_stage_inst_dmem_n14246), .ZN(MEM_stage_inst_dmem_n14243) );
NAND2_X1 MEM_stage_inst_dmem_U10979 ( .A1(MEM_stage_inst_dmem_n14241), .A2(MEM_stage_inst_dmem_n14240), .ZN(MEM_stage_inst_dmem_n12126) );
NAND2_X1 MEM_stage_inst_dmem_U10978 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n14247), .ZN(MEM_stage_inst_dmem_n14240) );
NAND2_X1 MEM_stage_inst_dmem_U10977 ( .A1(MEM_stage_inst_dmem_ram_803), .A2(MEM_stage_inst_dmem_n14246), .ZN(MEM_stage_inst_dmem_n14241) );
NAND2_X1 MEM_stage_inst_dmem_U10976 ( .A1(MEM_stage_inst_dmem_n14239), .A2(MEM_stage_inst_dmem_n14238), .ZN(MEM_stage_inst_dmem_n12127) );
NAND2_X1 MEM_stage_inst_dmem_U10975 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n14247), .ZN(MEM_stage_inst_dmem_n14238) );
NAND2_X1 MEM_stage_inst_dmem_U10974 ( .A1(MEM_stage_inst_dmem_ram_804), .A2(MEM_stage_inst_dmem_n14246), .ZN(MEM_stage_inst_dmem_n14239) );
NAND2_X1 MEM_stage_inst_dmem_U10973 ( .A1(MEM_stage_inst_dmem_n14237), .A2(MEM_stage_inst_dmem_n14236), .ZN(MEM_stage_inst_dmem_n12128) );
NAND2_X1 MEM_stage_inst_dmem_U10972 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n14247), .ZN(MEM_stage_inst_dmem_n14236) );
NAND2_X1 MEM_stage_inst_dmem_U10971 ( .A1(MEM_stage_inst_dmem_ram_805), .A2(MEM_stage_inst_dmem_n14246), .ZN(MEM_stage_inst_dmem_n14237) );
NAND2_X1 MEM_stage_inst_dmem_U10970 ( .A1(MEM_stage_inst_dmem_n14235), .A2(MEM_stage_inst_dmem_n14234), .ZN(MEM_stage_inst_dmem_n12129) );
NAND2_X1 MEM_stage_inst_dmem_U10969 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n14247), .ZN(MEM_stage_inst_dmem_n14234) );
NAND2_X1 MEM_stage_inst_dmem_U10968 ( .A1(MEM_stage_inst_dmem_ram_806), .A2(MEM_stage_inst_dmem_n14246), .ZN(MEM_stage_inst_dmem_n14235) );
NAND2_X1 MEM_stage_inst_dmem_U10967 ( .A1(MEM_stage_inst_dmem_n14233), .A2(MEM_stage_inst_dmem_n14232), .ZN(MEM_stage_inst_dmem_n12130) );
NAND2_X1 MEM_stage_inst_dmem_U10966 ( .A1(MEM_stage_inst_dmem_n17), .A2(MEM_stage_inst_dmem_n14247), .ZN(MEM_stage_inst_dmem_n14232) );
NAND2_X1 MEM_stage_inst_dmem_U10965 ( .A1(MEM_stage_inst_dmem_ram_807), .A2(MEM_stage_inst_dmem_n14246), .ZN(MEM_stage_inst_dmem_n14233) );
NAND2_X1 MEM_stage_inst_dmem_U10964 ( .A1(MEM_stage_inst_dmem_n14231), .A2(MEM_stage_inst_dmem_n14230), .ZN(MEM_stage_inst_dmem_n12131) );
NAND2_X1 MEM_stage_inst_dmem_U10963 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n14247), .ZN(MEM_stage_inst_dmem_n14230) );
NAND2_X1 MEM_stage_inst_dmem_U10962 ( .A1(MEM_stage_inst_dmem_ram_808), .A2(MEM_stage_inst_dmem_n14246), .ZN(MEM_stage_inst_dmem_n14231) );
NAND2_X1 MEM_stage_inst_dmem_U10961 ( .A1(MEM_stage_inst_dmem_n14229), .A2(MEM_stage_inst_dmem_n14228), .ZN(MEM_stage_inst_dmem_n12132) );
NAND2_X1 MEM_stage_inst_dmem_U10960 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n14247), .ZN(MEM_stage_inst_dmem_n14228) );
NAND2_X1 MEM_stage_inst_dmem_U10959 ( .A1(MEM_stage_inst_dmem_ram_809), .A2(MEM_stage_inst_dmem_n14246), .ZN(MEM_stage_inst_dmem_n14229) );
NAND2_X1 MEM_stage_inst_dmem_U10958 ( .A1(MEM_stage_inst_dmem_n14227), .A2(MEM_stage_inst_dmem_n14226), .ZN(MEM_stage_inst_dmem_n12133) );
NAND2_X1 MEM_stage_inst_dmem_U10957 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n14247), .ZN(MEM_stage_inst_dmem_n14226) );
NAND2_X1 MEM_stage_inst_dmem_U10956 ( .A1(MEM_stage_inst_dmem_ram_810), .A2(MEM_stage_inst_dmem_n14246), .ZN(MEM_stage_inst_dmem_n14227) );
NAND2_X1 MEM_stage_inst_dmem_U10955 ( .A1(MEM_stage_inst_dmem_n14225), .A2(MEM_stage_inst_dmem_n14224), .ZN(MEM_stage_inst_dmem_n12134) );
NAND2_X1 MEM_stage_inst_dmem_U10954 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n14247), .ZN(MEM_stage_inst_dmem_n14224) );
NAND2_X1 MEM_stage_inst_dmem_U10953 ( .A1(MEM_stage_inst_dmem_ram_811), .A2(MEM_stage_inst_dmem_n14246), .ZN(MEM_stage_inst_dmem_n14225) );
NAND2_X1 MEM_stage_inst_dmem_U10952 ( .A1(MEM_stage_inst_dmem_n14223), .A2(MEM_stage_inst_dmem_n14222), .ZN(MEM_stage_inst_dmem_n12135) );
NAND2_X1 MEM_stage_inst_dmem_U10951 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n14247), .ZN(MEM_stage_inst_dmem_n14222) );
NAND2_X1 MEM_stage_inst_dmem_U10950 ( .A1(MEM_stage_inst_dmem_ram_812), .A2(MEM_stage_inst_dmem_n14246), .ZN(MEM_stage_inst_dmem_n14223) );
NAND2_X1 MEM_stage_inst_dmem_U10949 ( .A1(MEM_stage_inst_dmem_n14221), .A2(MEM_stage_inst_dmem_n14220), .ZN(MEM_stage_inst_dmem_n12136) );
NAND2_X1 MEM_stage_inst_dmem_U10948 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n14247), .ZN(MEM_stage_inst_dmem_n14220) );
NAND2_X1 MEM_stage_inst_dmem_U10947 ( .A1(MEM_stage_inst_dmem_ram_813), .A2(MEM_stage_inst_dmem_n14246), .ZN(MEM_stage_inst_dmem_n14221) );
NAND2_X1 MEM_stage_inst_dmem_U10946 ( .A1(MEM_stage_inst_dmem_n14219), .A2(MEM_stage_inst_dmem_n14218), .ZN(MEM_stage_inst_dmem_n12137) );
NAND2_X1 MEM_stage_inst_dmem_U10945 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n14247), .ZN(MEM_stage_inst_dmem_n14218) );
NAND2_X1 MEM_stage_inst_dmem_U10944 ( .A1(MEM_stage_inst_dmem_ram_814), .A2(MEM_stage_inst_dmem_n14246), .ZN(MEM_stage_inst_dmem_n14219) );
NAND2_X1 MEM_stage_inst_dmem_U10943 ( .A1(MEM_stage_inst_dmem_n14217), .A2(MEM_stage_inst_dmem_n14216), .ZN(MEM_stage_inst_dmem_n12138) );
NAND2_X1 MEM_stage_inst_dmem_U10942 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n14247), .ZN(MEM_stage_inst_dmem_n14216) );
INV_X1 MEM_stage_inst_dmem_U10941 ( .A(MEM_stage_inst_dmem_n14246), .ZN(MEM_stage_inst_dmem_n14247) );
NAND2_X1 MEM_stage_inst_dmem_U10940 ( .A1(MEM_stage_inst_dmem_ram_815), .A2(MEM_stage_inst_dmem_n14246), .ZN(MEM_stage_inst_dmem_n14217) );
NAND2_X1 MEM_stage_inst_dmem_U10939 ( .A1(MEM_stage_inst_dmem_n21394), .A2(MEM_stage_inst_dmem_n14284), .ZN(MEM_stage_inst_dmem_n14246) );
NAND2_X1 MEM_stage_inst_dmem_U10938 ( .A1(MEM_stage_inst_dmem_n14215), .A2(MEM_stage_inst_dmem_n14214), .ZN(MEM_stage_inst_dmem_n12139) );
NAND2_X1 MEM_stage_inst_dmem_U10937 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n14213), .ZN(MEM_stage_inst_dmem_n14214) );
NAND2_X1 MEM_stage_inst_dmem_U10936 ( .A1(MEM_stage_inst_dmem_ram_816), .A2(MEM_stage_inst_dmem_n14212), .ZN(MEM_stage_inst_dmem_n14215) );
NAND2_X1 MEM_stage_inst_dmem_U10935 ( .A1(MEM_stage_inst_dmem_n14211), .A2(MEM_stage_inst_dmem_n14210), .ZN(MEM_stage_inst_dmem_n12140) );
NAND2_X1 MEM_stage_inst_dmem_U10934 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n14213), .ZN(MEM_stage_inst_dmem_n14210) );
NAND2_X1 MEM_stage_inst_dmem_U10933 ( .A1(MEM_stage_inst_dmem_ram_817), .A2(MEM_stage_inst_dmem_n14212), .ZN(MEM_stage_inst_dmem_n14211) );
NAND2_X1 MEM_stage_inst_dmem_U10932 ( .A1(MEM_stage_inst_dmem_n14209), .A2(MEM_stage_inst_dmem_n14208), .ZN(MEM_stage_inst_dmem_n12141) );
NAND2_X1 MEM_stage_inst_dmem_U10931 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n14213), .ZN(MEM_stage_inst_dmem_n14208) );
NAND2_X1 MEM_stage_inst_dmem_U10930 ( .A1(MEM_stage_inst_dmem_ram_818), .A2(MEM_stage_inst_dmem_n14212), .ZN(MEM_stage_inst_dmem_n14209) );
NAND2_X1 MEM_stage_inst_dmem_U10929 ( .A1(MEM_stage_inst_dmem_n14207), .A2(MEM_stage_inst_dmem_n14206), .ZN(MEM_stage_inst_dmem_n12142) );
NAND2_X1 MEM_stage_inst_dmem_U10928 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n14213), .ZN(MEM_stage_inst_dmem_n14206) );
NAND2_X1 MEM_stage_inst_dmem_U10927 ( .A1(MEM_stage_inst_dmem_ram_819), .A2(MEM_stage_inst_dmem_n14212), .ZN(MEM_stage_inst_dmem_n14207) );
NAND2_X1 MEM_stage_inst_dmem_U10926 ( .A1(MEM_stage_inst_dmem_n14205), .A2(MEM_stage_inst_dmem_n14204), .ZN(MEM_stage_inst_dmem_n12143) );
NAND2_X1 MEM_stage_inst_dmem_U10925 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n14213), .ZN(MEM_stage_inst_dmem_n14204) );
NAND2_X1 MEM_stage_inst_dmem_U10924 ( .A1(MEM_stage_inst_dmem_ram_820), .A2(MEM_stage_inst_dmem_n14212), .ZN(MEM_stage_inst_dmem_n14205) );
NAND2_X1 MEM_stage_inst_dmem_U10923 ( .A1(MEM_stage_inst_dmem_n14203), .A2(MEM_stage_inst_dmem_n14202), .ZN(MEM_stage_inst_dmem_n12144) );
NAND2_X1 MEM_stage_inst_dmem_U10922 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n14213), .ZN(MEM_stage_inst_dmem_n14202) );
NAND2_X1 MEM_stage_inst_dmem_U10921 ( .A1(MEM_stage_inst_dmem_ram_821), .A2(MEM_stage_inst_dmem_n14212), .ZN(MEM_stage_inst_dmem_n14203) );
NAND2_X1 MEM_stage_inst_dmem_U10920 ( .A1(MEM_stage_inst_dmem_n14201), .A2(MEM_stage_inst_dmem_n14200), .ZN(MEM_stage_inst_dmem_n12145) );
NAND2_X1 MEM_stage_inst_dmem_U10919 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n14213), .ZN(MEM_stage_inst_dmem_n14200) );
NAND2_X1 MEM_stage_inst_dmem_U10918 ( .A1(MEM_stage_inst_dmem_ram_822), .A2(MEM_stage_inst_dmem_n14212), .ZN(MEM_stage_inst_dmem_n14201) );
NAND2_X1 MEM_stage_inst_dmem_U10917 ( .A1(MEM_stage_inst_dmem_n14199), .A2(MEM_stage_inst_dmem_n14198), .ZN(MEM_stage_inst_dmem_n12146) );
NAND2_X1 MEM_stage_inst_dmem_U10916 ( .A1(MEM_stage_inst_dmem_n18), .A2(MEM_stage_inst_dmem_n14213), .ZN(MEM_stage_inst_dmem_n14198) );
NAND2_X1 MEM_stage_inst_dmem_U10915 ( .A1(MEM_stage_inst_dmem_ram_823), .A2(MEM_stage_inst_dmem_n14212), .ZN(MEM_stage_inst_dmem_n14199) );
NAND2_X1 MEM_stage_inst_dmem_U10914 ( .A1(MEM_stage_inst_dmem_n14197), .A2(MEM_stage_inst_dmem_n14196), .ZN(MEM_stage_inst_dmem_n12147) );
NAND2_X1 MEM_stage_inst_dmem_U10913 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n14213), .ZN(MEM_stage_inst_dmem_n14196) );
NAND2_X1 MEM_stage_inst_dmem_U10912 ( .A1(MEM_stage_inst_dmem_ram_824), .A2(MEM_stage_inst_dmem_n14212), .ZN(MEM_stage_inst_dmem_n14197) );
NAND2_X1 MEM_stage_inst_dmem_U10911 ( .A1(MEM_stage_inst_dmem_n14195), .A2(MEM_stage_inst_dmem_n14194), .ZN(MEM_stage_inst_dmem_n12148) );
NAND2_X1 MEM_stage_inst_dmem_U10910 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n14213), .ZN(MEM_stage_inst_dmem_n14194) );
NAND2_X1 MEM_stage_inst_dmem_U10909 ( .A1(MEM_stage_inst_dmem_ram_825), .A2(MEM_stage_inst_dmem_n14212), .ZN(MEM_stage_inst_dmem_n14195) );
NAND2_X1 MEM_stage_inst_dmem_U10908 ( .A1(MEM_stage_inst_dmem_n14193), .A2(MEM_stage_inst_dmem_n14192), .ZN(MEM_stage_inst_dmem_n12149) );
NAND2_X1 MEM_stage_inst_dmem_U10907 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n14213), .ZN(MEM_stage_inst_dmem_n14192) );
NAND2_X1 MEM_stage_inst_dmem_U10906 ( .A1(MEM_stage_inst_dmem_ram_826), .A2(MEM_stage_inst_dmem_n14212), .ZN(MEM_stage_inst_dmem_n14193) );
NAND2_X1 MEM_stage_inst_dmem_U10905 ( .A1(MEM_stage_inst_dmem_n14191), .A2(MEM_stage_inst_dmem_n14190), .ZN(MEM_stage_inst_dmem_n12150) );
NAND2_X1 MEM_stage_inst_dmem_U10904 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n14213), .ZN(MEM_stage_inst_dmem_n14190) );
NAND2_X1 MEM_stage_inst_dmem_U10903 ( .A1(MEM_stage_inst_dmem_ram_827), .A2(MEM_stage_inst_dmem_n14212), .ZN(MEM_stage_inst_dmem_n14191) );
NAND2_X1 MEM_stage_inst_dmem_U10902 ( .A1(MEM_stage_inst_dmem_n14189), .A2(MEM_stage_inst_dmem_n14188), .ZN(MEM_stage_inst_dmem_n12151) );
NAND2_X1 MEM_stage_inst_dmem_U10901 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n14213), .ZN(MEM_stage_inst_dmem_n14188) );
NAND2_X1 MEM_stage_inst_dmem_U10900 ( .A1(MEM_stage_inst_dmem_ram_828), .A2(MEM_stage_inst_dmem_n14212), .ZN(MEM_stage_inst_dmem_n14189) );
NAND2_X1 MEM_stage_inst_dmem_U10899 ( .A1(MEM_stage_inst_dmem_n14187), .A2(MEM_stage_inst_dmem_n14186), .ZN(MEM_stage_inst_dmem_n12152) );
NAND2_X1 MEM_stage_inst_dmem_U10898 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n14213), .ZN(MEM_stage_inst_dmem_n14186) );
NAND2_X1 MEM_stage_inst_dmem_U10897 ( .A1(MEM_stage_inst_dmem_ram_829), .A2(MEM_stage_inst_dmem_n14212), .ZN(MEM_stage_inst_dmem_n14187) );
NAND2_X1 MEM_stage_inst_dmem_U10896 ( .A1(MEM_stage_inst_dmem_n14185), .A2(MEM_stage_inst_dmem_n14184), .ZN(MEM_stage_inst_dmem_n12153) );
NAND2_X1 MEM_stage_inst_dmem_U10895 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n14213), .ZN(MEM_stage_inst_dmem_n14184) );
NAND2_X1 MEM_stage_inst_dmem_U10894 ( .A1(MEM_stage_inst_dmem_ram_830), .A2(MEM_stage_inst_dmem_n14212), .ZN(MEM_stage_inst_dmem_n14185) );
NAND2_X1 MEM_stage_inst_dmem_U10893 ( .A1(MEM_stage_inst_dmem_n14183), .A2(MEM_stage_inst_dmem_n14182), .ZN(MEM_stage_inst_dmem_n12154) );
NAND2_X1 MEM_stage_inst_dmem_U10892 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n14213), .ZN(MEM_stage_inst_dmem_n14182) );
NAND2_X1 MEM_stage_inst_dmem_U10891 ( .A1(MEM_stage_inst_dmem_ram_831), .A2(MEM_stage_inst_dmem_n14212), .ZN(MEM_stage_inst_dmem_n14183) );
NAND2_X1 MEM_stage_inst_dmem_U10890 ( .A1(MEM_stage_inst_dmem_n21359), .A2(MEM_stage_inst_dmem_n14284), .ZN(MEM_stage_inst_dmem_n14212) );
NAND2_X1 MEM_stage_inst_dmem_U10889 ( .A1(MEM_stage_inst_dmem_n14181), .A2(MEM_stage_inst_dmem_n14180), .ZN(MEM_stage_inst_dmem_n12155) );
NAND2_X1 MEM_stage_inst_dmem_U10888 ( .A1(MEM_stage_inst_dmem_n15145), .A2(MEM_stage_inst_dmem_n14179), .ZN(MEM_stage_inst_dmem_n14180) );
NAND2_X1 MEM_stage_inst_dmem_U10887 ( .A1(MEM_stage_inst_dmem_ram_832), .A2(MEM_stage_inst_dmem_n14178), .ZN(MEM_stage_inst_dmem_n14181) );
NAND2_X1 MEM_stage_inst_dmem_U10886 ( .A1(MEM_stage_inst_dmem_n14177), .A2(MEM_stage_inst_dmem_n14176), .ZN(MEM_stage_inst_dmem_n12156) );
NAND2_X1 MEM_stage_inst_dmem_U10885 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n14179), .ZN(MEM_stage_inst_dmem_n14176) );
NAND2_X1 MEM_stage_inst_dmem_U10884 ( .A1(MEM_stage_inst_dmem_ram_833), .A2(MEM_stage_inst_dmem_n14178), .ZN(MEM_stage_inst_dmem_n14177) );
NAND2_X1 MEM_stage_inst_dmem_U10883 ( .A1(MEM_stage_inst_dmem_n14175), .A2(MEM_stage_inst_dmem_n14174), .ZN(MEM_stage_inst_dmem_n12157) );
NAND2_X1 MEM_stage_inst_dmem_U10882 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n14179), .ZN(MEM_stage_inst_dmem_n14174) );
NAND2_X1 MEM_stage_inst_dmem_U10881 ( .A1(MEM_stage_inst_dmem_ram_834), .A2(MEM_stage_inst_dmem_n14178), .ZN(MEM_stage_inst_dmem_n14175) );
NAND2_X1 MEM_stage_inst_dmem_U10880 ( .A1(MEM_stage_inst_dmem_n14173), .A2(MEM_stage_inst_dmem_n14172), .ZN(MEM_stage_inst_dmem_n12158) );
NAND2_X1 MEM_stage_inst_dmem_U10879 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n14179), .ZN(MEM_stage_inst_dmem_n14172) );
NAND2_X1 MEM_stage_inst_dmem_U10878 ( .A1(MEM_stage_inst_dmem_ram_835), .A2(MEM_stage_inst_dmem_n14178), .ZN(MEM_stage_inst_dmem_n14173) );
NAND2_X1 MEM_stage_inst_dmem_U10877 ( .A1(MEM_stage_inst_dmem_n14171), .A2(MEM_stage_inst_dmem_n14170), .ZN(MEM_stage_inst_dmem_n12159) );
NAND2_X1 MEM_stage_inst_dmem_U10876 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n14179), .ZN(MEM_stage_inst_dmem_n14170) );
NAND2_X1 MEM_stage_inst_dmem_U10875 ( .A1(MEM_stage_inst_dmem_ram_836), .A2(MEM_stage_inst_dmem_n14178), .ZN(MEM_stage_inst_dmem_n14171) );
NAND2_X1 MEM_stage_inst_dmem_U10874 ( .A1(MEM_stage_inst_dmem_n14169), .A2(MEM_stage_inst_dmem_n14168), .ZN(MEM_stage_inst_dmem_n12160) );
NAND2_X1 MEM_stage_inst_dmem_U10873 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n14179), .ZN(MEM_stage_inst_dmem_n14168) );
NAND2_X1 MEM_stage_inst_dmem_U10872 ( .A1(MEM_stage_inst_dmem_ram_837), .A2(MEM_stage_inst_dmem_n14178), .ZN(MEM_stage_inst_dmem_n14169) );
NAND2_X1 MEM_stage_inst_dmem_U10871 ( .A1(MEM_stage_inst_dmem_n14167), .A2(MEM_stage_inst_dmem_n14166), .ZN(MEM_stage_inst_dmem_n12161) );
NAND2_X1 MEM_stage_inst_dmem_U10870 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n14179), .ZN(MEM_stage_inst_dmem_n14166) );
NAND2_X1 MEM_stage_inst_dmem_U10869 ( .A1(MEM_stage_inst_dmem_ram_838), .A2(MEM_stage_inst_dmem_n14178), .ZN(MEM_stage_inst_dmem_n14167) );
NAND2_X1 MEM_stage_inst_dmem_U10868 ( .A1(MEM_stage_inst_dmem_n14165), .A2(MEM_stage_inst_dmem_n14164), .ZN(MEM_stage_inst_dmem_n12162) );
NAND2_X1 MEM_stage_inst_dmem_U10867 ( .A1(MEM_stage_inst_dmem_n17), .A2(MEM_stage_inst_dmem_n14179), .ZN(MEM_stage_inst_dmem_n14164) );
NAND2_X1 MEM_stage_inst_dmem_U10866 ( .A1(MEM_stage_inst_dmem_ram_839), .A2(MEM_stage_inst_dmem_n14178), .ZN(MEM_stage_inst_dmem_n14165) );
NAND2_X1 MEM_stage_inst_dmem_U10865 ( .A1(MEM_stage_inst_dmem_n14163), .A2(MEM_stage_inst_dmem_n14162), .ZN(MEM_stage_inst_dmem_n12163) );
NAND2_X1 MEM_stage_inst_dmem_U10864 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n14179), .ZN(MEM_stage_inst_dmem_n14162) );
NAND2_X1 MEM_stage_inst_dmem_U10863 ( .A1(MEM_stage_inst_dmem_ram_840), .A2(MEM_stage_inst_dmem_n14178), .ZN(MEM_stage_inst_dmem_n14163) );
NAND2_X1 MEM_stage_inst_dmem_U10862 ( .A1(MEM_stage_inst_dmem_n14161), .A2(MEM_stage_inst_dmem_n14160), .ZN(MEM_stage_inst_dmem_n12164) );
NAND2_X1 MEM_stage_inst_dmem_U10861 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n14179), .ZN(MEM_stage_inst_dmem_n14160) );
NAND2_X1 MEM_stage_inst_dmem_U10860 ( .A1(MEM_stage_inst_dmem_ram_841), .A2(MEM_stage_inst_dmem_n14178), .ZN(MEM_stage_inst_dmem_n14161) );
NAND2_X1 MEM_stage_inst_dmem_U10859 ( .A1(MEM_stage_inst_dmem_n14159), .A2(MEM_stage_inst_dmem_n14158), .ZN(MEM_stage_inst_dmem_n12165) );
NAND2_X1 MEM_stage_inst_dmem_U10858 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n14179), .ZN(MEM_stage_inst_dmem_n14158) );
NAND2_X1 MEM_stage_inst_dmem_U10857 ( .A1(MEM_stage_inst_dmem_ram_842), .A2(MEM_stage_inst_dmem_n14178), .ZN(MEM_stage_inst_dmem_n14159) );
NAND2_X1 MEM_stage_inst_dmem_U10856 ( .A1(MEM_stage_inst_dmem_n14157), .A2(MEM_stage_inst_dmem_n14156), .ZN(MEM_stage_inst_dmem_n12166) );
NAND2_X1 MEM_stage_inst_dmem_U10855 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n14179), .ZN(MEM_stage_inst_dmem_n14156) );
NAND2_X1 MEM_stage_inst_dmem_U10854 ( .A1(MEM_stage_inst_dmem_ram_843), .A2(MEM_stage_inst_dmem_n14178), .ZN(MEM_stage_inst_dmem_n14157) );
NAND2_X1 MEM_stage_inst_dmem_U10853 ( .A1(MEM_stage_inst_dmem_n14155), .A2(MEM_stage_inst_dmem_n14154), .ZN(MEM_stage_inst_dmem_n12167) );
NAND2_X1 MEM_stage_inst_dmem_U10852 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n14179), .ZN(MEM_stage_inst_dmem_n14154) );
NAND2_X1 MEM_stage_inst_dmem_U10851 ( .A1(MEM_stage_inst_dmem_ram_844), .A2(MEM_stage_inst_dmem_n14178), .ZN(MEM_stage_inst_dmem_n14155) );
NAND2_X1 MEM_stage_inst_dmem_U10850 ( .A1(MEM_stage_inst_dmem_n14153), .A2(MEM_stage_inst_dmem_n14152), .ZN(MEM_stage_inst_dmem_n12168) );
NAND2_X1 MEM_stage_inst_dmem_U10849 ( .A1(MEM_stage_inst_dmem_n15116), .A2(MEM_stage_inst_dmem_n14179), .ZN(MEM_stage_inst_dmem_n14152) );
NAND2_X1 MEM_stage_inst_dmem_U10848 ( .A1(MEM_stage_inst_dmem_ram_845), .A2(MEM_stage_inst_dmem_n14178), .ZN(MEM_stage_inst_dmem_n14153) );
NAND2_X1 MEM_stage_inst_dmem_U10847 ( .A1(MEM_stage_inst_dmem_n14151), .A2(MEM_stage_inst_dmem_n14150), .ZN(MEM_stage_inst_dmem_n12169) );
NAND2_X1 MEM_stage_inst_dmem_U10846 ( .A1(MEM_stage_inst_dmem_n15113), .A2(MEM_stage_inst_dmem_n14179), .ZN(MEM_stage_inst_dmem_n14150) );
NAND2_X1 MEM_stage_inst_dmem_U10845 ( .A1(MEM_stage_inst_dmem_ram_846), .A2(MEM_stage_inst_dmem_n14178), .ZN(MEM_stage_inst_dmem_n14151) );
NAND2_X1 MEM_stage_inst_dmem_U10844 ( .A1(MEM_stage_inst_dmem_n14149), .A2(MEM_stage_inst_dmem_n14148), .ZN(MEM_stage_inst_dmem_n12170) );
NAND2_X1 MEM_stage_inst_dmem_U10843 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n14179), .ZN(MEM_stage_inst_dmem_n14148) );
INV_X1 MEM_stage_inst_dmem_U10842 ( .A(MEM_stage_inst_dmem_n14178), .ZN(MEM_stage_inst_dmem_n14179) );
NAND2_X1 MEM_stage_inst_dmem_U10841 ( .A1(MEM_stage_inst_dmem_ram_847), .A2(MEM_stage_inst_dmem_n14178), .ZN(MEM_stage_inst_dmem_n14149) );
NAND2_X1 MEM_stage_inst_dmem_U10840 ( .A1(MEM_stage_inst_dmem_n21319), .A2(MEM_stage_inst_dmem_n14284), .ZN(MEM_stage_inst_dmem_n14178) );
NAND2_X1 MEM_stage_inst_dmem_U10839 ( .A1(MEM_stage_inst_dmem_n14147), .A2(MEM_stage_inst_dmem_n14146), .ZN(MEM_stage_inst_dmem_n12171) );
NAND2_X1 MEM_stage_inst_dmem_U10838 ( .A1(MEM_stage_inst_dmem_n14732), .A2(MEM_stage_inst_dmem_n14145), .ZN(MEM_stage_inst_dmem_n14146) );
NAND2_X1 MEM_stage_inst_dmem_U10837 ( .A1(MEM_stage_inst_dmem_ram_848), .A2(MEM_stage_inst_dmem_n14144), .ZN(MEM_stage_inst_dmem_n14147) );
NAND2_X1 MEM_stage_inst_dmem_U10836 ( .A1(MEM_stage_inst_dmem_n14143), .A2(MEM_stage_inst_dmem_n14142), .ZN(MEM_stage_inst_dmem_n12172) );
NAND2_X1 MEM_stage_inst_dmem_U10835 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n14145), .ZN(MEM_stage_inst_dmem_n14142) );
NAND2_X1 MEM_stage_inst_dmem_U10834 ( .A1(MEM_stage_inst_dmem_ram_849), .A2(MEM_stage_inst_dmem_n14144), .ZN(MEM_stage_inst_dmem_n14143) );
NAND2_X1 MEM_stage_inst_dmem_U10833 ( .A1(MEM_stage_inst_dmem_n14141), .A2(MEM_stage_inst_dmem_n14140), .ZN(MEM_stage_inst_dmem_n12173) );
NAND2_X1 MEM_stage_inst_dmem_U10832 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n14145), .ZN(MEM_stage_inst_dmem_n14140) );
NAND2_X1 MEM_stage_inst_dmem_U10831 ( .A1(MEM_stage_inst_dmem_ram_850), .A2(MEM_stage_inst_dmem_n14144), .ZN(MEM_stage_inst_dmem_n14141) );
NAND2_X1 MEM_stage_inst_dmem_U10830 ( .A1(MEM_stage_inst_dmem_n14139), .A2(MEM_stage_inst_dmem_n14138), .ZN(MEM_stage_inst_dmem_n12174) );
NAND2_X1 MEM_stage_inst_dmem_U10829 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n14145), .ZN(MEM_stage_inst_dmem_n14138) );
NAND2_X1 MEM_stage_inst_dmem_U10828 ( .A1(MEM_stage_inst_dmem_ram_851), .A2(MEM_stage_inst_dmem_n14144), .ZN(MEM_stage_inst_dmem_n14139) );
NAND2_X1 MEM_stage_inst_dmem_U10827 ( .A1(MEM_stage_inst_dmem_n14137), .A2(MEM_stage_inst_dmem_n14136), .ZN(MEM_stage_inst_dmem_n12175) );
NAND2_X1 MEM_stage_inst_dmem_U10826 ( .A1(MEM_stage_inst_dmem_n16784), .A2(MEM_stage_inst_dmem_n14145), .ZN(MEM_stage_inst_dmem_n14136) );
NAND2_X1 MEM_stage_inst_dmem_U10825 ( .A1(MEM_stage_inst_dmem_ram_852), .A2(MEM_stage_inst_dmem_n14144), .ZN(MEM_stage_inst_dmem_n14137) );
NAND2_X1 MEM_stage_inst_dmem_U10824 ( .A1(MEM_stage_inst_dmem_n14135), .A2(MEM_stage_inst_dmem_n14134), .ZN(MEM_stage_inst_dmem_n12176) );
NAND2_X1 MEM_stage_inst_dmem_U10823 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n14145), .ZN(MEM_stage_inst_dmem_n14134) );
NAND2_X1 MEM_stage_inst_dmem_U10822 ( .A1(MEM_stage_inst_dmem_ram_853), .A2(MEM_stage_inst_dmem_n14144), .ZN(MEM_stage_inst_dmem_n14135) );
NAND2_X1 MEM_stage_inst_dmem_U10821 ( .A1(MEM_stage_inst_dmem_n14133), .A2(MEM_stage_inst_dmem_n14132), .ZN(MEM_stage_inst_dmem_n12177) );
NAND2_X1 MEM_stage_inst_dmem_U10820 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n14145), .ZN(MEM_stage_inst_dmem_n14132) );
NAND2_X1 MEM_stage_inst_dmem_U10819 ( .A1(MEM_stage_inst_dmem_ram_854), .A2(MEM_stage_inst_dmem_n14144), .ZN(MEM_stage_inst_dmem_n14133) );
NAND2_X1 MEM_stage_inst_dmem_U10818 ( .A1(MEM_stage_inst_dmem_n14131), .A2(MEM_stage_inst_dmem_n14130), .ZN(MEM_stage_inst_dmem_n12178) );
NAND2_X1 MEM_stage_inst_dmem_U10817 ( .A1(MEM_stage_inst_dmem_n18), .A2(MEM_stage_inst_dmem_n14145), .ZN(MEM_stage_inst_dmem_n14130) );
NAND2_X1 MEM_stage_inst_dmem_U10816 ( .A1(MEM_stage_inst_dmem_ram_855), .A2(MEM_stage_inst_dmem_n14144), .ZN(MEM_stage_inst_dmem_n14131) );
NAND2_X1 MEM_stage_inst_dmem_U10815 ( .A1(MEM_stage_inst_dmem_n14129), .A2(MEM_stage_inst_dmem_n14128), .ZN(MEM_stage_inst_dmem_n12179) );
NAND2_X1 MEM_stage_inst_dmem_U10814 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n14145), .ZN(MEM_stage_inst_dmem_n14128) );
NAND2_X1 MEM_stage_inst_dmem_U10813 ( .A1(MEM_stage_inst_dmem_ram_856), .A2(MEM_stage_inst_dmem_n14144), .ZN(MEM_stage_inst_dmem_n14129) );
NAND2_X1 MEM_stage_inst_dmem_U10812 ( .A1(MEM_stage_inst_dmem_n14127), .A2(MEM_stage_inst_dmem_n14126), .ZN(MEM_stage_inst_dmem_n12180) );
NAND2_X1 MEM_stage_inst_dmem_U10811 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n14145), .ZN(MEM_stage_inst_dmem_n14126) );
NAND2_X1 MEM_stage_inst_dmem_U10810 ( .A1(MEM_stage_inst_dmem_ram_857), .A2(MEM_stage_inst_dmem_n14144), .ZN(MEM_stage_inst_dmem_n14127) );
NAND2_X1 MEM_stage_inst_dmem_U10809 ( .A1(MEM_stage_inst_dmem_n14125), .A2(MEM_stage_inst_dmem_n14124), .ZN(MEM_stage_inst_dmem_n12181) );
NAND2_X1 MEM_stage_inst_dmem_U10808 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n14145), .ZN(MEM_stage_inst_dmem_n14124) );
NAND2_X1 MEM_stage_inst_dmem_U10807 ( .A1(MEM_stage_inst_dmem_ram_858), .A2(MEM_stage_inst_dmem_n14144), .ZN(MEM_stage_inst_dmem_n14125) );
NAND2_X1 MEM_stage_inst_dmem_U10806 ( .A1(MEM_stage_inst_dmem_n14123), .A2(MEM_stage_inst_dmem_n14122), .ZN(MEM_stage_inst_dmem_n12182) );
NAND2_X1 MEM_stage_inst_dmem_U10805 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n14145), .ZN(MEM_stage_inst_dmem_n14122) );
NAND2_X1 MEM_stage_inst_dmem_U10804 ( .A1(MEM_stage_inst_dmem_ram_859), .A2(MEM_stage_inst_dmem_n14144), .ZN(MEM_stage_inst_dmem_n14123) );
NAND2_X1 MEM_stage_inst_dmem_U10803 ( .A1(MEM_stage_inst_dmem_n14121), .A2(MEM_stage_inst_dmem_n14120), .ZN(MEM_stage_inst_dmem_n12183) );
NAND2_X1 MEM_stage_inst_dmem_U10802 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n14145), .ZN(MEM_stage_inst_dmem_n14120) );
NAND2_X1 MEM_stage_inst_dmem_U10801 ( .A1(MEM_stage_inst_dmem_ram_860), .A2(MEM_stage_inst_dmem_n14144), .ZN(MEM_stage_inst_dmem_n14121) );
NAND2_X1 MEM_stage_inst_dmem_U10800 ( .A1(MEM_stage_inst_dmem_n14119), .A2(MEM_stage_inst_dmem_n14118), .ZN(MEM_stage_inst_dmem_n12184) );
NAND2_X1 MEM_stage_inst_dmem_U10799 ( .A1(MEM_stage_inst_dmem_n116), .A2(MEM_stage_inst_dmem_n14145), .ZN(MEM_stage_inst_dmem_n14118) );
NAND2_X1 MEM_stage_inst_dmem_U10798 ( .A1(MEM_stage_inst_dmem_ram_861), .A2(MEM_stage_inst_dmem_n14144), .ZN(MEM_stage_inst_dmem_n14119) );
NAND2_X1 MEM_stage_inst_dmem_U10797 ( .A1(MEM_stage_inst_dmem_n14117), .A2(MEM_stage_inst_dmem_n14116), .ZN(MEM_stage_inst_dmem_n12185) );
NAND2_X1 MEM_stage_inst_dmem_U10796 ( .A1(MEM_stage_inst_dmem_n14696), .A2(MEM_stage_inst_dmem_n14145), .ZN(MEM_stage_inst_dmem_n14116) );
NAND2_X1 MEM_stage_inst_dmem_U10795 ( .A1(MEM_stage_inst_dmem_ram_862), .A2(MEM_stage_inst_dmem_n14144), .ZN(MEM_stage_inst_dmem_n14117) );
NAND2_X1 MEM_stage_inst_dmem_U10794 ( .A1(MEM_stage_inst_dmem_n14115), .A2(MEM_stage_inst_dmem_n14114), .ZN(MEM_stage_inst_dmem_n12186) );
NAND2_X1 MEM_stage_inst_dmem_U10793 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n14145), .ZN(MEM_stage_inst_dmem_n14114) );
INV_X1 MEM_stage_inst_dmem_U10792 ( .A(MEM_stage_inst_dmem_n14144), .ZN(MEM_stage_inst_dmem_n14145) );
NAND2_X1 MEM_stage_inst_dmem_U10791 ( .A1(MEM_stage_inst_dmem_ram_863), .A2(MEM_stage_inst_dmem_n14144), .ZN(MEM_stage_inst_dmem_n14115) );
NAND2_X1 MEM_stage_inst_dmem_U10790 ( .A1(MEM_stage_inst_dmem_n21284), .A2(MEM_stage_inst_dmem_n14284), .ZN(MEM_stage_inst_dmem_n14144) );
NAND2_X1 MEM_stage_inst_dmem_U10789 ( .A1(MEM_stage_inst_dmem_n14113), .A2(MEM_stage_inst_dmem_n14112), .ZN(MEM_stage_inst_dmem_n12187) );
NAND2_X1 MEM_stage_inst_dmem_U10788 ( .A1(MEM_stage_inst_dmem_n19275), .A2(MEM_stage_inst_dmem_n14111), .ZN(MEM_stage_inst_dmem_n14112) );
NAND2_X1 MEM_stage_inst_dmem_U10787 ( .A1(MEM_stage_inst_dmem_ram_864), .A2(MEM_stage_inst_dmem_n14110), .ZN(MEM_stage_inst_dmem_n14113) );
NAND2_X1 MEM_stage_inst_dmem_U10786 ( .A1(MEM_stage_inst_dmem_n14109), .A2(MEM_stage_inst_dmem_n14108), .ZN(MEM_stage_inst_dmem_n12188) );
NAND2_X1 MEM_stage_inst_dmem_U10785 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n14111), .ZN(MEM_stage_inst_dmem_n14108) );
NAND2_X1 MEM_stage_inst_dmem_U10784 ( .A1(MEM_stage_inst_dmem_ram_865), .A2(MEM_stage_inst_dmem_n14110), .ZN(MEM_stage_inst_dmem_n14109) );
NAND2_X1 MEM_stage_inst_dmem_U10783 ( .A1(MEM_stage_inst_dmem_n14107), .A2(MEM_stage_inst_dmem_n14106), .ZN(MEM_stage_inst_dmem_n12189) );
NAND2_X1 MEM_stage_inst_dmem_U10782 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n14111), .ZN(MEM_stage_inst_dmem_n14106) );
NAND2_X1 MEM_stage_inst_dmem_U10781 ( .A1(MEM_stage_inst_dmem_ram_866), .A2(MEM_stage_inst_dmem_n14110), .ZN(MEM_stage_inst_dmem_n14107) );
NAND2_X1 MEM_stage_inst_dmem_U10780 ( .A1(MEM_stage_inst_dmem_n14105), .A2(MEM_stage_inst_dmem_n14104), .ZN(MEM_stage_inst_dmem_n12190) );
NAND2_X1 MEM_stage_inst_dmem_U10779 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n14111), .ZN(MEM_stage_inst_dmem_n14104) );
NAND2_X1 MEM_stage_inst_dmem_U10778 ( .A1(MEM_stage_inst_dmem_ram_867), .A2(MEM_stage_inst_dmem_n14110), .ZN(MEM_stage_inst_dmem_n14105) );
NAND2_X1 MEM_stage_inst_dmem_U10777 ( .A1(MEM_stage_inst_dmem_n14103), .A2(MEM_stage_inst_dmem_n14102), .ZN(MEM_stage_inst_dmem_n12191) );
NAND2_X1 MEM_stage_inst_dmem_U10776 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n14111), .ZN(MEM_stage_inst_dmem_n14102) );
NAND2_X1 MEM_stage_inst_dmem_U10775 ( .A1(MEM_stage_inst_dmem_ram_868), .A2(MEM_stage_inst_dmem_n14110), .ZN(MEM_stage_inst_dmem_n14103) );
NAND2_X1 MEM_stage_inst_dmem_U10774 ( .A1(MEM_stage_inst_dmem_n14101), .A2(MEM_stage_inst_dmem_n14100), .ZN(MEM_stage_inst_dmem_n12192) );
NAND2_X1 MEM_stage_inst_dmem_U10773 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n14111), .ZN(MEM_stage_inst_dmem_n14100) );
NAND2_X1 MEM_stage_inst_dmem_U10772 ( .A1(MEM_stage_inst_dmem_ram_869), .A2(MEM_stage_inst_dmem_n14110), .ZN(MEM_stage_inst_dmem_n14101) );
NAND2_X1 MEM_stage_inst_dmem_U10771 ( .A1(MEM_stage_inst_dmem_n14099), .A2(MEM_stage_inst_dmem_n14098), .ZN(MEM_stage_inst_dmem_n12193) );
NAND2_X1 MEM_stage_inst_dmem_U10770 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n14111), .ZN(MEM_stage_inst_dmem_n14098) );
NAND2_X1 MEM_stage_inst_dmem_U10769 ( .A1(MEM_stage_inst_dmem_ram_870), .A2(MEM_stage_inst_dmem_n14110), .ZN(MEM_stage_inst_dmem_n14099) );
NAND2_X1 MEM_stage_inst_dmem_U10768 ( .A1(MEM_stage_inst_dmem_n14097), .A2(MEM_stage_inst_dmem_n14096), .ZN(MEM_stage_inst_dmem_n12194) );
NAND2_X1 MEM_stage_inst_dmem_U10767 ( .A1(MEM_stage_inst_dmem_n17), .A2(MEM_stage_inst_dmem_n14111), .ZN(MEM_stage_inst_dmem_n14096) );
NAND2_X1 MEM_stage_inst_dmem_U10766 ( .A1(MEM_stage_inst_dmem_ram_871), .A2(MEM_stage_inst_dmem_n14110), .ZN(MEM_stage_inst_dmem_n14097) );
NAND2_X1 MEM_stage_inst_dmem_U10765 ( .A1(MEM_stage_inst_dmem_n14095), .A2(MEM_stage_inst_dmem_n14094), .ZN(MEM_stage_inst_dmem_n12195) );
NAND2_X1 MEM_stage_inst_dmem_U10764 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n14111), .ZN(MEM_stage_inst_dmem_n14094) );
NAND2_X1 MEM_stage_inst_dmem_U10763 ( .A1(MEM_stage_inst_dmem_ram_872), .A2(MEM_stage_inst_dmem_n14110), .ZN(MEM_stage_inst_dmem_n14095) );
NAND2_X1 MEM_stage_inst_dmem_U10762 ( .A1(MEM_stage_inst_dmem_n14093), .A2(MEM_stage_inst_dmem_n14092), .ZN(MEM_stage_inst_dmem_n12196) );
NAND2_X1 MEM_stage_inst_dmem_U10761 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n14111), .ZN(MEM_stage_inst_dmem_n14092) );
NAND2_X1 MEM_stage_inst_dmem_U10760 ( .A1(MEM_stage_inst_dmem_ram_873), .A2(MEM_stage_inst_dmem_n14110), .ZN(MEM_stage_inst_dmem_n14093) );
NAND2_X1 MEM_stage_inst_dmem_U10759 ( .A1(MEM_stage_inst_dmem_n14091), .A2(MEM_stage_inst_dmem_n14090), .ZN(MEM_stage_inst_dmem_n12197) );
NAND2_X1 MEM_stage_inst_dmem_U10758 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n14111), .ZN(MEM_stage_inst_dmem_n14090) );
NAND2_X1 MEM_stage_inst_dmem_U10757 ( .A1(MEM_stage_inst_dmem_ram_874), .A2(MEM_stage_inst_dmem_n14110), .ZN(MEM_stage_inst_dmem_n14091) );
NAND2_X1 MEM_stage_inst_dmem_U10756 ( .A1(MEM_stage_inst_dmem_n14089), .A2(MEM_stage_inst_dmem_n14088), .ZN(MEM_stage_inst_dmem_n12198) );
NAND2_X1 MEM_stage_inst_dmem_U10755 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n14111), .ZN(MEM_stage_inst_dmem_n14088) );
NAND2_X1 MEM_stage_inst_dmem_U10754 ( .A1(MEM_stage_inst_dmem_ram_875), .A2(MEM_stage_inst_dmem_n14110), .ZN(MEM_stage_inst_dmem_n14089) );
NAND2_X1 MEM_stage_inst_dmem_U10753 ( .A1(MEM_stage_inst_dmem_n14087), .A2(MEM_stage_inst_dmem_n14086), .ZN(MEM_stage_inst_dmem_n12199) );
NAND2_X1 MEM_stage_inst_dmem_U10752 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n14111), .ZN(MEM_stage_inst_dmem_n14086) );
NAND2_X1 MEM_stage_inst_dmem_U10751 ( .A1(MEM_stage_inst_dmem_ram_876), .A2(MEM_stage_inst_dmem_n14110), .ZN(MEM_stage_inst_dmem_n14087) );
NAND2_X1 MEM_stage_inst_dmem_U10750 ( .A1(MEM_stage_inst_dmem_n14085), .A2(MEM_stage_inst_dmem_n14084), .ZN(MEM_stage_inst_dmem_n12200) );
NAND2_X1 MEM_stage_inst_dmem_U10749 ( .A1(MEM_stage_inst_dmem_n19242), .A2(MEM_stage_inst_dmem_n14111), .ZN(MEM_stage_inst_dmem_n14084) );
NAND2_X1 MEM_stage_inst_dmem_U10748 ( .A1(MEM_stage_inst_dmem_ram_877), .A2(MEM_stage_inst_dmem_n14110), .ZN(MEM_stage_inst_dmem_n14085) );
NAND2_X1 MEM_stage_inst_dmem_U10747 ( .A1(MEM_stage_inst_dmem_n14083), .A2(MEM_stage_inst_dmem_n14082), .ZN(MEM_stage_inst_dmem_n12201) );
NAND2_X1 MEM_stage_inst_dmem_U10746 ( .A1(MEM_stage_inst_dmem_n115), .A2(MEM_stage_inst_dmem_n14111), .ZN(MEM_stage_inst_dmem_n14082) );
NAND2_X1 MEM_stage_inst_dmem_U10745 ( .A1(MEM_stage_inst_dmem_ram_878), .A2(MEM_stage_inst_dmem_n14110), .ZN(MEM_stage_inst_dmem_n14083) );
NAND2_X1 MEM_stage_inst_dmem_U10744 ( .A1(MEM_stage_inst_dmem_n14081), .A2(MEM_stage_inst_dmem_n14080), .ZN(MEM_stage_inst_dmem_n12202) );
NAND2_X1 MEM_stage_inst_dmem_U10743 ( .A1(MEM_stage_inst_dmem_n16343), .A2(MEM_stage_inst_dmem_n14111), .ZN(MEM_stage_inst_dmem_n14080) );
INV_X1 MEM_stage_inst_dmem_U10742 ( .A(MEM_stage_inst_dmem_n14110), .ZN(MEM_stage_inst_dmem_n14111) );
NAND2_X1 MEM_stage_inst_dmem_U10741 ( .A1(MEM_stage_inst_dmem_ram_879), .A2(MEM_stage_inst_dmem_n14110), .ZN(MEM_stage_inst_dmem_n14081) );
NAND2_X1 MEM_stage_inst_dmem_U10740 ( .A1(MEM_stage_inst_dmem_n21249), .A2(MEM_stage_inst_dmem_n14284), .ZN(MEM_stage_inst_dmem_n14110) );
NAND2_X1 MEM_stage_inst_dmem_U10739 ( .A1(MEM_stage_inst_dmem_n14079), .A2(MEM_stage_inst_dmem_n14078), .ZN(MEM_stage_inst_dmem_n12203) );
NAND2_X1 MEM_stage_inst_dmem_U10738 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n14077), .ZN(MEM_stage_inst_dmem_n14078) );
NAND2_X1 MEM_stage_inst_dmem_U10737 ( .A1(MEM_stage_inst_dmem_ram_880), .A2(MEM_stage_inst_dmem_n14076), .ZN(MEM_stage_inst_dmem_n14079) );
NAND2_X1 MEM_stage_inst_dmem_U10736 ( .A1(MEM_stage_inst_dmem_n14075), .A2(MEM_stage_inst_dmem_n14074), .ZN(MEM_stage_inst_dmem_n12204) );
NAND2_X1 MEM_stage_inst_dmem_U10735 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n14077), .ZN(MEM_stage_inst_dmem_n14074) );
NAND2_X1 MEM_stage_inst_dmem_U10734 ( .A1(MEM_stage_inst_dmem_ram_881), .A2(MEM_stage_inst_dmem_n14076), .ZN(MEM_stage_inst_dmem_n14075) );
NAND2_X1 MEM_stage_inst_dmem_U10733 ( .A1(MEM_stage_inst_dmem_n14073), .A2(MEM_stage_inst_dmem_n14072), .ZN(MEM_stage_inst_dmem_n12205) );
NAND2_X1 MEM_stage_inst_dmem_U10732 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n14077), .ZN(MEM_stage_inst_dmem_n14072) );
NAND2_X1 MEM_stage_inst_dmem_U10731 ( .A1(MEM_stage_inst_dmem_ram_882), .A2(MEM_stage_inst_dmem_n14076), .ZN(MEM_stage_inst_dmem_n14073) );
NAND2_X1 MEM_stage_inst_dmem_U10730 ( .A1(MEM_stage_inst_dmem_n14071), .A2(MEM_stage_inst_dmem_n14070), .ZN(MEM_stage_inst_dmem_n12206) );
NAND2_X1 MEM_stage_inst_dmem_U10729 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n14077), .ZN(MEM_stage_inst_dmem_n14070) );
NAND2_X1 MEM_stage_inst_dmem_U10728 ( .A1(MEM_stage_inst_dmem_ram_883), .A2(MEM_stage_inst_dmem_n14076), .ZN(MEM_stage_inst_dmem_n14071) );
NAND2_X1 MEM_stage_inst_dmem_U10727 ( .A1(MEM_stage_inst_dmem_n14069), .A2(MEM_stage_inst_dmem_n14068), .ZN(MEM_stage_inst_dmem_n12207) );
NAND2_X1 MEM_stage_inst_dmem_U10726 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n14077), .ZN(MEM_stage_inst_dmem_n14068) );
NAND2_X1 MEM_stage_inst_dmem_U10725 ( .A1(MEM_stage_inst_dmem_ram_884), .A2(MEM_stage_inst_dmem_n14076), .ZN(MEM_stage_inst_dmem_n14069) );
NAND2_X1 MEM_stage_inst_dmem_U10724 ( .A1(MEM_stage_inst_dmem_n14067), .A2(MEM_stage_inst_dmem_n14066), .ZN(MEM_stage_inst_dmem_n12208) );
NAND2_X1 MEM_stage_inst_dmem_U10723 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n14077), .ZN(MEM_stage_inst_dmem_n14066) );
NAND2_X1 MEM_stage_inst_dmem_U10722 ( .A1(MEM_stage_inst_dmem_ram_885), .A2(MEM_stage_inst_dmem_n14076), .ZN(MEM_stage_inst_dmem_n14067) );
NAND2_X1 MEM_stage_inst_dmem_U10721 ( .A1(MEM_stage_inst_dmem_n14065), .A2(MEM_stage_inst_dmem_n14064), .ZN(MEM_stage_inst_dmem_n12209) );
NAND2_X1 MEM_stage_inst_dmem_U10720 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n14077), .ZN(MEM_stage_inst_dmem_n14064) );
NAND2_X1 MEM_stage_inst_dmem_U10719 ( .A1(MEM_stage_inst_dmem_ram_886), .A2(MEM_stage_inst_dmem_n14076), .ZN(MEM_stage_inst_dmem_n14065) );
NAND2_X1 MEM_stage_inst_dmem_U10718 ( .A1(MEM_stage_inst_dmem_n14063), .A2(MEM_stage_inst_dmem_n14062), .ZN(MEM_stage_inst_dmem_n12210) );
NAND2_X1 MEM_stage_inst_dmem_U10717 ( .A1(MEM_stage_inst_dmem_n18), .A2(MEM_stage_inst_dmem_n14077), .ZN(MEM_stage_inst_dmem_n14062) );
NAND2_X1 MEM_stage_inst_dmem_U10716 ( .A1(MEM_stage_inst_dmem_ram_887), .A2(MEM_stage_inst_dmem_n14076), .ZN(MEM_stage_inst_dmem_n14063) );
NAND2_X1 MEM_stage_inst_dmem_U10715 ( .A1(MEM_stage_inst_dmem_n14061), .A2(MEM_stage_inst_dmem_n14060), .ZN(MEM_stage_inst_dmem_n12211) );
NAND2_X1 MEM_stage_inst_dmem_U10714 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n14077), .ZN(MEM_stage_inst_dmem_n14060) );
NAND2_X1 MEM_stage_inst_dmem_U10713 ( .A1(MEM_stage_inst_dmem_ram_888), .A2(MEM_stage_inst_dmem_n14076), .ZN(MEM_stage_inst_dmem_n14061) );
NAND2_X1 MEM_stage_inst_dmem_U10712 ( .A1(MEM_stage_inst_dmem_n14059), .A2(MEM_stage_inst_dmem_n14058), .ZN(MEM_stage_inst_dmem_n12212) );
NAND2_X1 MEM_stage_inst_dmem_U10711 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n14077), .ZN(MEM_stage_inst_dmem_n14058) );
NAND2_X1 MEM_stage_inst_dmem_U10710 ( .A1(MEM_stage_inst_dmem_ram_889), .A2(MEM_stage_inst_dmem_n14076), .ZN(MEM_stage_inst_dmem_n14059) );
NAND2_X1 MEM_stage_inst_dmem_U10709 ( .A1(MEM_stage_inst_dmem_n14057), .A2(MEM_stage_inst_dmem_n14056), .ZN(MEM_stage_inst_dmem_n12213) );
NAND2_X1 MEM_stage_inst_dmem_U10708 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n14077), .ZN(MEM_stage_inst_dmem_n14056) );
NAND2_X1 MEM_stage_inst_dmem_U10707 ( .A1(MEM_stage_inst_dmem_ram_890), .A2(MEM_stage_inst_dmem_n14076), .ZN(MEM_stage_inst_dmem_n14057) );
NAND2_X1 MEM_stage_inst_dmem_U10706 ( .A1(MEM_stage_inst_dmem_n14055), .A2(MEM_stage_inst_dmem_n14054), .ZN(MEM_stage_inst_dmem_n12214) );
NAND2_X1 MEM_stage_inst_dmem_U10705 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n14077), .ZN(MEM_stage_inst_dmem_n14054) );
NAND2_X1 MEM_stage_inst_dmem_U10704 ( .A1(MEM_stage_inst_dmem_ram_891), .A2(MEM_stage_inst_dmem_n14076), .ZN(MEM_stage_inst_dmem_n14055) );
NAND2_X1 MEM_stage_inst_dmem_U10703 ( .A1(MEM_stage_inst_dmem_n14053), .A2(MEM_stage_inst_dmem_n14052), .ZN(MEM_stage_inst_dmem_n12215) );
NAND2_X1 MEM_stage_inst_dmem_U10702 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n14077), .ZN(MEM_stage_inst_dmem_n14052) );
NAND2_X1 MEM_stage_inst_dmem_U10701 ( .A1(MEM_stage_inst_dmem_ram_892), .A2(MEM_stage_inst_dmem_n14076), .ZN(MEM_stage_inst_dmem_n14053) );
NAND2_X1 MEM_stage_inst_dmem_U10700 ( .A1(MEM_stage_inst_dmem_n14051), .A2(MEM_stage_inst_dmem_n14050), .ZN(MEM_stage_inst_dmem_n12216) );
NAND2_X1 MEM_stage_inst_dmem_U10699 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n14077), .ZN(MEM_stage_inst_dmem_n14050) );
NAND2_X1 MEM_stage_inst_dmem_U10698 ( .A1(MEM_stage_inst_dmem_ram_893), .A2(MEM_stage_inst_dmem_n14076), .ZN(MEM_stage_inst_dmem_n14051) );
NAND2_X1 MEM_stage_inst_dmem_U10697 ( .A1(MEM_stage_inst_dmem_n14049), .A2(MEM_stage_inst_dmem_n14048), .ZN(MEM_stage_inst_dmem_n12217) );
NAND2_X1 MEM_stage_inst_dmem_U10696 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n14077), .ZN(MEM_stage_inst_dmem_n14048) );
NAND2_X1 MEM_stage_inst_dmem_U10695 ( .A1(MEM_stage_inst_dmem_ram_894), .A2(MEM_stage_inst_dmem_n14076), .ZN(MEM_stage_inst_dmem_n14049) );
NAND2_X1 MEM_stage_inst_dmem_U10694 ( .A1(MEM_stage_inst_dmem_n14047), .A2(MEM_stage_inst_dmem_n14046), .ZN(MEM_stage_inst_dmem_n12218) );
NAND2_X1 MEM_stage_inst_dmem_U10693 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n14077), .ZN(MEM_stage_inst_dmem_n14046) );
INV_X1 MEM_stage_inst_dmem_U10692 ( .A(MEM_stage_inst_dmem_n14076), .ZN(MEM_stage_inst_dmem_n14077) );
NAND2_X1 MEM_stage_inst_dmem_U10691 ( .A1(MEM_stage_inst_dmem_ram_895), .A2(MEM_stage_inst_dmem_n14076), .ZN(MEM_stage_inst_dmem_n14047) );
NAND2_X1 MEM_stage_inst_dmem_U10690 ( .A1(MEM_stage_inst_dmem_n21214), .A2(MEM_stage_inst_dmem_n14284), .ZN(MEM_stage_inst_dmem_n14076) );
NAND2_X1 MEM_stage_inst_dmem_U10689 ( .A1(MEM_stage_inst_dmem_n14045), .A2(MEM_stage_inst_dmem_n14044), .ZN(MEM_stage_inst_dmem_n12219) );
NAND2_X1 MEM_stage_inst_dmem_U10688 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n14043), .ZN(MEM_stage_inst_dmem_n14044) );
NAND2_X1 MEM_stage_inst_dmem_U10687 ( .A1(MEM_stage_inst_dmem_ram_896), .A2(MEM_stage_inst_dmem_n14042), .ZN(MEM_stage_inst_dmem_n14045) );
NAND2_X1 MEM_stage_inst_dmem_U10686 ( .A1(MEM_stage_inst_dmem_n14041), .A2(MEM_stage_inst_dmem_n14040), .ZN(MEM_stage_inst_dmem_n12220) );
NAND2_X1 MEM_stage_inst_dmem_U10685 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n14043), .ZN(MEM_stage_inst_dmem_n14040) );
NAND2_X1 MEM_stage_inst_dmem_U10684 ( .A1(MEM_stage_inst_dmem_ram_897), .A2(MEM_stage_inst_dmem_n14042), .ZN(MEM_stage_inst_dmem_n14041) );
NAND2_X1 MEM_stage_inst_dmem_U10683 ( .A1(MEM_stage_inst_dmem_n14039), .A2(MEM_stage_inst_dmem_n14038), .ZN(MEM_stage_inst_dmem_n12221) );
NAND2_X1 MEM_stage_inst_dmem_U10682 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n14043), .ZN(MEM_stage_inst_dmem_n14038) );
NAND2_X1 MEM_stage_inst_dmem_U10681 ( .A1(MEM_stage_inst_dmem_ram_898), .A2(MEM_stage_inst_dmem_n14042), .ZN(MEM_stage_inst_dmem_n14039) );
NAND2_X1 MEM_stage_inst_dmem_U10680 ( .A1(MEM_stage_inst_dmem_n14037), .A2(MEM_stage_inst_dmem_n14036), .ZN(MEM_stage_inst_dmem_n12222) );
NAND2_X1 MEM_stage_inst_dmem_U10679 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n14043), .ZN(MEM_stage_inst_dmem_n14036) );
NAND2_X1 MEM_stage_inst_dmem_U10678 ( .A1(MEM_stage_inst_dmem_ram_899), .A2(MEM_stage_inst_dmem_n14042), .ZN(MEM_stage_inst_dmem_n14037) );
NAND2_X1 MEM_stage_inst_dmem_U10677 ( .A1(MEM_stage_inst_dmem_n14035), .A2(MEM_stage_inst_dmem_n14034), .ZN(MEM_stage_inst_dmem_n12223) );
NAND2_X1 MEM_stage_inst_dmem_U10676 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n14043), .ZN(MEM_stage_inst_dmem_n14034) );
NAND2_X1 MEM_stage_inst_dmem_U10675 ( .A1(MEM_stage_inst_dmem_ram_900), .A2(MEM_stage_inst_dmem_n14042), .ZN(MEM_stage_inst_dmem_n14035) );
NAND2_X1 MEM_stage_inst_dmem_U10674 ( .A1(MEM_stage_inst_dmem_n14033), .A2(MEM_stage_inst_dmem_n14032), .ZN(MEM_stage_inst_dmem_n12224) );
NAND2_X1 MEM_stage_inst_dmem_U10673 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n14043), .ZN(MEM_stage_inst_dmem_n14032) );
NAND2_X1 MEM_stage_inst_dmem_U10672 ( .A1(MEM_stage_inst_dmem_ram_901), .A2(MEM_stage_inst_dmem_n14042), .ZN(MEM_stage_inst_dmem_n14033) );
NAND2_X1 MEM_stage_inst_dmem_U10671 ( .A1(MEM_stage_inst_dmem_n14031), .A2(MEM_stage_inst_dmem_n14030), .ZN(MEM_stage_inst_dmem_n12225) );
NAND2_X1 MEM_stage_inst_dmem_U10670 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n14043), .ZN(MEM_stage_inst_dmem_n14030) );
NAND2_X1 MEM_stage_inst_dmem_U10669 ( .A1(MEM_stage_inst_dmem_ram_902), .A2(MEM_stage_inst_dmem_n14042), .ZN(MEM_stage_inst_dmem_n14031) );
NAND2_X1 MEM_stage_inst_dmem_U10668 ( .A1(MEM_stage_inst_dmem_n14029), .A2(MEM_stage_inst_dmem_n14028), .ZN(MEM_stage_inst_dmem_n12226) );
NAND2_X1 MEM_stage_inst_dmem_U10667 ( .A1(MEM_stage_inst_dmem_n17), .A2(MEM_stage_inst_dmem_n14043), .ZN(MEM_stage_inst_dmem_n14028) );
NAND2_X1 MEM_stage_inst_dmem_U10666 ( .A1(MEM_stage_inst_dmem_ram_903), .A2(MEM_stage_inst_dmem_n14042), .ZN(MEM_stage_inst_dmem_n14029) );
NAND2_X1 MEM_stage_inst_dmem_U10665 ( .A1(MEM_stage_inst_dmem_n14027), .A2(MEM_stage_inst_dmem_n14026), .ZN(MEM_stage_inst_dmem_n12227) );
NAND2_X1 MEM_stage_inst_dmem_U10664 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n14043), .ZN(MEM_stage_inst_dmem_n14026) );
NAND2_X1 MEM_stage_inst_dmem_U10663 ( .A1(MEM_stage_inst_dmem_ram_904), .A2(MEM_stage_inst_dmem_n14042), .ZN(MEM_stage_inst_dmem_n14027) );
NAND2_X1 MEM_stage_inst_dmem_U10662 ( .A1(MEM_stage_inst_dmem_n14025), .A2(MEM_stage_inst_dmem_n14024), .ZN(MEM_stage_inst_dmem_n12228) );
NAND2_X1 MEM_stage_inst_dmem_U10661 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n14043), .ZN(MEM_stage_inst_dmem_n14024) );
NAND2_X1 MEM_stage_inst_dmem_U10660 ( .A1(MEM_stage_inst_dmem_ram_905), .A2(MEM_stage_inst_dmem_n14042), .ZN(MEM_stage_inst_dmem_n14025) );
NAND2_X1 MEM_stage_inst_dmem_U10659 ( .A1(MEM_stage_inst_dmem_n14023), .A2(MEM_stage_inst_dmem_n14022), .ZN(MEM_stage_inst_dmem_n12229) );
NAND2_X1 MEM_stage_inst_dmem_U10658 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n14043), .ZN(MEM_stage_inst_dmem_n14022) );
NAND2_X1 MEM_stage_inst_dmem_U10657 ( .A1(MEM_stage_inst_dmem_ram_906), .A2(MEM_stage_inst_dmem_n14042), .ZN(MEM_stage_inst_dmem_n14023) );
NAND2_X1 MEM_stage_inst_dmem_U10656 ( .A1(MEM_stage_inst_dmem_n14021), .A2(MEM_stage_inst_dmem_n14020), .ZN(MEM_stage_inst_dmem_n12230) );
NAND2_X1 MEM_stage_inst_dmem_U10655 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n14043), .ZN(MEM_stage_inst_dmem_n14020) );
NAND2_X1 MEM_stage_inst_dmem_U10654 ( .A1(MEM_stage_inst_dmem_ram_907), .A2(MEM_stage_inst_dmem_n14042), .ZN(MEM_stage_inst_dmem_n14021) );
NAND2_X1 MEM_stage_inst_dmem_U10653 ( .A1(MEM_stage_inst_dmem_n14019), .A2(MEM_stage_inst_dmem_n14018), .ZN(MEM_stage_inst_dmem_n12231) );
NAND2_X1 MEM_stage_inst_dmem_U10652 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n14043), .ZN(MEM_stage_inst_dmem_n14018) );
NAND2_X1 MEM_stage_inst_dmem_U10651 ( .A1(MEM_stage_inst_dmem_ram_908), .A2(MEM_stage_inst_dmem_n14042), .ZN(MEM_stage_inst_dmem_n14019) );
NAND2_X1 MEM_stage_inst_dmem_U10650 ( .A1(MEM_stage_inst_dmem_n14017), .A2(MEM_stage_inst_dmem_n14016), .ZN(MEM_stage_inst_dmem_n12232) );
NAND2_X1 MEM_stage_inst_dmem_U10649 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n14043), .ZN(MEM_stage_inst_dmem_n14016) );
NAND2_X1 MEM_stage_inst_dmem_U10648 ( .A1(MEM_stage_inst_dmem_ram_909), .A2(MEM_stage_inst_dmem_n14042), .ZN(MEM_stage_inst_dmem_n14017) );
NAND2_X1 MEM_stage_inst_dmem_U10647 ( .A1(MEM_stage_inst_dmem_n14015), .A2(MEM_stage_inst_dmem_n14014), .ZN(MEM_stage_inst_dmem_n12233) );
NAND2_X1 MEM_stage_inst_dmem_U10646 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n14043), .ZN(MEM_stage_inst_dmem_n14014) );
NAND2_X1 MEM_stage_inst_dmem_U10645 ( .A1(MEM_stage_inst_dmem_ram_910), .A2(MEM_stage_inst_dmem_n14042), .ZN(MEM_stage_inst_dmem_n14015) );
NAND2_X1 MEM_stage_inst_dmem_U10644 ( .A1(MEM_stage_inst_dmem_n14013), .A2(MEM_stage_inst_dmem_n14012), .ZN(MEM_stage_inst_dmem_n12234) );
NAND2_X1 MEM_stage_inst_dmem_U10643 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n14043), .ZN(MEM_stage_inst_dmem_n14012) );
INV_X1 MEM_stage_inst_dmem_U10642 ( .A(MEM_stage_inst_dmem_n14042), .ZN(MEM_stage_inst_dmem_n14043) );
NAND2_X1 MEM_stage_inst_dmem_U10641 ( .A1(MEM_stage_inst_dmem_ram_911), .A2(MEM_stage_inst_dmem_n14042), .ZN(MEM_stage_inst_dmem_n14013) );
NAND2_X1 MEM_stage_inst_dmem_U10640 ( .A1(MEM_stage_inst_dmem_n21179), .A2(MEM_stage_inst_dmem_n14284), .ZN(MEM_stage_inst_dmem_n14042) );
NAND2_X1 MEM_stage_inst_dmem_U10639 ( .A1(MEM_stage_inst_dmem_n14011), .A2(MEM_stage_inst_dmem_n14010), .ZN(MEM_stage_inst_dmem_n12235) );
NAND2_X1 MEM_stage_inst_dmem_U10638 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n14009), .ZN(MEM_stage_inst_dmem_n14010) );
NAND2_X1 MEM_stage_inst_dmem_U10637 ( .A1(MEM_stage_inst_dmem_ram_912), .A2(MEM_stage_inst_dmem_n14008), .ZN(MEM_stage_inst_dmem_n14011) );
NAND2_X1 MEM_stage_inst_dmem_U10636 ( .A1(MEM_stage_inst_dmem_n14007), .A2(MEM_stage_inst_dmem_n14006), .ZN(MEM_stage_inst_dmem_n12236) );
NAND2_X1 MEM_stage_inst_dmem_U10635 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n14009), .ZN(MEM_stage_inst_dmem_n14006) );
NAND2_X1 MEM_stage_inst_dmem_U10634 ( .A1(MEM_stage_inst_dmem_ram_913), .A2(MEM_stage_inst_dmem_n14008), .ZN(MEM_stage_inst_dmem_n14007) );
NAND2_X1 MEM_stage_inst_dmem_U10633 ( .A1(MEM_stage_inst_dmem_n14005), .A2(MEM_stage_inst_dmem_n14004), .ZN(MEM_stage_inst_dmem_n12237) );
NAND2_X1 MEM_stage_inst_dmem_U10632 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n14009), .ZN(MEM_stage_inst_dmem_n14004) );
NAND2_X1 MEM_stage_inst_dmem_U10631 ( .A1(MEM_stage_inst_dmem_ram_914), .A2(MEM_stage_inst_dmem_n14008), .ZN(MEM_stage_inst_dmem_n14005) );
NAND2_X1 MEM_stage_inst_dmem_U10630 ( .A1(MEM_stage_inst_dmem_n14003), .A2(MEM_stage_inst_dmem_n14002), .ZN(MEM_stage_inst_dmem_n12238) );
NAND2_X1 MEM_stage_inst_dmem_U10629 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n14009), .ZN(MEM_stage_inst_dmem_n14002) );
NAND2_X1 MEM_stage_inst_dmem_U10628 ( .A1(MEM_stage_inst_dmem_ram_915), .A2(MEM_stage_inst_dmem_n14008), .ZN(MEM_stage_inst_dmem_n14003) );
NAND2_X1 MEM_stage_inst_dmem_U10627 ( .A1(MEM_stage_inst_dmem_n14001), .A2(MEM_stage_inst_dmem_n14000), .ZN(MEM_stage_inst_dmem_n12239) );
NAND2_X1 MEM_stage_inst_dmem_U10626 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n14009), .ZN(MEM_stage_inst_dmem_n14000) );
NAND2_X1 MEM_stage_inst_dmem_U10625 ( .A1(MEM_stage_inst_dmem_ram_916), .A2(MEM_stage_inst_dmem_n14008), .ZN(MEM_stage_inst_dmem_n14001) );
NAND2_X1 MEM_stage_inst_dmem_U10624 ( .A1(MEM_stage_inst_dmem_n13999), .A2(MEM_stage_inst_dmem_n13998), .ZN(MEM_stage_inst_dmem_n12240) );
NAND2_X1 MEM_stage_inst_dmem_U10623 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n14009), .ZN(MEM_stage_inst_dmem_n13998) );
NAND2_X1 MEM_stage_inst_dmem_U10622 ( .A1(MEM_stage_inst_dmem_ram_917), .A2(MEM_stage_inst_dmem_n14008), .ZN(MEM_stage_inst_dmem_n13999) );
NAND2_X1 MEM_stage_inst_dmem_U10621 ( .A1(MEM_stage_inst_dmem_n13997), .A2(MEM_stage_inst_dmem_n13996), .ZN(MEM_stage_inst_dmem_n12241) );
NAND2_X1 MEM_stage_inst_dmem_U10620 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n14009), .ZN(MEM_stage_inst_dmem_n13996) );
NAND2_X1 MEM_stage_inst_dmem_U10619 ( .A1(MEM_stage_inst_dmem_ram_918), .A2(MEM_stage_inst_dmem_n14008), .ZN(MEM_stage_inst_dmem_n13997) );
NAND2_X1 MEM_stage_inst_dmem_U10618 ( .A1(MEM_stage_inst_dmem_n13995), .A2(MEM_stage_inst_dmem_n13994), .ZN(MEM_stage_inst_dmem_n12242) );
NAND2_X1 MEM_stage_inst_dmem_U10617 ( .A1(MEM_stage_inst_dmem_n18), .A2(MEM_stage_inst_dmem_n14009), .ZN(MEM_stage_inst_dmem_n13994) );
NAND2_X1 MEM_stage_inst_dmem_U10616 ( .A1(MEM_stage_inst_dmem_ram_919), .A2(MEM_stage_inst_dmem_n14008), .ZN(MEM_stage_inst_dmem_n13995) );
NAND2_X1 MEM_stage_inst_dmem_U10615 ( .A1(MEM_stage_inst_dmem_n13993), .A2(MEM_stage_inst_dmem_n13992), .ZN(MEM_stage_inst_dmem_n12243) );
NAND2_X1 MEM_stage_inst_dmem_U10614 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n14009), .ZN(MEM_stage_inst_dmem_n13992) );
NAND2_X1 MEM_stage_inst_dmem_U10613 ( .A1(MEM_stage_inst_dmem_ram_920), .A2(MEM_stage_inst_dmem_n14008), .ZN(MEM_stage_inst_dmem_n13993) );
NAND2_X1 MEM_stage_inst_dmem_U10612 ( .A1(MEM_stage_inst_dmem_n13991), .A2(MEM_stage_inst_dmem_n13990), .ZN(MEM_stage_inst_dmem_n12244) );
NAND2_X1 MEM_stage_inst_dmem_U10611 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n14009), .ZN(MEM_stage_inst_dmem_n13990) );
NAND2_X1 MEM_stage_inst_dmem_U10610 ( .A1(MEM_stage_inst_dmem_ram_921), .A2(MEM_stage_inst_dmem_n14008), .ZN(MEM_stage_inst_dmem_n13991) );
NAND2_X1 MEM_stage_inst_dmem_U10609 ( .A1(MEM_stage_inst_dmem_n13989), .A2(MEM_stage_inst_dmem_n13988), .ZN(MEM_stage_inst_dmem_n12245) );
NAND2_X1 MEM_stage_inst_dmem_U10608 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n14009), .ZN(MEM_stage_inst_dmem_n13988) );
NAND2_X1 MEM_stage_inst_dmem_U10607 ( .A1(MEM_stage_inst_dmem_ram_922), .A2(MEM_stage_inst_dmem_n14008), .ZN(MEM_stage_inst_dmem_n13989) );
NAND2_X1 MEM_stage_inst_dmem_U10606 ( .A1(MEM_stage_inst_dmem_n13987), .A2(MEM_stage_inst_dmem_n13986), .ZN(MEM_stage_inst_dmem_n12246) );
NAND2_X1 MEM_stage_inst_dmem_U10605 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n14009), .ZN(MEM_stage_inst_dmem_n13986) );
NAND2_X1 MEM_stage_inst_dmem_U10604 ( .A1(MEM_stage_inst_dmem_ram_923), .A2(MEM_stage_inst_dmem_n14008), .ZN(MEM_stage_inst_dmem_n13987) );
NAND2_X1 MEM_stage_inst_dmem_U10603 ( .A1(MEM_stage_inst_dmem_n13985), .A2(MEM_stage_inst_dmem_n13984), .ZN(MEM_stage_inst_dmem_n12247) );
NAND2_X1 MEM_stage_inst_dmem_U10602 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n14009), .ZN(MEM_stage_inst_dmem_n13984) );
NAND2_X1 MEM_stage_inst_dmem_U10601 ( .A1(MEM_stage_inst_dmem_ram_924), .A2(MEM_stage_inst_dmem_n14008), .ZN(MEM_stage_inst_dmem_n13985) );
NAND2_X1 MEM_stage_inst_dmem_U10600 ( .A1(MEM_stage_inst_dmem_n13983), .A2(MEM_stage_inst_dmem_n13982), .ZN(MEM_stage_inst_dmem_n12248) );
NAND2_X1 MEM_stage_inst_dmem_U10599 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n14009), .ZN(MEM_stage_inst_dmem_n13982) );
NAND2_X1 MEM_stage_inst_dmem_U10598 ( .A1(MEM_stage_inst_dmem_ram_925), .A2(MEM_stage_inst_dmem_n14008), .ZN(MEM_stage_inst_dmem_n13983) );
NAND2_X1 MEM_stage_inst_dmem_U10597 ( .A1(MEM_stage_inst_dmem_n13981), .A2(MEM_stage_inst_dmem_n13980), .ZN(MEM_stage_inst_dmem_n12249) );
NAND2_X1 MEM_stage_inst_dmem_U10596 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n14009), .ZN(MEM_stage_inst_dmem_n13980) );
NAND2_X1 MEM_stage_inst_dmem_U10595 ( .A1(MEM_stage_inst_dmem_ram_926), .A2(MEM_stage_inst_dmem_n14008), .ZN(MEM_stage_inst_dmem_n13981) );
NAND2_X1 MEM_stage_inst_dmem_U10594 ( .A1(MEM_stage_inst_dmem_n13979), .A2(MEM_stage_inst_dmem_n13978), .ZN(MEM_stage_inst_dmem_n12250) );
NAND2_X1 MEM_stage_inst_dmem_U10593 ( .A1(MEM_stage_inst_dmem_n16343), .A2(MEM_stage_inst_dmem_n14009), .ZN(MEM_stage_inst_dmem_n13978) );
INV_X1 MEM_stage_inst_dmem_U10592 ( .A(MEM_stage_inst_dmem_n14008), .ZN(MEM_stage_inst_dmem_n14009) );
NAND2_X1 MEM_stage_inst_dmem_U10591 ( .A1(MEM_stage_inst_dmem_ram_927), .A2(MEM_stage_inst_dmem_n14008), .ZN(MEM_stage_inst_dmem_n13979) );
NAND2_X1 MEM_stage_inst_dmem_U10590 ( .A1(MEM_stage_inst_dmem_n21144), .A2(MEM_stage_inst_dmem_n14284), .ZN(MEM_stage_inst_dmem_n14008) );
NAND2_X1 MEM_stage_inst_dmem_U10589 ( .A1(MEM_stage_inst_dmem_n13977), .A2(MEM_stage_inst_dmem_n13976), .ZN(MEM_stage_inst_dmem_n12251) );
NAND2_X1 MEM_stage_inst_dmem_U10588 ( .A1(MEM_stage_inst_dmem_n15145), .A2(MEM_stage_inst_dmem_n13975), .ZN(MEM_stage_inst_dmem_n13976) );
NAND2_X1 MEM_stage_inst_dmem_U10587 ( .A1(MEM_stage_inst_dmem_ram_928), .A2(MEM_stage_inst_dmem_n13974), .ZN(MEM_stage_inst_dmem_n13977) );
NAND2_X1 MEM_stage_inst_dmem_U10586 ( .A1(MEM_stage_inst_dmem_n13973), .A2(MEM_stage_inst_dmem_n13972), .ZN(MEM_stage_inst_dmem_n12252) );
NAND2_X1 MEM_stage_inst_dmem_U10585 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n13975), .ZN(MEM_stage_inst_dmem_n13972) );
NAND2_X1 MEM_stage_inst_dmem_U10584 ( .A1(MEM_stage_inst_dmem_ram_929), .A2(MEM_stage_inst_dmem_n13974), .ZN(MEM_stage_inst_dmem_n13973) );
NAND2_X1 MEM_stage_inst_dmem_U10583 ( .A1(MEM_stage_inst_dmem_n13971), .A2(MEM_stage_inst_dmem_n13970), .ZN(MEM_stage_inst_dmem_n12253) );
NAND2_X1 MEM_stage_inst_dmem_U10582 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n13975), .ZN(MEM_stage_inst_dmem_n13970) );
NAND2_X1 MEM_stage_inst_dmem_U10581 ( .A1(MEM_stage_inst_dmem_ram_930), .A2(MEM_stage_inst_dmem_n13974), .ZN(MEM_stage_inst_dmem_n13971) );
NAND2_X1 MEM_stage_inst_dmem_U10580 ( .A1(MEM_stage_inst_dmem_n13969), .A2(MEM_stage_inst_dmem_n13968), .ZN(MEM_stage_inst_dmem_n12254) );
NAND2_X1 MEM_stage_inst_dmem_U10579 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n13975), .ZN(MEM_stage_inst_dmem_n13968) );
NAND2_X1 MEM_stage_inst_dmem_U10578 ( .A1(MEM_stage_inst_dmem_ram_931), .A2(MEM_stage_inst_dmem_n13974), .ZN(MEM_stage_inst_dmem_n13969) );
NAND2_X1 MEM_stage_inst_dmem_U10577 ( .A1(MEM_stage_inst_dmem_n13967), .A2(MEM_stage_inst_dmem_n13966), .ZN(MEM_stage_inst_dmem_n12255) );
NAND2_X1 MEM_stage_inst_dmem_U10576 ( .A1(MEM_stage_inst_dmem_n16784), .A2(MEM_stage_inst_dmem_n13975), .ZN(MEM_stage_inst_dmem_n13966) );
NAND2_X1 MEM_stage_inst_dmem_U10575 ( .A1(MEM_stage_inst_dmem_ram_932), .A2(MEM_stage_inst_dmem_n13974), .ZN(MEM_stage_inst_dmem_n13967) );
NAND2_X1 MEM_stage_inst_dmem_U10574 ( .A1(MEM_stage_inst_dmem_n13965), .A2(MEM_stage_inst_dmem_n13964), .ZN(MEM_stage_inst_dmem_n12256) );
NAND2_X1 MEM_stage_inst_dmem_U10573 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n13975), .ZN(MEM_stage_inst_dmem_n13964) );
NAND2_X1 MEM_stage_inst_dmem_U10572 ( .A1(MEM_stage_inst_dmem_ram_933), .A2(MEM_stage_inst_dmem_n13974), .ZN(MEM_stage_inst_dmem_n13965) );
NAND2_X1 MEM_stage_inst_dmem_U10571 ( .A1(MEM_stage_inst_dmem_n13963), .A2(MEM_stage_inst_dmem_n13962), .ZN(MEM_stage_inst_dmem_n12257) );
NAND2_X1 MEM_stage_inst_dmem_U10570 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n13975), .ZN(MEM_stage_inst_dmem_n13962) );
NAND2_X1 MEM_stage_inst_dmem_U10569 ( .A1(MEM_stage_inst_dmem_ram_934), .A2(MEM_stage_inst_dmem_n13974), .ZN(MEM_stage_inst_dmem_n13963) );
NAND2_X1 MEM_stage_inst_dmem_U10568 ( .A1(MEM_stage_inst_dmem_n13961), .A2(MEM_stage_inst_dmem_n13960), .ZN(MEM_stage_inst_dmem_n12258) );
NAND2_X1 MEM_stage_inst_dmem_U10567 ( .A1(MEM_stage_inst_dmem_n17), .A2(MEM_stage_inst_dmem_n13975), .ZN(MEM_stage_inst_dmem_n13960) );
NAND2_X1 MEM_stage_inst_dmem_U10566 ( .A1(MEM_stage_inst_dmem_ram_935), .A2(MEM_stage_inst_dmem_n13974), .ZN(MEM_stage_inst_dmem_n13961) );
NAND2_X1 MEM_stage_inst_dmem_U10565 ( .A1(MEM_stage_inst_dmem_n13959), .A2(MEM_stage_inst_dmem_n13958), .ZN(MEM_stage_inst_dmem_n12259) );
NAND2_X1 MEM_stage_inst_dmem_U10564 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n13975), .ZN(MEM_stage_inst_dmem_n13958) );
NAND2_X1 MEM_stage_inst_dmem_U10563 ( .A1(MEM_stage_inst_dmem_ram_936), .A2(MEM_stage_inst_dmem_n13974), .ZN(MEM_stage_inst_dmem_n13959) );
NAND2_X1 MEM_stage_inst_dmem_U10562 ( .A1(MEM_stage_inst_dmem_n13957), .A2(MEM_stage_inst_dmem_n13956), .ZN(MEM_stage_inst_dmem_n12260) );
NAND2_X1 MEM_stage_inst_dmem_U10561 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n13975), .ZN(MEM_stage_inst_dmem_n13956) );
NAND2_X1 MEM_stage_inst_dmem_U10560 ( .A1(MEM_stage_inst_dmem_ram_937), .A2(MEM_stage_inst_dmem_n13974), .ZN(MEM_stage_inst_dmem_n13957) );
NAND2_X1 MEM_stage_inst_dmem_U10559 ( .A1(MEM_stage_inst_dmem_n13955), .A2(MEM_stage_inst_dmem_n13954), .ZN(MEM_stage_inst_dmem_n12261) );
NAND2_X1 MEM_stage_inst_dmem_U10558 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n13975), .ZN(MEM_stage_inst_dmem_n13954) );
NAND2_X1 MEM_stage_inst_dmem_U10557 ( .A1(MEM_stage_inst_dmem_ram_938), .A2(MEM_stage_inst_dmem_n13974), .ZN(MEM_stage_inst_dmem_n13955) );
NAND2_X1 MEM_stage_inst_dmem_U10556 ( .A1(MEM_stage_inst_dmem_n13953), .A2(MEM_stage_inst_dmem_n13952), .ZN(MEM_stage_inst_dmem_n12262) );
NAND2_X1 MEM_stage_inst_dmem_U10555 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n13975), .ZN(MEM_stage_inst_dmem_n13952) );
NAND2_X1 MEM_stage_inst_dmem_U10554 ( .A1(MEM_stage_inst_dmem_ram_939), .A2(MEM_stage_inst_dmem_n13974), .ZN(MEM_stage_inst_dmem_n13953) );
NAND2_X1 MEM_stage_inst_dmem_U10553 ( .A1(MEM_stage_inst_dmem_n13951), .A2(MEM_stage_inst_dmem_n13950), .ZN(MEM_stage_inst_dmem_n12263) );
NAND2_X1 MEM_stage_inst_dmem_U10552 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n13975), .ZN(MEM_stage_inst_dmem_n13950) );
NAND2_X1 MEM_stage_inst_dmem_U10551 ( .A1(MEM_stage_inst_dmem_ram_940), .A2(MEM_stage_inst_dmem_n13974), .ZN(MEM_stage_inst_dmem_n13951) );
NAND2_X1 MEM_stage_inst_dmem_U10550 ( .A1(MEM_stage_inst_dmem_n13949), .A2(MEM_stage_inst_dmem_n13948), .ZN(MEM_stage_inst_dmem_n12264) );
NAND2_X1 MEM_stage_inst_dmem_U10549 ( .A1(MEM_stage_inst_dmem_n15116), .A2(MEM_stage_inst_dmem_n13975), .ZN(MEM_stage_inst_dmem_n13948) );
NAND2_X1 MEM_stage_inst_dmem_U10548 ( .A1(MEM_stage_inst_dmem_ram_941), .A2(MEM_stage_inst_dmem_n13974), .ZN(MEM_stage_inst_dmem_n13949) );
NAND2_X1 MEM_stage_inst_dmem_U10547 ( .A1(MEM_stage_inst_dmem_n13947), .A2(MEM_stage_inst_dmem_n13946), .ZN(MEM_stage_inst_dmem_n12265) );
NAND2_X1 MEM_stage_inst_dmem_U10546 ( .A1(MEM_stage_inst_dmem_n15113), .A2(MEM_stage_inst_dmem_n13975), .ZN(MEM_stage_inst_dmem_n13946) );
NAND2_X1 MEM_stage_inst_dmem_U10545 ( .A1(MEM_stage_inst_dmem_ram_942), .A2(MEM_stage_inst_dmem_n13974), .ZN(MEM_stage_inst_dmem_n13947) );
NAND2_X1 MEM_stage_inst_dmem_U10544 ( .A1(MEM_stage_inst_dmem_n13945), .A2(MEM_stage_inst_dmem_n13944), .ZN(MEM_stage_inst_dmem_n12266) );
NAND2_X1 MEM_stage_inst_dmem_U10543 ( .A1(MEM_stage_inst_dmem_n14693), .A2(MEM_stage_inst_dmem_n13975), .ZN(MEM_stage_inst_dmem_n13944) );
INV_X1 MEM_stage_inst_dmem_U10542 ( .A(MEM_stage_inst_dmem_n13974), .ZN(MEM_stage_inst_dmem_n13975) );
NAND2_X1 MEM_stage_inst_dmem_U10541 ( .A1(MEM_stage_inst_dmem_ram_943), .A2(MEM_stage_inst_dmem_n13974), .ZN(MEM_stage_inst_dmem_n13945) );
NAND2_X1 MEM_stage_inst_dmem_U10540 ( .A1(MEM_stage_inst_dmem_n21109), .A2(MEM_stage_inst_dmem_n14284), .ZN(MEM_stage_inst_dmem_n13974) );
NAND2_X1 MEM_stage_inst_dmem_U10539 ( .A1(MEM_stage_inst_dmem_n13943), .A2(MEM_stage_inst_dmem_n13942), .ZN(MEM_stage_inst_dmem_n12267) );
NAND2_X1 MEM_stage_inst_dmem_U10538 ( .A1(MEM_stage_inst_dmem_n14732), .A2(MEM_stage_inst_dmem_n13941), .ZN(MEM_stage_inst_dmem_n13942) );
NAND2_X1 MEM_stage_inst_dmem_U10537 ( .A1(MEM_stage_inst_dmem_ram_944), .A2(MEM_stage_inst_dmem_n13940), .ZN(MEM_stage_inst_dmem_n13943) );
NAND2_X1 MEM_stage_inst_dmem_U10536 ( .A1(MEM_stage_inst_dmem_n13939), .A2(MEM_stage_inst_dmem_n13938), .ZN(MEM_stage_inst_dmem_n12268) );
NAND2_X1 MEM_stage_inst_dmem_U10535 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n13941), .ZN(MEM_stage_inst_dmem_n13938) );
NAND2_X1 MEM_stage_inst_dmem_U10534 ( .A1(MEM_stage_inst_dmem_ram_945), .A2(MEM_stage_inst_dmem_n13940), .ZN(MEM_stage_inst_dmem_n13939) );
NAND2_X1 MEM_stage_inst_dmem_U10533 ( .A1(MEM_stage_inst_dmem_n13937), .A2(MEM_stage_inst_dmem_n13936), .ZN(MEM_stage_inst_dmem_n12269) );
NAND2_X1 MEM_stage_inst_dmem_U10532 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n13941), .ZN(MEM_stage_inst_dmem_n13936) );
NAND2_X1 MEM_stage_inst_dmem_U10531 ( .A1(MEM_stage_inst_dmem_ram_946), .A2(MEM_stage_inst_dmem_n13940), .ZN(MEM_stage_inst_dmem_n13937) );
NAND2_X1 MEM_stage_inst_dmem_U10530 ( .A1(MEM_stage_inst_dmem_n13935), .A2(MEM_stage_inst_dmem_n13934), .ZN(MEM_stage_inst_dmem_n12270) );
NAND2_X1 MEM_stage_inst_dmem_U10529 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n13941), .ZN(MEM_stage_inst_dmem_n13934) );
NAND2_X1 MEM_stage_inst_dmem_U10528 ( .A1(MEM_stage_inst_dmem_ram_947), .A2(MEM_stage_inst_dmem_n13940), .ZN(MEM_stage_inst_dmem_n13935) );
NAND2_X1 MEM_stage_inst_dmem_U10527 ( .A1(MEM_stage_inst_dmem_n13933), .A2(MEM_stage_inst_dmem_n13932), .ZN(MEM_stage_inst_dmem_n12271) );
NAND2_X1 MEM_stage_inst_dmem_U10526 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n13941), .ZN(MEM_stage_inst_dmem_n13932) );
NAND2_X1 MEM_stage_inst_dmem_U10525 ( .A1(MEM_stage_inst_dmem_ram_948), .A2(MEM_stage_inst_dmem_n13940), .ZN(MEM_stage_inst_dmem_n13933) );
NAND2_X1 MEM_stage_inst_dmem_U10524 ( .A1(MEM_stage_inst_dmem_n13931), .A2(MEM_stage_inst_dmem_n13930), .ZN(MEM_stage_inst_dmem_n12272) );
NAND2_X1 MEM_stage_inst_dmem_U10523 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n13941), .ZN(MEM_stage_inst_dmem_n13930) );
NAND2_X1 MEM_stage_inst_dmem_U10522 ( .A1(MEM_stage_inst_dmem_ram_949), .A2(MEM_stage_inst_dmem_n13940), .ZN(MEM_stage_inst_dmem_n13931) );
NAND2_X1 MEM_stage_inst_dmem_U10521 ( .A1(MEM_stage_inst_dmem_n13929), .A2(MEM_stage_inst_dmem_n13928), .ZN(MEM_stage_inst_dmem_n12273) );
NAND2_X1 MEM_stage_inst_dmem_U10520 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n13941), .ZN(MEM_stage_inst_dmem_n13928) );
NAND2_X1 MEM_stage_inst_dmem_U10519 ( .A1(MEM_stage_inst_dmem_ram_950), .A2(MEM_stage_inst_dmem_n13940), .ZN(MEM_stage_inst_dmem_n13929) );
NAND2_X1 MEM_stage_inst_dmem_U10518 ( .A1(MEM_stage_inst_dmem_n13927), .A2(MEM_stage_inst_dmem_n13926), .ZN(MEM_stage_inst_dmem_n12274) );
NAND2_X1 MEM_stage_inst_dmem_U10517 ( .A1(MEM_stage_inst_dmem_n18), .A2(MEM_stage_inst_dmem_n13941), .ZN(MEM_stage_inst_dmem_n13926) );
NAND2_X1 MEM_stage_inst_dmem_U10516 ( .A1(MEM_stage_inst_dmem_ram_951), .A2(MEM_stage_inst_dmem_n13940), .ZN(MEM_stage_inst_dmem_n13927) );
NAND2_X1 MEM_stage_inst_dmem_U10515 ( .A1(MEM_stage_inst_dmem_n13925), .A2(MEM_stage_inst_dmem_n13924), .ZN(MEM_stage_inst_dmem_n12275) );
NAND2_X1 MEM_stage_inst_dmem_U10514 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n13941), .ZN(MEM_stage_inst_dmem_n13924) );
NAND2_X1 MEM_stage_inst_dmem_U10513 ( .A1(MEM_stage_inst_dmem_ram_952), .A2(MEM_stage_inst_dmem_n13940), .ZN(MEM_stage_inst_dmem_n13925) );
NAND2_X1 MEM_stage_inst_dmem_U10512 ( .A1(MEM_stage_inst_dmem_n13923), .A2(MEM_stage_inst_dmem_n13922), .ZN(MEM_stage_inst_dmem_n12276) );
NAND2_X1 MEM_stage_inst_dmem_U10511 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n13941), .ZN(MEM_stage_inst_dmem_n13922) );
NAND2_X1 MEM_stage_inst_dmem_U10510 ( .A1(MEM_stage_inst_dmem_ram_953), .A2(MEM_stage_inst_dmem_n13940), .ZN(MEM_stage_inst_dmem_n13923) );
NAND2_X1 MEM_stage_inst_dmem_U10509 ( .A1(MEM_stage_inst_dmem_n13921), .A2(MEM_stage_inst_dmem_n13920), .ZN(MEM_stage_inst_dmem_n12277) );
NAND2_X1 MEM_stage_inst_dmem_U10508 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n13941), .ZN(MEM_stage_inst_dmem_n13920) );
NAND2_X1 MEM_stage_inst_dmem_U10507 ( .A1(MEM_stage_inst_dmem_ram_954), .A2(MEM_stage_inst_dmem_n13940), .ZN(MEM_stage_inst_dmem_n13921) );
NAND2_X1 MEM_stage_inst_dmem_U10506 ( .A1(MEM_stage_inst_dmem_n13919), .A2(MEM_stage_inst_dmem_n13918), .ZN(MEM_stage_inst_dmem_n12278) );
NAND2_X1 MEM_stage_inst_dmem_U10505 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n13941), .ZN(MEM_stage_inst_dmem_n13918) );
NAND2_X1 MEM_stage_inst_dmem_U10504 ( .A1(MEM_stage_inst_dmem_ram_955), .A2(MEM_stage_inst_dmem_n13940), .ZN(MEM_stage_inst_dmem_n13919) );
NAND2_X1 MEM_stage_inst_dmem_U10503 ( .A1(MEM_stage_inst_dmem_n13917), .A2(MEM_stage_inst_dmem_n13916), .ZN(MEM_stage_inst_dmem_n12279) );
NAND2_X1 MEM_stage_inst_dmem_U10502 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n13941), .ZN(MEM_stage_inst_dmem_n13916) );
NAND2_X1 MEM_stage_inst_dmem_U10501 ( .A1(MEM_stage_inst_dmem_ram_956), .A2(MEM_stage_inst_dmem_n13940), .ZN(MEM_stage_inst_dmem_n13917) );
NAND2_X1 MEM_stage_inst_dmem_U10500 ( .A1(MEM_stage_inst_dmem_n13915), .A2(MEM_stage_inst_dmem_n13914), .ZN(MEM_stage_inst_dmem_n12280) );
NAND2_X1 MEM_stage_inst_dmem_U10499 ( .A1(MEM_stage_inst_dmem_n116), .A2(MEM_stage_inst_dmem_n13941), .ZN(MEM_stage_inst_dmem_n13914) );
NAND2_X1 MEM_stage_inst_dmem_U10498 ( .A1(MEM_stage_inst_dmem_ram_957), .A2(MEM_stage_inst_dmem_n13940), .ZN(MEM_stage_inst_dmem_n13915) );
NAND2_X1 MEM_stage_inst_dmem_U10497 ( .A1(MEM_stage_inst_dmem_n13913), .A2(MEM_stage_inst_dmem_n13912), .ZN(MEM_stage_inst_dmem_n12281) );
NAND2_X1 MEM_stage_inst_dmem_U10496 ( .A1(MEM_stage_inst_dmem_n14696), .A2(MEM_stage_inst_dmem_n13941), .ZN(MEM_stage_inst_dmem_n13912) );
NAND2_X1 MEM_stage_inst_dmem_U10495 ( .A1(MEM_stage_inst_dmem_ram_958), .A2(MEM_stage_inst_dmem_n13940), .ZN(MEM_stage_inst_dmem_n13913) );
NAND2_X1 MEM_stage_inst_dmem_U10494 ( .A1(MEM_stage_inst_dmem_n13911), .A2(MEM_stage_inst_dmem_n13910), .ZN(MEM_stage_inst_dmem_n12282) );
NAND2_X1 MEM_stage_inst_dmem_U10493 ( .A1(MEM_stage_inst_dmem_n16343), .A2(MEM_stage_inst_dmem_n13941), .ZN(MEM_stage_inst_dmem_n13910) );
NAND2_X1 MEM_stage_inst_dmem_U10492 ( .A1(MEM_stage_inst_dmem_ram_959), .A2(MEM_stage_inst_dmem_n13940), .ZN(MEM_stage_inst_dmem_n13911) );
NAND2_X1 MEM_stage_inst_dmem_U10491 ( .A1(MEM_stage_inst_dmem_n21074), .A2(MEM_stage_inst_dmem_n14284), .ZN(MEM_stage_inst_dmem_n13940) );
NAND2_X1 MEM_stage_inst_dmem_U10490 ( .A1(MEM_stage_inst_dmem_n13909), .A2(MEM_stage_inst_dmem_n13908), .ZN(MEM_stage_inst_dmem_n12283) );
NAND2_X1 MEM_stage_inst_dmem_U10489 ( .A1(MEM_stage_inst_dmem_n15145), .A2(MEM_stage_inst_dmem_n13907), .ZN(MEM_stage_inst_dmem_n13908) );
NAND2_X1 MEM_stage_inst_dmem_U10488 ( .A1(MEM_stage_inst_dmem_ram_960), .A2(MEM_stage_inst_dmem_n13906), .ZN(MEM_stage_inst_dmem_n13909) );
NAND2_X1 MEM_stage_inst_dmem_U10487 ( .A1(MEM_stage_inst_dmem_n13905), .A2(MEM_stage_inst_dmem_n13904), .ZN(MEM_stage_inst_dmem_n12284) );
NAND2_X1 MEM_stage_inst_dmem_U10486 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n13907), .ZN(MEM_stage_inst_dmem_n13904) );
NAND2_X1 MEM_stage_inst_dmem_U10485 ( .A1(MEM_stage_inst_dmem_ram_961), .A2(MEM_stage_inst_dmem_n13906), .ZN(MEM_stage_inst_dmem_n13905) );
NAND2_X1 MEM_stage_inst_dmem_U10484 ( .A1(MEM_stage_inst_dmem_n13902), .A2(MEM_stage_inst_dmem_n13901), .ZN(MEM_stage_inst_dmem_n12285) );
NAND2_X1 MEM_stage_inst_dmem_U10483 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n13907), .ZN(MEM_stage_inst_dmem_n13901) );
NAND2_X1 MEM_stage_inst_dmem_U10482 ( .A1(MEM_stage_inst_dmem_ram_962), .A2(MEM_stage_inst_dmem_n13906), .ZN(MEM_stage_inst_dmem_n13902) );
NAND2_X1 MEM_stage_inst_dmem_U10481 ( .A1(MEM_stage_inst_dmem_n13899), .A2(MEM_stage_inst_dmem_n13898), .ZN(MEM_stage_inst_dmem_n12286) );
NAND2_X1 MEM_stage_inst_dmem_U10480 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n13907), .ZN(MEM_stage_inst_dmem_n13898) );
NAND2_X1 MEM_stage_inst_dmem_U10479 ( .A1(MEM_stage_inst_dmem_ram_963), .A2(MEM_stage_inst_dmem_n13906), .ZN(MEM_stage_inst_dmem_n13899) );
NAND2_X1 MEM_stage_inst_dmem_U10478 ( .A1(MEM_stage_inst_dmem_n13896), .A2(MEM_stage_inst_dmem_n13895), .ZN(MEM_stage_inst_dmem_n12287) );
NAND2_X1 MEM_stage_inst_dmem_U10477 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n13907), .ZN(MEM_stage_inst_dmem_n13895) );
NAND2_X1 MEM_stage_inst_dmem_U10476 ( .A1(MEM_stage_inst_dmem_ram_964), .A2(MEM_stage_inst_dmem_n13906), .ZN(MEM_stage_inst_dmem_n13896) );
NAND2_X1 MEM_stage_inst_dmem_U10475 ( .A1(MEM_stage_inst_dmem_n13894), .A2(MEM_stage_inst_dmem_n13893), .ZN(MEM_stage_inst_dmem_n12288) );
NAND2_X1 MEM_stage_inst_dmem_U10474 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n13907), .ZN(MEM_stage_inst_dmem_n13893) );
NAND2_X1 MEM_stage_inst_dmem_U10473 ( .A1(MEM_stage_inst_dmem_ram_965), .A2(MEM_stage_inst_dmem_n13906), .ZN(MEM_stage_inst_dmem_n13894) );
NAND2_X1 MEM_stage_inst_dmem_U10472 ( .A1(MEM_stage_inst_dmem_n13891), .A2(MEM_stage_inst_dmem_n13890), .ZN(MEM_stage_inst_dmem_n12289) );
NAND2_X1 MEM_stage_inst_dmem_U10471 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n13907), .ZN(MEM_stage_inst_dmem_n13890) );
NAND2_X1 MEM_stage_inst_dmem_U10470 ( .A1(MEM_stage_inst_dmem_ram_966), .A2(MEM_stage_inst_dmem_n13906), .ZN(MEM_stage_inst_dmem_n13891) );
NAND2_X1 MEM_stage_inst_dmem_U10469 ( .A1(MEM_stage_inst_dmem_n13888), .A2(MEM_stage_inst_dmem_n13887), .ZN(MEM_stage_inst_dmem_n12290) );
NAND2_X1 MEM_stage_inst_dmem_U10468 ( .A1(MEM_stage_inst_dmem_n13886), .A2(MEM_stage_inst_dmem_n13907), .ZN(MEM_stage_inst_dmem_n13887) );
NAND2_X1 MEM_stage_inst_dmem_U10467 ( .A1(MEM_stage_inst_dmem_ram_967), .A2(MEM_stage_inst_dmem_n13906), .ZN(MEM_stage_inst_dmem_n13888) );
NAND2_X1 MEM_stage_inst_dmem_U10466 ( .A1(MEM_stage_inst_dmem_n13885), .A2(MEM_stage_inst_dmem_n13884), .ZN(MEM_stage_inst_dmem_n12291) );
NAND2_X1 MEM_stage_inst_dmem_U10465 ( .A1(MEM_stage_inst_dmem_n13883), .A2(MEM_stage_inst_dmem_n13907), .ZN(MEM_stage_inst_dmem_n13884) );
NAND2_X1 MEM_stage_inst_dmem_U10464 ( .A1(MEM_stage_inst_dmem_ram_968), .A2(MEM_stage_inst_dmem_n13906), .ZN(MEM_stage_inst_dmem_n13885) );
NAND2_X1 MEM_stage_inst_dmem_U10463 ( .A1(MEM_stage_inst_dmem_n13882), .A2(MEM_stage_inst_dmem_n13881), .ZN(MEM_stage_inst_dmem_n12292) );
NAND2_X1 MEM_stage_inst_dmem_U10462 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n13907), .ZN(MEM_stage_inst_dmem_n13881) );
NAND2_X1 MEM_stage_inst_dmem_U10461 ( .A1(MEM_stage_inst_dmem_ram_969), .A2(MEM_stage_inst_dmem_n13906), .ZN(MEM_stage_inst_dmem_n13882) );
NAND2_X1 MEM_stage_inst_dmem_U10460 ( .A1(MEM_stage_inst_dmem_n13879), .A2(MEM_stage_inst_dmem_n13878), .ZN(MEM_stage_inst_dmem_n12293) );
NAND2_X1 MEM_stage_inst_dmem_U10459 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n13907), .ZN(MEM_stage_inst_dmem_n13878) );
NAND2_X1 MEM_stage_inst_dmem_U10458 ( .A1(MEM_stage_inst_dmem_ram_970), .A2(MEM_stage_inst_dmem_n13906), .ZN(MEM_stage_inst_dmem_n13879) );
NAND2_X1 MEM_stage_inst_dmem_U10457 ( .A1(MEM_stage_inst_dmem_n13876), .A2(MEM_stage_inst_dmem_n13875), .ZN(MEM_stage_inst_dmem_n12294) );
NAND2_X1 MEM_stage_inst_dmem_U10456 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n13907), .ZN(MEM_stage_inst_dmem_n13875) );
NAND2_X1 MEM_stage_inst_dmem_U10455 ( .A1(MEM_stage_inst_dmem_ram_971), .A2(MEM_stage_inst_dmem_n13906), .ZN(MEM_stage_inst_dmem_n13876) );
NAND2_X1 MEM_stage_inst_dmem_U10454 ( .A1(MEM_stage_inst_dmem_n13873), .A2(MEM_stage_inst_dmem_n13872), .ZN(MEM_stage_inst_dmem_n12295) );
NAND2_X1 MEM_stage_inst_dmem_U10453 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n13907), .ZN(MEM_stage_inst_dmem_n13872) );
NAND2_X1 MEM_stage_inst_dmem_U10452 ( .A1(MEM_stage_inst_dmem_ram_972), .A2(MEM_stage_inst_dmem_n13906), .ZN(MEM_stage_inst_dmem_n13873) );
NAND2_X1 MEM_stage_inst_dmem_U10451 ( .A1(MEM_stage_inst_dmem_n13870), .A2(MEM_stage_inst_dmem_n13869), .ZN(MEM_stage_inst_dmem_n12296) );
NAND2_X1 MEM_stage_inst_dmem_U10450 ( .A1(MEM_stage_inst_dmem_n15116), .A2(MEM_stage_inst_dmem_n13907), .ZN(MEM_stage_inst_dmem_n13869) );
NAND2_X1 MEM_stage_inst_dmem_U10449 ( .A1(MEM_stage_inst_dmem_ram_973), .A2(MEM_stage_inst_dmem_n13906), .ZN(MEM_stage_inst_dmem_n13870) );
NAND2_X1 MEM_stage_inst_dmem_U10448 ( .A1(MEM_stage_inst_dmem_n13868), .A2(MEM_stage_inst_dmem_n13867), .ZN(MEM_stage_inst_dmem_n12297) );
NAND2_X1 MEM_stage_inst_dmem_U10447 ( .A1(MEM_stage_inst_dmem_n15113), .A2(MEM_stage_inst_dmem_n13907), .ZN(MEM_stage_inst_dmem_n13867) );
NAND2_X1 MEM_stage_inst_dmem_U10446 ( .A1(MEM_stage_inst_dmem_ram_974), .A2(MEM_stage_inst_dmem_n13906), .ZN(MEM_stage_inst_dmem_n13868) );
NAND2_X1 MEM_stage_inst_dmem_U10445 ( .A1(MEM_stage_inst_dmem_n13866), .A2(MEM_stage_inst_dmem_n13865), .ZN(MEM_stage_inst_dmem_n12298) );
NAND2_X1 MEM_stage_inst_dmem_U10444 ( .A1(MEM_stage_inst_dmem_n21320), .A2(MEM_stage_inst_dmem_n13907), .ZN(MEM_stage_inst_dmem_n13865) );
INV_X1 MEM_stage_inst_dmem_U10443 ( .A(MEM_stage_inst_dmem_n13906), .ZN(MEM_stage_inst_dmem_n13907) );
NAND2_X1 MEM_stage_inst_dmem_U10442 ( .A1(MEM_stage_inst_dmem_ram_975), .A2(MEM_stage_inst_dmem_n13906), .ZN(MEM_stage_inst_dmem_n13866) );
NAND2_X1 MEM_stage_inst_dmem_U10441 ( .A1(MEM_stage_inst_dmem_n21039), .A2(MEM_stage_inst_dmem_n14284), .ZN(MEM_stage_inst_dmem_n13906) );
NAND2_X1 MEM_stage_inst_dmem_U10440 ( .A1(MEM_stage_inst_dmem_n13864), .A2(MEM_stage_inst_dmem_n13863), .ZN(MEM_stage_inst_dmem_n12299) );
NAND2_X1 MEM_stage_inst_dmem_U10439 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n13862), .ZN(MEM_stage_inst_dmem_n13863) );
NAND2_X1 MEM_stage_inst_dmem_U10438 ( .A1(MEM_stage_inst_dmem_ram_976), .A2(MEM_stage_inst_dmem_n13861), .ZN(MEM_stage_inst_dmem_n13864) );
NAND2_X1 MEM_stage_inst_dmem_U10437 ( .A1(MEM_stage_inst_dmem_n13860), .A2(MEM_stage_inst_dmem_n13859), .ZN(MEM_stage_inst_dmem_n12300) );
NAND2_X1 MEM_stage_inst_dmem_U10436 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n13862), .ZN(MEM_stage_inst_dmem_n13859) );
NAND2_X1 MEM_stage_inst_dmem_U10435 ( .A1(MEM_stage_inst_dmem_ram_977), .A2(MEM_stage_inst_dmem_n13861), .ZN(MEM_stage_inst_dmem_n13860) );
NAND2_X1 MEM_stage_inst_dmem_U10434 ( .A1(MEM_stage_inst_dmem_n13858), .A2(MEM_stage_inst_dmem_n13857), .ZN(MEM_stage_inst_dmem_n12301) );
NAND2_X1 MEM_stage_inst_dmem_U10433 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n13862), .ZN(MEM_stage_inst_dmem_n13857) );
NAND2_X1 MEM_stage_inst_dmem_U10432 ( .A1(MEM_stage_inst_dmem_ram_978), .A2(MEM_stage_inst_dmem_n13861), .ZN(MEM_stage_inst_dmem_n13858) );
NAND2_X1 MEM_stage_inst_dmem_U10431 ( .A1(MEM_stage_inst_dmem_n13856), .A2(MEM_stage_inst_dmem_n13855), .ZN(MEM_stage_inst_dmem_n12302) );
NAND2_X1 MEM_stage_inst_dmem_U10430 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n13862), .ZN(MEM_stage_inst_dmem_n13855) );
NAND2_X1 MEM_stage_inst_dmem_U10429 ( .A1(MEM_stage_inst_dmem_ram_979), .A2(MEM_stage_inst_dmem_n13861), .ZN(MEM_stage_inst_dmem_n13856) );
NAND2_X1 MEM_stage_inst_dmem_U10428 ( .A1(MEM_stage_inst_dmem_n13854), .A2(MEM_stage_inst_dmem_n13853), .ZN(MEM_stage_inst_dmem_n12303) );
NAND2_X1 MEM_stage_inst_dmem_U10427 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n13862), .ZN(MEM_stage_inst_dmem_n13853) );
NAND2_X1 MEM_stage_inst_dmem_U10426 ( .A1(MEM_stage_inst_dmem_ram_980), .A2(MEM_stage_inst_dmem_n13861), .ZN(MEM_stage_inst_dmem_n13854) );
NAND2_X1 MEM_stage_inst_dmem_U10425 ( .A1(MEM_stage_inst_dmem_n13852), .A2(MEM_stage_inst_dmem_n13851), .ZN(MEM_stage_inst_dmem_n12304) );
NAND2_X1 MEM_stage_inst_dmem_U10424 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n13862), .ZN(MEM_stage_inst_dmem_n13851) );
NAND2_X1 MEM_stage_inst_dmem_U10423 ( .A1(MEM_stage_inst_dmem_ram_981), .A2(MEM_stage_inst_dmem_n13861), .ZN(MEM_stage_inst_dmem_n13852) );
NAND2_X1 MEM_stage_inst_dmem_U10422 ( .A1(MEM_stage_inst_dmem_n13850), .A2(MEM_stage_inst_dmem_n13849), .ZN(MEM_stage_inst_dmem_n12305) );
NAND2_X1 MEM_stage_inst_dmem_U10421 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n13862), .ZN(MEM_stage_inst_dmem_n13849) );
NAND2_X1 MEM_stage_inst_dmem_U10420 ( .A1(MEM_stage_inst_dmem_ram_982), .A2(MEM_stage_inst_dmem_n13861), .ZN(MEM_stage_inst_dmem_n13850) );
NAND2_X1 MEM_stage_inst_dmem_U10419 ( .A1(MEM_stage_inst_dmem_n13848), .A2(MEM_stage_inst_dmem_n13847), .ZN(MEM_stage_inst_dmem_n12306) );
NAND2_X1 MEM_stage_inst_dmem_U10418 ( .A1(MEM_stage_inst_dmem_n13886), .A2(MEM_stage_inst_dmem_n13862), .ZN(MEM_stage_inst_dmem_n13847) );
NAND2_X1 MEM_stage_inst_dmem_U10417 ( .A1(MEM_stage_inst_dmem_ram_983), .A2(MEM_stage_inst_dmem_n13861), .ZN(MEM_stage_inst_dmem_n13848) );
NAND2_X1 MEM_stage_inst_dmem_U10416 ( .A1(MEM_stage_inst_dmem_n13846), .A2(MEM_stage_inst_dmem_n13845), .ZN(MEM_stage_inst_dmem_n12307) );
NAND2_X1 MEM_stage_inst_dmem_U10415 ( .A1(MEM_stage_inst_dmem_n13883), .A2(MEM_stage_inst_dmem_n13862), .ZN(MEM_stage_inst_dmem_n13845) );
NAND2_X1 MEM_stage_inst_dmem_U10414 ( .A1(MEM_stage_inst_dmem_ram_984), .A2(MEM_stage_inst_dmem_n13861), .ZN(MEM_stage_inst_dmem_n13846) );
NAND2_X1 MEM_stage_inst_dmem_U10413 ( .A1(MEM_stage_inst_dmem_n13844), .A2(MEM_stage_inst_dmem_n13843), .ZN(MEM_stage_inst_dmem_n12308) );
NAND2_X1 MEM_stage_inst_dmem_U10412 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n13862), .ZN(MEM_stage_inst_dmem_n13843) );
NAND2_X1 MEM_stage_inst_dmem_U10411 ( .A1(MEM_stage_inst_dmem_ram_985), .A2(MEM_stage_inst_dmem_n13861), .ZN(MEM_stage_inst_dmem_n13844) );
NAND2_X1 MEM_stage_inst_dmem_U10410 ( .A1(MEM_stage_inst_dmem_n13842), .A2(MEM_stage_inst_dmem_n13841), .ZN(MEM_stage_inst_dmem_n12309) );
NAND2_X1 MEM_stage_inst_dmem_U10409 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n13862), .ZN(MEM_stage_inst_dmem_n13841) );
NAND2_X1 MEM_stage_inst_dmem_U10408 ( .A1(MEM_stage_inst_dmem_ram_986), .A2(MEM_stage_inst_dmem_n13861), .ZN(MEM_stage_inst_dmem_n13842) );
NAND2_X1 MEM_stage_inst_dmem_U10407 ( .A1(MEM_stage_inst_dmem_n13840), .A2(MEM_stage_inst_dmem_n13839), .ZN(MEM_stage_inst_dmem_n12310) );
NAND2_X1 MEM_stage_inst_dmem_U10406 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n13862), .ZN(MEM_stage_inst_dmem_n13839) );
NAND2_X1 MEM_stage_inst_dmem_U10405 ( .A1(MEM_stage_inst_dmem_ram_987), .A2(MEM_stage_inst_dmem_n13861), .ZN(MEM_stage_inst_dmem_n13840) );
NAND2_X1 MEM_stage_inst_dmem_U10404 ( .A1(MEM_stage_inst_dmem_n13838), .A2(MEM_stage_inst_dmem_n13837), .ZN(MEM_stage_inst_dmem_n12311) );
NAND2_X1 MEM_stage_inst_dmem_U10403 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n13862), .ZN(MEM_stage_inst_dmem_n13837) );
NAND2_X1 MEM_stage_inst_dmem_U10402 ( .A1(MEM_stage_inst_dmem_ram_988), .A2(MEM_stage_inst_dmem_n13861), .ZN(MEM_stage_inst_dmem_n13838) );
NAND2_X1 MEM_stage_inst_dmem_U10401 ( .A1(MEM_stage_inst_dmem_n13836), .A2(MEM_stage_inst_dmem_n13835), .ZN(MEM_stage_inst_dmem_n12312) );
NAND2_X1 MEM_stage_inst_dmem_U10400 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n13862), .ZN(MEM_stage_inst_dmem_n13835) );
NAND2_X1 MEM_stage_inst_dmem_U10399 ( .A1(MEM_stage_inst_dmem_ram_989), .A2(MEM_stage_inst_dmem_n13861), .ZN(MEM_stage_inst_dmem_n13836) );
NAND2_X1 MEM_stage_inst_dmem_U10398 ( .A1(MEM_stage_inst_dmem_n13834), .A2(MEM_stage_inst_dmem_n13833), .ZN(MEM_stage_inst_dmem_n12313) );
NAND2_X1 MEM_stage_inst_dmem_U10397 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n13862), .ZN(MEM_stage_inst_dmem_n13833) );
NAND2_X1 MEM_stage_inst_dmem_U10396 ( .A1(MEM_stage_inst_dmem_ram_990), .A2(MEM_stage_inst_dmem_n13861), .ZN(MEM_stage_inst_dmem_n13834) );
NAND2_X1 MEM_stage_inst_dmem_U10395 ( .A1(MEM_stage_inst_dmem_n13832), .A2(MEM_stage_inst_dmem_n13831), .ZN(MEM_stage_inst_dmem_n12314) );
NAND2_X1 MEM_stage_inst_dmem_U10394 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n13862), .ZN(MEM_stage_inst_dmem_n13831) );
INV_X1 MEM_stage_inst_dmem_U10393 ( .A(MEM_stage_inst_dmem_n13861), .ZN(MEM_stage_inst_dmem_n13862) );
NAND2_X1 MEM_stage_inst_dmem_U10392 ( .A1(MEM_stage_inst_dmem_ram_991), .A2(MEM_stage_inst_dmem_n13861), .ZN(MEM_stage_inst_dmem_n13832) );
NAND2_X1 MEM_stage_inst_dmem_U10391 ( .A1(MEM_stage_inst_dmem_n21004), .A2(MEM_stage_inst_dmem_n14284), .ZN(MEM_stage_inst_dmem_n13861) );
NAND2_X1 MEM_stage_inst_dmem_U10390 ( .A1(MEM_stage_inst_dmem_n13830), .A2(MEM_stage_inst_dmem_n13829), .ZN(MEM_stage_inst_dmem_n12315) );
NAND2_X1 MEM_stage_inst_dmem_U10389 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n13828), .ZN(MEM_stage_inst_dmem_n13829) );
NAND2_X1 MEM_stage_inst_dmem_U10388 ( .A1(MEM_stage_inst_dmem_ram_992), .A2(MEM_stage_inst_dmem_n13827), .ZN(MEM_stage_inst_dmem_n13830) );
NAND2_X1 MEM_stage_inst_dmem_U10387 ( .A1(MEM_stage_inst_dmem_n13826), .A2(MEM_stage_inst_dmem_n13825), .ZN(MEM_stage_inst_dmem_n12316) );
NAND2_X1 MEM_stage_inst_dmem_U10386 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n13828), .ZN(MEM_stage_inst_dmem_n13825) );
NAND2_X1 MEM_stage_inst_dmem_U10385 ( .A1(MEM_stage_inst_dmem_ram_993), .A2(MEM_stage_inst_dmem_n13827), .ZN(MEM_stage_inst_dmem_n13826) );
NAND2_X1 MEM_stage_inst_dmem_U10384 ( .A1(MEM_stage_inst_dmem_n13824), .A2(MEM_stage_inst_dmem_n13823), .ZN(MEM_stage_inst_dmem_n12317) );
NAND2_X1 MEM_stage_inst_dmem_U10383 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n13828), .ZN(MEM_stage_inst_dmem_n13823) );
NAND2_X1 MEM_stage_inst_dmem_U10382 ( .A1(MEM_stage_inst_dmem_ram_994), .A2(MEM_stage_inst_dmem_n13827), .ZN(MEM_stage_inst_dmem_n13824) );
NAND2_X1 MEM_stage_inst_dmem_U10381 ( .A1(MEM_stage_inst_dmem_n13822), .A2(MEM_stage_inst_dmem_n13821), .ZN(MEM_stage_inst_dmem_n12318) );
NAND2_X1 MEM_stage_inst_dmem_U10380 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n13828), .ZN(MEM_stage_inst_dmem_n13821) );
NAND2_X1 MEM_stage_inst_dmem_U10379 ( .A1(MEM_stage_inst_dmem_ram_995), .A2(MEM_stage_inst_dmem_n13827), .ZN(MEM_stage_inst_dmem_n13822) );
NAND2_X1 MEM_stage_inst_dmem_U10378 ( .A1(MEM_stage_inst_dmem_n13820), .A2(MEM_stage_inst_dmem_n13819), .ZN(MEM_stage_inst_dmem_n12319) );
NAND2_X1 MEM_stage_inst_dmem_U10377 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n13828), .ZN(MEM_stage_inst_dmem_n13819) );
NAND2_X1 MEM_stage_inst_dmem_U10376 ( .A1(MEM_stage_inst_dmem_ram_996), .A2(MEM_stage_inst_dmem_n13827), .ZN(MEM_stage_inst_dmem_n13820) );
NAND2_X1 MEM_stage_inst_dmem_U10375 ( .A1(MEM_stage_inst_dmem_n13818), .A2(MEM_stage_inst_dmem_n13817), .ZN(MEM_stage_inst_dmem_n12320) );
NAND2_X1 MEM_stage_inst_dmem_U10374 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n13828), .ZN(MEM_stage_inst_dmem_n13817) );
NAND2_X1 MEM_stage_inst_dmem_U10373 ( .A1(MEM_stage_inst_dmem_ram_997), .A2(MEM_stage_inst_dmem_n13827), .ZN(MEM_stage_inst_dmem_n13818) );
NAND2_X1 MEM_stage_inst_dmem_U10372 ( .A1(MEM_stage_inst_dmem_n13816), .A2(MEM_stage_inst_dmem_n13815), .ZN(MEM_stage_inst_dmem_n12321) );
NAND2_X1 MEM_stage_inst_dmem_U10371 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n13828), .ZN(MEM_stage_inst_dmem_n13815) );
NAND2_X1 MEM_stage_inst_dmem_U10370 ( .A1(MEM_stage_inst_dmem_ram_998), .A2(MEM_stage_inst_dmem_n13827), .ZN(MEM_stage_inst_dmem_n13816) );
NAND2_X1 MEM_stage_inst_dmem_U10369 ( .A1(MEM_stage_inst_dmem_n13814), .A2(MEM_stage_inst_dmem_n13813), .ZN(MEM_stage_inst_dmem_n12322) );
NAND2_X1 MEM_stage_inst_dmem_U10368 ( .A1(MEM_stage_inst_dmem_n13886), .A2(MEM_stage_inst_dmem_n13828), .ZN(MEM_stage_inst_dmem_n13813) );
NAND2_X1 MEM_stage_inst_dmem_U10367 ( .A1(MEM_stage_inst_dmem_ram_999), .A2(MEM_stage_inst_dmem_n13827), .ZN(MEM_stage_inst_dmem_n13814) );
NAND2_X1 MEM_stage_inst_dmem_U10366 ( .A1(MEM_stage_inst_dmem_n13812), .A2(MEM_stage_inst_dmem_n13811), .ZN(MEM_stage_inst_dmem_n12323) );
NAND2_X1 MEM_stage_inst_dmem_U10365 ( .A1(MEM_stage_inst_dmem_n13883), .A2(MEM_stage_inst_dmem_n13828), .ZN(MEM_stage_inst_dmem_n13811) );
NAND2_X1 MEM_stage_inst_dmem_U10364 ( .A1(MEM_stage_inst_dmem_ram_1000), .A2(MEM_stage_inst_dmem_n13827), .ZN(MEM_stage_inst_dmem_n13812) );
NAND2_X1 MEM_stage_inst_dmem_U10363 ( .A1(MEM_stage_inst_dmem_n13810), .A2(MEM_stage_inst_dmem_n13809), .ZN(MEM_stage_inst_dmem_n12324) );
NAND2_X1 MEM_stage_inst_dmem_U10362 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n13828), .ZN(MEM_stage_inst_dmem_n13809) );
NAND2_X1 MEM_stage_inst_dmem_U10361 ( .A1(MEM_stage_inst_dmem_ram_1001), .A2(MEM_stage_inst_dmem_n13827), .ZN(MEM_stage_inst_dmem_n13810) );
NAND2_X1 MEM_stage_inst_dmem_U10360 ( .A1(MEM_stage_inst_dmem_n13808), .A2(MEM_stage_inst_dmem_n13807), .ZN(MEM_stage_inst_dmem_n12325) );
NAND2_X1 MEM_stage_inst_dmem_U10359 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n13828), .ZN(MEM_stage_inst_dmem_n13807) );
NAND2_X1 MEM_stage_inst_dmem_U10358 ( .A1(MEM_stage_inst_dmem_ram_1002), .A2(MEM_stage_inst_dmem_n13827), .ZN(MEM_stage_inst_dmem_n13808) );
NAND2_X1 MEM_stage_inst_dmem_U10357 ( .A1(MEM_stage_inst_dmem_n13806), .A2(MEM_stage_inst_dmem_n13805), .ZN(MEM_stage_inst_dmem_n12326) );
NAND2_X1 MEM_stage_inst_dmem_U10356 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n13828), .ZN(MEM_stage_inst_dmem_n13805) );
NAND2_X1 MEM_stage_inst_dmem_U10355 ( .A1(MEM_stage_inst_dmem_ram_1003), .A2(MEM_stage_inst_dmem_n13827), .ZN(MEM_stage_inst_dmem_n13806) );
NAND2_X1 MEM_stage_inst_dmem_U10354 ( .A1(MEM_stage_inst_dmem_n13804), .A2(MEM_stage_inst_dmem_n13803), .ZN(MEM_stage_inst_dmem_n12327) );
NAND2_X1 MEM_stage_inst_dmem_U10353 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n13828), .ZN(MEM_stage_inst_dmem_n13803) );
NAND2_X1 MEM_stage_inst_dmem_U10352 ( .A1(MEM_stage_inst_dmem_ram_1004), .A2(MEM_stage_inst_dmem_n13827), .ZN(MEM_stage_inst_dmem_n13804) );
NAND2_X1 MEM_stage_inst_dmem_U10351 ( .A1(MEM_stage_inst_dmem_n13802), .A2(MEM_stage_inst_dmem_n13801), .ZN(MEM_stage_inst_dmem_n12328) );
NAND2_X1 MEM_stage_inst_dmem_U10350 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n13828), .ZN(MEM_stage_inst_dmem_n13801) );
NAND2_X1 MEM_stage_inst_dmem_U10349 ( .A1(MEM_stage_inst_dmem_ram_1005), .A2(MEM_stage_inst_dmem_n13827), .ZN(MEM_stage_inst_dmem_n13802) );
NAND2_X1 MEM_stage_inst_dmem_U10348 ( .A1(MEM_stage_inst_dmem_n13800), .A2(MEM_stage_inst_dmem_n13799), .ZN(MEM_stage_inst_dmem_n12329) );
NAND2_X1 MEM_stage_inst_dmem_U10347 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n13828), .ZN(MEM_stage_inst_dmem_n13799) );
NAND2_X1 MEM_stage_inst_dmem_U10346 ( .A1(MEM_stage_inst_dmem_ram_1006), .A2(MEM_stage_inst_dmem_n13827), .ZN(MEM_stage_inst_dmem_n13800) );
NAND2_X1 MEM_stage_inst_dmem_U10345 ( .A1(MEM_stage_inst_dmem_n13798), .A2(MEM_stage_inst_dmem_n13797), .ZN(MEM_stage_inst_dmem_n12330) );
NAND2_X1 MEM_stage_inst_dmem_U10344 ( .A1(MEM_stage_inst_dmem_n14693), .A2(MEM_stage_inst_dmem_n13828), .ZN(MEM_stage_inst_dmem_n13797) );
INV_X1 MEM_stage_inst_dmem_U10343 ( .A(MEM_stage_inst_dmem_n13827), .ZN(MEM_stage_inst_dmem_n13828) );
NAND2_X1 MEM_stage_inst_dmem_U10342 ( .A1(MEM_stage_inst_dmem_ram_1007), .A2(MEM_stage_inst_dmem_n13827), .ZN(MEM_stage_inst_dmem_n13798) );
NAND2_X1 MEM_stage_inst_dmem_U10341 ( .A1(MEM_stage_inst_dmem_n20969), .A2(MEM_stage_inst_dmem_n14284), .ZN(MEM_stage_inst_dmem_n13827) );
NAND2_X1 MEM_stage_inst_dmem_U10340 ( .A1(MEM_stage_inst_dmem_n13796), .A2(MEM_stage_inst_dmem_n13795), .ZN(MEM_stage_inst_dmem_n12331) );
NAND2_X1 MEM_stage_inst_dmem_U10339 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n13794), .ZN(MEM_stage_inst_dmem_n13795) );
NAND2_X1 MEM_stage_inst_dmem_U10338 ( .A1(MEM_stage_inst_dmem_ram_1008), .A2(MEM_stage_inst_dmem_n13793), .ZN(MEM_stage_inst_dmem_n13796) );
NAND2_X1 MEM_stage_inst_dmem_U10337 ( .A1(MEM_stage_inst_dmem_n13792), .A2(MEM_stage_inst_dmem_n13791), .ZN(MEM_stage_inst_dmem_n12332) );
NAND2_X1 MEM_stage_inst_dmem_U10336 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n13794), .ZN(MEM_stage_inst_dmem_n13791) );
NAND2_X1 MEM_stage_inst_dmem_U10335 ( .A1(MEM_stage_inst_dmem_ram_1009), .A2(MEM_stage_inst_dmem_n13793), .ZN(MEM_stage_inst_dmem_n13792) );
NAND2_X1 MEM_stage_inst_dmem_U10334 ( .A1(MEM_stage_inst_dmem_n13790), .A2(MEM_stage_inst_dmem_n13789), .ZN(MEM_stage_inst_dmem_n12333) );
NAND2_X1 MEM_stage_inst_dmem_U10333 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n13794), .ZN(MEM_stage_inst_dmem_n13789) );
NAND2_X1 MEM_stage_inst_dmem_U10332 ( .A1(MEM_stage_inst_dmem_ram_1010), .A2(MEM_stage_inst_dmem_n13793), .ZN(MEM_stage_inst_dmem_n13790) );
NAND2_X1 MEM_stage_inst_dmem_U10331 ( .A1(MEM_stage_inst_dmem_n13788), .A2(MEM_stage_inst_dmem_n13787), .ZN(MEM_stage_inst_dmem_n12334) );
NAND2_X1 MEM_stage_inst_dmem_U10330 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n13794), .ZN(MEM_stage_inst_dmem_n13787) );
NAND2_X1 MEM_stage_inst_dmem_U10329 ( .A1(MEM_stage_inst_dmem_ram_1011), .A2(MEM_stage_inst_dmem_n13793), .ZN(MEM_stage_inst_dmem_n13788) );
NAND2_X1 MEM_stage_inst_dmem_U10328 ( .A1(MEM_stage_inst_dmem_n13786), .A2(MEM_stage_inst_dmem_n13785), .ZN(MEM_stage_inst_dmem_n12335) );
NAND2_X1 MEM_stage_inst_dmem_U10327 ( .A1(EX_pipeline_reg_out_9), .A2(MEM_stage_inst_dmem_n13794), .ZN(MEM_stage_inst_dmem_n13785) );
NAND2_X1 MEM_stage_inst_dmem_U10326 ( .A1(MEM_stage_inst_dmem_ram_1012), .A2(MEM_stage_inst_dmem_n13793), .ZN(MEM_stage_inst_dmem_n13786) );
NAND2_X1 MEM_stage_inst_dmem_U10325 ( .A1(MEM_stage_inst_dmem_n13784), .A2(MEM_stage_inst_dmem_n13783), .ZN(MEM_stage_inst_dmem_n12336) );
NAND2_X1 MEM_stage_inst_dmem_U10324 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n13794), .ZN(MEM_stage_inst_dmem_n13783) );
NAND2_X1 MEM_stage_inst_dmem_U10323 ( .A1(MEM_stage_inst_dmem_ram_1013), .A2(MEM_stage_inst_dmem_n13793), .ZN(MEM_stage_inst_dmem_n13784) );
NAND2_X1 MEM_stage_inst_dmem_U10322 ( .A1(MEM_stage_inst_dmem_n13782), .A2(MEM_stage_inst_dmem_n13781), .ZN(MEM_stage_inst_dmem_n12337) );
NAND2_X1 MEM_stage_inst_dmem_U10321 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n13794), .ZN(MEM_stage_inst_dmem_n13781) );
NAND2_X1 MEM_stage_inst_dmem_U10320 ( .A1(MEM_stage_inst_dmem_ram_1014), .A2(MEM_stage_inst_dmem_n13793), .ZN(MEM_stage_inst_dmem_n13782) );
NAND2_X1 MEM_stage_inst_dmem_U10319 ( .A1(MEM_stage_inst_dmem_n13780), .A2(MEM_stage_inst_dmem_n13779), .ZN(MEM_stage_inst_dmem_n12338) );
NAND2_X1 MEM_stage_inst_dmem_U10318 ( .A1(MEM_stage_inst_dmem_n13886), .A2(MEM_stage_inst_dmem_n13794), .ZN(MEM_stage_inst_dmem_n13779) );
NAND2_X1 MEM_stage_inst_dmem_U10317 ( .A1(MEM_stage_inst_dmem_ram_1015), .A2(MEM_stage_inst_dmem_n13793), .ZN(MEM_stage_inst_dmem_n13780) );
NAND2_X1 MEM_stage_inst_dmem_U10316 ( .A1(MEM_stage_inst_dmem_n13778), .A2(MEM_stage_inst_dmem_n13777), .ZN(MEM_stage_inst_dmem_n12339) );
NAND2_X1 MEM_stage_inst_dmem_U10315 ( .A1(MEM_stage_inst_dmem_n13883), .A2(MEM_stage_inst_dmem_n13794), .ZN(MEM_stage_inst_dmem_n13777) );
NAND2_X1 MEM_stage_inst_dmem_U10314 ( .A1(MEM_stage_inst_dmem_ram_1016), .A2(MEM_stage_inst_dmem_n13793), .ZN(MEM_stage_inst_dmem_n13778) );
NAND2_X1 MEM_stage_inst_dmem_U10313 ( .A1(MEM_stage_inst_dmem_n13776), .A2(MEM_stage_inst_dmem_n13775), .ZN(MEM_stage_inst_dmem_n12340) );
NAND2_X1 MEM_stage_inst_dmem_U10312 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n13794), .ZN(MEM_stage_inst_dmem_n13775) );
NAND2_X1 MEM_stage_inst_dmem_U10311 ( .A1(MEM_stage_inst_dmem_ram_1017), .A2(MEM_stage_inst_dmem_n13793), .ZN(MEM_stage_inst_dmem_n13776) );
NAND2_X1 MEM_stage_inst_dmem_U10310 ( .A1(MEM_stage_inst_dmem_n13774), .A2(MEM_stage_inst_dmem_n13773), .ZN(MEM_stage_inst_dmem_n12341) );
NAND2_X1 MEM_stage_inst_dmem_U10309 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n13794), .ZN(MEM_stage_inst_dmem_n13773) );
NAND2_X1 MEM_stage_inst_dmem_U10308 ( .A1(MEM_stage_inst_dmem_ram_1018), .A2(MEM_stage_inst_dmem_n13793), .ZN(MEM_stage_inst_dmem_n13774) );
NAND2_X1 MEM_stage_inst_dmem_U10307 ( .A1(MEM_stage_inst_dmem_n13772), .A2(MEM_stage_inst_dmem_n13771), .ZN(MEM_stage_inst_dmem_n12342) );
NAND2_X1 MEM_stage_inst_dmem_U10306 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n13794), .ZN(MEM_stage_inst_dmem_n13771) );
NAND2_X1 MEM_stage_inst_dmem_U10305 ( .A1(MEM_stage_inst_dmem_ram_1019), .A2(MEM_stage_inst_dmem_n13793), .ZN(MEM_stage_inst_dmem_n13772) );
NAND2_X1 MEM_stage_inst_dmem_U10304 ( .A1(MEM_stage_inst_dmem_n13770), .A2(MEM_stage_inst_dmem_n13769), .ZN(MEM_stage_inst_dmem_n12343) );
NAND2_X1 MEM_stage_inst_dmem_U10303 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n13794), .ZN(MEM_stage_inst_dmem_n13769) );
NAND2_X1 MEM_stage_inst_dmem_U10302 ( .A1(MEM_stage_inst_dmem_ram_1020), .A2(MEM_stage_inst_dmem_n13793), .ZN(MEM_stage_inst_dmem_n13770) );
NAND2_X1 MEM_stage_inst_dmem_U10301 ( .A1(MEM_stage_inst_dmem_n13768), .A2(MEM_stage_inst_dmem_n13767), .ZN(MEM_stage_inst_dmem_n12344) );
NAND2_X1 MEM_stage_inst_dmem_U10300 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n13794), .ZN(MEM_stage_inst_dmem_n13767) );
NAND2_X1 MEM_stage_inst_dmem_U10299 ( .A1(MEM_stage_inst_dmem_ram_1021), .A2(MEM_stage_inst_dmem_n13793), .ZN(MEM_stage_inst_dmem_n13768) );
NAND2_X1 MEM_stage_inst_dmem_U10298 ( .A1(MEM_stage_inst_dmem_n13766), .A2(MEM_stage_inst_dmem_n13765), .ZN(MEM_stage_inst_dmem_n12345) );
NAND2_X1 MEM_stage_inst_dmem_U10297 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n13794), .ZN(MEM_stage_inst_dmem_n13765) );
NAND2_X1 MEM_stage_inst_dmem_U10296 ( .A1(MEM_stage_inst_dmem_ram_1022), .A2(MEM_stage_inst_dmem_n13793), .ZN(MEM_stage_inst_dmem_n13766) );
NAND2_X1 MEM_stage_inst_dmem_U10295 ( .A1(MEM_stage_inst_dmem_n13764), .A2(MEM_stage_inst_dmem_n13763), .ZN(MEM_stage_inst_dmem_n12346) );
NAND2_X1 MEM_stage_inst_dmem_U10294 ( .A1(MEM_stage_inst_dmem_n16343), .A2(MEM_stage_inst_dmem_n13794), .ZN(MEM_stage_inst_dmem_n13763) );
INV_X1 MEM_stage_inst_dmem_U10293 ( .A(MEM_stage_inst_dmem_n13793), .ZN(MEM_stage_inst_dmem_n13794) );
NAND2_X1 MEM_stage_inst_dmem_U10292 ( .A1(MEM_stage_inst_dmem_ram_1023), .A2(MEM_stage_inst_dmem_n13793), .ZN(MEM_stage_inst_dmem_n13764) );
NAND2_X1 MEM_stage_inst_dmem_U10291 ( .A1(MEM_stage_inst_dmem_n20934), .A2(MEM_stage_inst_dmem_n14284), .ZN(MEM_stage_inst_dmem_n13793) );
NOR2_X2 MEM_stage_inst_dmem_U10290 ( .A1(MEM_stage_inst_dmem_n15968), .A2(MEM_stage_inst_dmem_n18718), .ZN(MEM_stage_inst_dmem_n14284) );
NAND2_X1 MEM_stage_inst_dmem_U10289 ( .A1(EX_pipeline_reg_out_28), .A2(MEM_stage_inst_dmem_n15966), .ZN(MEM_stage_inst_dmem_n18718) );
NAND2_X1 MEM_stage_inst_dmem_U10288 ( .A1(MEM_stage_inst_dmem_n13762), .A2(MEM_stage_inst_dmem_n13761), .ZN(MEM_stage_inst_dmem_n12347) );
NAND2_X1 MEM_stage_inst_dmem_U10287 ( .A1(MEM_stage_inst_dmem_n15145), .A2(MEM_stage_inst_dmem_n13760), .ZN(MEM_stage_inst_dmem_n13761) );
NAND2_X1 MEM_stage_inst_dmem_U10286 ( .A1(MEM_stage_inst_dmem_ram_0), .A2(MEM_stage_inst_dmem_n13759), .ZN(MEM_stage_inst_dmem_n13762) );
NAND2_X1 MEM_stage_inst_dmem_U10285 ( .A1(MEM_stage_inst_dmem_n13758), .A2(MEM_stage_inst_dmem_n13757), .ZN(MEM_stage_inst_dmem_n12348) );
NAND2_X1 MEM_stage_inst_dmem_U10284 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n13760), .ZN(MEM_stage_inst_dmem_n13757) );
NAND2_X1 MEM_stage_inst_dmem_U10283 ( .A1(MEM_stage_inst_dmem_ram_1), .A2(MEM_stage_inst_dmem_n13759), .ZN(MEM_stage_inst_dmem_n13758) );
NAND2_X1 MEM_stage_inst_dmem_U10282 ( .A1(MEM_stage_inst_dmem_n13756), .A2(MEM_stage_inst_dmem_n13755), .ZN(MEM_stage_inst_dmem_n12349) );
NAND2_X1 MEM_stage_inst_dmem_U10281 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n13760), .ZN(MEM_stage_inst_dmem_n13755) );
NAND2_X1 MEM_stage_inst_dmem_U10280 ( .A1(MEM_stage_inst_dmem_ram_2), .A2(MEM_stage_inst_dmem_n13759), .ZN(MEM_stage_inst_dmem_n13756) );
NAND2_X1 MEM_stage_inst_dmem_U10279 ( .A1(MEM_stage_inst_dmem_n13754), .A2(MEM_stage_inst_dmem_n13753), .ZN(MEM_stage_inst_dmem_n12350) );
NAND2_X1 MEM_stage_inst_dmem_U10278 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n13760), .ZN(MEM_stage_inst_dmem_n13753) );
NAND2_X1 MEM_stage_inst_dmem_U10277 ( .A1(MEM_stage_inst_dmem_ram_3), .A2(MEM_stage_inst_dmem_n13759), .ZN(MEM_stage_inst_dmem_n13754) );
NAND2_X1 MEM_stage_inst_dmem_U10276 ( .A1(MEM_stage_inst_dmem_n13752), .A2(MEM_stage_inst_dmem_n13751), .ZN(MEM_stage_inst_dmem_n12351) );
NAND2_X1 MEM_stage_inst_dmem_U10275 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n13760), .ZN(MEM_stage_inst_dmem_n13751) );
NAND2_X1 MEM_stage_inst_dmem_U10274 ( .A1(MEM_stage_inst_dmem_ram_4), .A2(MEM_stage_inst_dmem_n13759), .ZN(MEM_stage_inst_dmem_n13752) );
NAND2_X1 MEM_stage_inst_dmem_U10273 ( .A1(MEM_stage_inst_dmem_n13750), .A2(MEM_stage_inst_dmem_n13749), .ZN(MEM_stage_inst_dmem_n12352) );
NAND2_X1 MEM_stage_inst_dmem_U10272 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n13760), .ZN(MEM_stage_inst_dmem_n13749) );
NAND2_X1 MEM_stage_inst_dmem_U10271 ( .A1(MEM_stage_inst_dmem_ram_5), .A2(MEM_stage_inst_dmem_n13759), .ZN(MEM_stage_inst_dmem_n13750) );
NAND2_X1 MEM_stage_inst_dmem_U10270 ( .A1(MEM_stage_inst_dmem_n13748), .A2(MEM_stage_inst_dmem_n13747), .ZN(MEM_stage_inst_dmem_n12353) );
NAND2_X1 MEM_stage_inst_dmem_U10269 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n13760), .ZN(MEM_stage_inst_dmem_n13747) );
NAND2_X1 MEM_stage_inst_dmem_U10268 ( .A1(MEM_stage_inst_dmem_ram_6), .A2(MEM_stage_inst_dmem_n13759), .ZN(MEM_stage_inst_dmem_n13748) );
NAND2_X1 MEM_stage_inst_dmem_U10267 ( .A1(MEM_stage_inst_dmem_n13746), .A2(MEM_stage_inst_dmem_n13745), .ZN(MEM_stage_inst_dmem_n12354) );
NAND2_X1 MEM_stage_inst_dmem_U10266 ( .A1(MEM_stage_inst_dmem_n13886), .A2(MEM_stage_inst_dmem_n13760), .ZN(MEM_stage_inst_dmem_n13745) );
NAND2_X1 MEM_stage_inst_dmem_U10265 ( .A1(MEM_stage_inst_dmem_ram_7), .A2(MEM_stage_inst_dmem_n13759), .ZN(MEM_stage_inst_dmem_n13746) );
NAND2_X1 MEM_stage_inst_dmem_U10264 ( .A1(MEM_stage_inst_dmem_n13744), .A2(MEM_stage_inst_dmem_n13743), .ZN(MEM_stage_inst_dmem_n12355) );
NAND2_X1 MEM_stage_inst_dmem_U10263 ( .A1(MEM_stage_inst_dmem_n13883), .A2(MEM_stage_inst_dmem_n13760), .ZN(MEM_stage_inst_dmem_n13743) );
NAND2_X1 MEM_stage_inst_dmem_U10262 ( .A1(MEM_stage_inst_dmem_ram_8), .A2(MEM_stage_inst_dmem_n13759), .ZN(MEM_stage_inst_dmem_n13744) );
NAND2_X1 MEM_stage_inst_dmem_U10261 ( .A1(MEM_stage_inst_dmem_n13742), .A2(MEM_stage_inst_dmem_n13741), .ZN(MEM_stage_inst_dmem_n12356) );
NAND2_X1 MEM_stage_inst_dmem_U10260 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n13760), .ZN(MEM_stage_inst_dmem_n13741) );
NAND2_X1 MEM_stage_inst_dmem_U10259 ( .A1(MEM_stage_inst_dmem_ram_9), .A2(MEM_stage_inst_dmem_n13759), .ZN(MEM_stage_inst_dmem_n13742) );
NAND2_X1 MEM_stage_inst_dmem_U10258 ( .A1(MEM_stage_inst_dmem_n13740), .A2(MEM_stage_inst_dmem_n13739), .ZN(MEM_stage_inst_dmem_n12357) );
NAND2_X1 MEM_stage_inst_dmem_U10257 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n13760), .ZN(MEM_stage_inst_dmem_n13739) );
NAND2_X1 MEM_stage_inst_dmem_U10256 ( .A1(MEM_stage_inst_dmem_ram_10), .A2(MEM_stage_inst_dmem_n13759), .ZN(MEM_stage_inst_dmem_n13740) );
NAND2_X1 MEM_stage_inst_dmem_U10255 ( .A1(MEM_stage_inst_dmem_n13738), .A2(MEM_stage_inst_dmem_n13737), .ZN(MEM_stage_inst_dmem_n12358) );
NAND2_X1 MEM_stage_inst_dmem_U10254 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n13760), .ZN(MEM_stage_inst_dmem_n13737) );
NAND2_X1 MEM_stage_inst_dmem_U10253 ( .A1(MEM_stage_inst_dmem_ram_11), .A2(MEM_stage_inst_dmem_n13759), .ZN(MEM_stage_inst_dmem_n13738) );
NAND2_X1 MEM_stage_inst_dmem_U10252 ( .A1(MEM_stage_inst_dmem_n13736), .A2(MEM_stage_inst_dmem_n13735), .ZN(MEM_stage_inst_dmem_n12359) );
NAND2_X1 MEM_stage_inst_dmem_U10251 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n13760), .ZN(MEM_stage_inst_dmem_n13735) );
NAND2_X1 MEM_stage_inst_dmem_U10250 ( .A1(MEM_stage_inst_dmem_ram_12), .A2(MEM_stage_inst_dmem_n13759), .ZN(MEM_stage_inst_dmem_n13736) );
NAND2_X1 MEM_stage_inst_dmem_U10249 ( .A1(MEM_stage_inst_dmem_n13734), .A2(MEM_stage_inst_dmem_n13733), .ZN(MEM_stage_inst_dmem_n12360) );
NAND2_X1 MEM_stage_inst_dmem_U10248 ( .A1(MEM_stage_inst_dmem_n15116), .A2(MEM_stage_inst_dmem_n13760), .ZN(MEM_stage_inst_dmem_n13733) );
NAND2_X1 MEM_stage_inst_dmem_U10247 ( .A1(MEM_stage_inst_dmem_ram_13), .A2(MEM_stage_inst_dmem_n13759), .ZN(MEM_stage_inst_dmem_n13734) );
NAND2_X1 MEM_stage_inst_dmem_U10246 ( .A1(MEM_stage_inst_dmem_n13732), .A2(MEM_stage_inst_dmem_n13731), .ZN(MEM_stage_inst_dmem_n12361) );
NAND2_X1 MEM_stage_inst_dmem_U10245 ( .A1(MEM_stage_inst_dmem_n15113), .A2(MEM_stage_inst_dmem_n13760), .ZN(MEM_stage_inst_dmem_n13731) );
NAND2_X1 MEM_stage_inst_dmem_U10244 ( .A1(MEM_stage_inst_dmem_ram_14), .A2(MEM_stage_inst_dmem_n13759), .ZN(MEM_stage_inst_dmem_n13732) );
NAND2_X1 MEM_stage_inst_dmem_U10243 ( .A1(MEM_stage_inst_dmem_n13730), .A2(MEM_stage_inst_dmem_n13729), .ZN(MEM_stage_inst_dmem_n12362) );
NAND2_X1 MEM_stage_inst_dmem_U10242 ( .A1(MEM_stage_inst_dmem_n14693), .A2(MEM_stage_inst_dmem_n13760), .ZN(MEM_stage_inst_dmem_n13729) );
INV_X1 MEM_stage_inst_dmem_U10241 ( .A(MEM_stage_inst_dmem_n13759), .ZN(MEM_stage_inst_dmem_n13760) );
NAND2_X1 MEM_stage_inst_dmem_U10240 ( .A1(MEM_stage_inst_dmem_ram_15), .A2(MEM_stage_inst_dmem_n13759), .ZN(MEM_stage_inst_dmem_n13730) );
NAND2_X1 MEM_stage_inst_dmem_U10239 ( .A1(MEM_stage_inst_dmem_n21465), .A2(MEM_stage_inst_dmem_n13728), .ZN(MEM_stage_inst_dmem_n13759) );
NAND2_X1 MEM_stage_inst_dmem_U10238 ( .A1(MEM_stage_inst_dmem_n13727), .A2(MEM_stage_inst_dmem_n13726), .ZN(MEM_stage_inst_dmem_n12363) );
NAND2_X1 MEM_stage_inst_dmem_U10237 ( .A1(MEM_stage_inst_dmem_n14732), .A2(MEM_stage_inst_dmem_n13725), .ZN(MEM_stage_inst_dmem_n13726) );
NAND2_X1 MEM_stage_inst_dmem_U10236 ( .A1(MEM_stage_inst_dmem_ram_16), .A2(MEM_stage_inst_dmem_n13724), .ZN(MEM_stage_inst_dmem_n13727) );
NAND2_X1 MEM_stage_inst_dmem_U10235 ( .A1(MEM_stage_inst_dmem_n13723), .A2(MEM_stage_inst_dmem_n13722), .ZN(MEM_stage_inst_dmem_n12364) );
NAND2_X1 MEM_stage_inst_dmem_U10234 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n13725), .ZN(MEM_stage_inst_dmem_n13722) );
NAND2_X1 MEM_stage_inst_dmem_U10233 ( .A1(MEM_stage_inst_dmem_ram_17), .A2(MEM_stage_inst_dmem_n13724), .ZN(MEM_stage_inst_dmem_n13723) );
NAND2_X1 MEM_stage_inst_dmem_U10232 ( .A1(MEM_stage_inst_dmem_n13721), .A2(MEM_stage_inst_dmem_n13720), .ZN(MEM_stage_inst_dmem_n12365) );
NAND2_X1 MEM_stage_inst_dmem_U10231 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n13725), .ZN(MEM_stage_inst_dmem_n13720) );
NAND2_X1 MEM_stage_inst_dmem_U10230 ( .A1(MEM_stage_inst_dmem_ram_18), .A2(MEM_stage_inst_dmem_n13724), .ZN(MEM_stage_inst_dmem_n13721) );
NAND2_X1 MEM_stage_inst_dmem_U10229 ( .A1(MEM_stage_inst_dmem_n13719), .A2(MEM_stage_inst_dmem_n13718), .ZN(MEM_stage_inst_dmem_n12366) );
NAND2_X1 MEM_stage_inst_dmem_U10228 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n13725), .ZN(MEM_stage_inst_dmem_n13718) );
NAND2_X1 MEM_stage_inst_dmem_U10227 ( .A1(MEM_stage_inst_dmem_ram_19), .A2(MEM_stage_inst_dmem_n13724), .ZN(MEM_stage_inst_dmem_n13719) );
NAND2_X1 MEM_stage_inst_dmem_U10226 ( .A1(MEM_stage_inst_dmem_n13717), .A2(MEM_stage_inst_dmem_n13716), .ZN(MEM_stage_inst_dmem_n12367) );
NAND2_X1 MEM_stage_inst_dmem_U10225 ( .A1(MEM_stage_inst_dmem_n16368), .A2(MEM_stage_inst_dmem_n13725), .ZN(MEM_stage_inst_dmem_n13716) );
NAND2_X1 MEM_stage_inst_dmem_U10224 ( .A1(MEM_stage_inst_dmem_ram_20), .A2(MEM_stage_inst_dmem_n13724), .ZN(MEM_stage_inst_dmem_n13717) );
NAND2_X1 MEM_stage_inst_dmem_U10223 ( .A1(MEM_stage_inst_dmem_n13715), .A2(MEM_stage_inst_dmem_n13714), .ZN(MEM_stage_inst_dmem_n12368) );
NAND2_X1 MEM_stage_inst_dmem_U10222 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n13725), .ZN(MEM_stage_inst_dmem_n13714) );
NAND2_X1 MEM_stage_inst_dmem_U10221 ( .A1(MEM_stage_inst_dmem_ram_21), .A2(MEM_stage_inst_dmem_n13724), .ZN(MEM_stage_inst_dmem_n13715) );
NAND2_X1 MEM_stage_inst_dmem_U10220 ( .A1(MEM_stage_inst_dmem_n13713), .A2(MEM_stage_inst_dmem_n13712), .ZN(MEM_stage_inst_dmem_n12369) );
NAND2_X1 MEM_stage_inst_dmem_U10219 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n13725), .ZN(MEM_stage_inst_dmem_n13712) );
NAND2_X1 MEM_stage_inst_dmem_U10218 ( .A1(MEM_stage_inst_dmem_ram_22), .A2(MEM_stage_inst_dmem_n13724), .ZN(MEM_stage_inst_dmem_n13713) );
NAND2_X1 MEM_stage_inst_dmem_U10217 ( .A1(MEM_stage_inst_dmem_n13711), .A2(MEM_stage_inst_dmem_n13710), .ZN(MEM_stage_inst_dmem_n12370) );
NAND2_X1 MEM_stage_inst_dmem_U10216 ( .A1(MEM_stage_inst_dmem_n13886), .A2(MEM_stage_inst_dmem_n13725), .ZN(MEM_stage_inst_dmem_n13710) );
NAND2_X1 MEM_stage_inst_dmem_U10215 ( .A1(MEM_stage_inst_dmem_ram_23), .A2(MEM_stage_inst_dmem_n13724), .ZN(MEM_stage_inst_dmem_n13711) );
NAND2_X1 MEM_stage_inst_dmem_U10214 ( .A1(MEM_stage_inst_dmem_n13709), .A2(MEM_stage_inst_dmem_n13708), .ZN(MEM_stage_inst_dmem_n12371) );
NAND2_X1 MEM_stage_inst_dmem_U10213 ( .A1(MEM_stage_inst_dmem_n13883), .A2(MEM_stage_inst_dmem_n13725), .ZN(MEM_stage_inst_dmem_n13708) );
NAND2_X1 MEM_stage_inst_dmem_U10212 ( .A1(MEM_stage_inst_dmem_ram_24), .A2(MEM_stage_inst_dmem_n13724), .ZN(MEM_stage_inst_dmem_n13709) );
NAND2_X1 MEM_stage_inst_dmem_U10211 ( .A1(MEM_stage_inst_dmem_n13707), .A2(MEM_stage_inst_dmem_n13706), .ZN(MEM_stage_inst_dmem_n12372) );
NAND2_X1 MEM_stage_inst_dmem_U10210 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n13725), .ZN(MEM_stage_inst_dmem_n13706) );
NAND2_X1 MEM_stage_inst_dmem_U10209 ( .A1(MEM_stage_inst_dmem_ram_25), .A2(MEM_stage_inst_dmem_n13724), .ZN(MEM_stage_inst_dmem_n13707) );
NAND2_X1 MEM_stage_inst_dmem_U10208 ( .A1(MEM_stage_inst_dmem_n13705), .A2(MEM_stage_inst_dmem_n13704), .ZN(MEM_stage_inst_dmem_n12373) );
NAND2_X1 MEM_stage_inst_dmem_U10207 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n13725), .ZN(MEM_stage_inst_dmem_n13704) );
NAND2_X1 MEM_stage_inst_dmem_U10206 ( .A1(MEM_stage_inst_dmem_ram_26), .A2(MEM_stage_inst_dmem_n13724), .ZN(MEM_stage_inst_dmem_n13705) );
NAND2_X1 MEM_stage_inst_dmem_U10205 ( .A1(MEM_stage_inst_dmem_n13703), .A2(MEM_stage_inst_dmem_n13702), .ZN(MEM_stage_inst_dmem_n12374) );
NAND2_X1 MEM_stage_inst_dmem_U10204 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n13725), .ZN(MEM_stage_inst_dmem_n13702) );
NAND2_X1 MEM_stage_inst_dmem_U10203 ( .A1(MEM_stage_inst_dmem_ram_27), .A2(MEM_stage_inst_dmem_n13724), .ZN(MEM_stage_inst_dmem_n13703) );
NAND2_X1 MEM_stage_inst_dmem_U10202 ( .A1(MEM_stage_inst_dmem_n13701), .A2(MEM_stage_inst_dmem_n13700), .ZN(MEM_stage_inst_dmem_n12375) );
NAND2_X1 MEM_stage_inst_dmem_U10201 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n13725), .ZN(MEM_stage_inst_dmem_n13700) );
NAND2_X1 MEM_stage_inst_dmem_U10200 ( .A1(MEM_stage_inst_dmem_ram_28), .A2(MEM_stage_inst_dmem_n13724), .ZN(MEM_stage_inst_dmem_n13701) );
NAND2_X1 MEM_stage_inst_dmem_U10199 ( .A1(MEM_stage_inst_dmem_n13699), .A2(MEM_stage_inst_dmem_n13698), .ZN(MEM_stage_inst_dmem_n12376) );
NAND2_X1 MEM_stage_inst_dmem_U10198 ( .A1(MEM_stage_inst_dmem_n116), .A2(MEM_stage_inst_dmem_n13725), .ZN(MEM_stage_inst_dmem_n13698) );
NAND2_X1 MEM_stage_inst_dmem_U10197 ( .A1(MEM_stage_inst_dmem_ram_29), .A2(MEM_stage_inst_dmem_n13724), .ZN(MEM_stage_inst_dmem_n13699) );
NAND2_X1 MEM_stage_inst_dmem_U10196 ( .A1(MEM_stage_inst_dmem_n13697), .A2(MEM_stage_inst_dmem_n13696), .ZN(MEM_stage_inst_dmem_n12377) );
NAND2_X1 MEM_stage_inst_dmem_U10195 ( .A1(MEM_stage_inst_dmem_n14696), .A2(MEM_stage_inst_dmem_n13725), .ZN(MEM_stage_inst_dmem_n13696) );
NAND2_X1 MEM_stage_inst_dmem_U10194 ( .A1(MEM_stage_inst_dmem_ram_30), .A2(MEM_stage_inst_dmem_n13724), .ZN(MEM_stage_inst_dmem_n13697) );
NAND2_X1 MEM_stage_inst_dmem_U10193 ( .A1(MEM_stage_inst_dmem_n13695), .A2(MEM_stage_inst_dmem_n13694), .ZN(MEM_stage_inst_dmem_n12378) );
NAND2_X1 MEM_stage_inst_dmem_U10192 ( .A1(MEM_stage_inst_dmem_n16343), .A2(MEM_stage_inst_dmem_n13725), .ZN(MEM_stage_inst_dmem_n13694) );
INV_X1 MEM_stage_inst_dmem_U10191 ( .A(MEM_stage_inst_dmem_n13724), .ZN(MEM_stage_inst_dmem_n13725) );
NAND2_X1 MEM_stage_inst_dmem_U10190 ( .A1(MEM_stage_inst_dmem_ram_31), .A2(MEM_stage_inst_dmem_n13724), .ZN(MEM_stage_inst_dmem_n13695) );
NAND2_X1 MEM_stage_inst_dmem_U10189 ( .A1(MEM_stage_inst_dmem_n21429), .A2(MEM_stage_inst_dmem_n13728), .ZN(MEM_stage_inst_dmem_n13724) );
NAND2_X1 MEM_stage_inst_dmem_U10188 ( .A1(MEM_stage_inst_dmem_n13693), .A2(MEM_stage_inst_dmem_n13692), .ZN(MEM_stage_inst_dmem_n12379) );
NAND2_X1 MEM_stage_inst_dmem_U10187 ( .A1(MEM_stage_inst_dmem_n19275), .A2(MEM_stage_inst_dmem_n13691), .ZN(MEM_stage_inst_dmem_n13692) );
NAND2_X1 MEM_stage_inst_dmem_U10186 ( .A1(MEM_stage_inst_dmem_ram_32), .A2(MEM_stage_inst_dmem_n13690), .ZN(MEM_stage_inst_dmem_n13693) );
NAND2_X1 MEM_stage_inst_dmem_U10185 ( .A1(MEM_stage_inst_dmem_n13689), .A2(MEM_stage_inst_dmem_n13688), .ZN(MEM_stage_inst_dmem_n12380) );
NAND2_X1 MEM_stage_inst_dmem_U10184 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n13691), .ZN(MEM_stage_inst_dmem_n13688) );
NAND2_X1 MEM_stage_inst_dmem_U10183 ( .A1(MEM_stage_inst_dmem_ram_33), .A2(MEM_stage_inst_dmem_n13690), .ZN(MEM_stage_inst_dmem_n13689) );
NAND2_X1 MEM_stage_inst_dmem_U10182 ( .A1(MEM_stage_inst_dmem_n13687), .A2(MEM_stage_inst_dmem_n13686), .ZN(MEM_stage_inst_dmem_n12381) );
NAND2_X1 MEM_stage_inst_dmem_U10181 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n13691), .ZN(MEM_stage_inst_dmem_n13686) );
NAND2_X1 MEM_stage_inst_dmem_U10180 ( .A1(MEM_stage_inst_dmem_ram_34), .A2(MEM_stage_inst_dmem_n13690), .ZN(MEM_stage_inst_dmem_n13687) );
NAND2_X1 MEM_stage_inst_dmem_U10179 ( .A1(MEM_stage_inst_dmem_n13685), .A2(MEM_stage_inst_dmem_n13684), .ZN(MEM_stage_inst_dmem_n12382) );
NAND2_X1 MEM_stage_inst_dmem_U10178 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n13691), .ZN(MEM_stage_inst_dmem_n13684) );
NAND2_X1 MEM_stage_inst_dmem_U10177 ( .A1(MEM_stage_inst_dmem_ram_35), .A2(MEM_stage_inst_dmem_n13690), .ZN(MEM_stage_inst_dmem_n13685) );
NAND2_X1 MEM_stage_inst_dmem_U10176 ( .A1(MEM_stage_inst_dmem_n13683), .A2(MEM_stage_inst_dmem_n13682), .ZN(MEM_stage_inst_dmem_n12383) );
NAND2_X1 MEM_stage_inst_dmem_U10175 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n13691), .ZN(MEM_stage_inst_dmem_n13682) );
NAND2_X1 MEM_stage_inst_dmem_U10174 ( .A1(MEM_stage_inst_dmem_ram_36), .A2(MEM_stage_inst_dmem_n13690), .ZN(MEM_stage_inst_dmem_n13683) );
NAND2_X1 MEM_stage_inst_dmem_U10173 ( .A1(MEM_stage_inst_dmem_n13681), .A2(MEM_stage_inst_dmem_n13680), .ZN(MEM_stage_inst_dmem_n12384) );
NAND2_X1 MEM_stage_inst_dmem_U10172 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n13691), .ZN(MEM_stage_inst_dmem_n13680) );
NAND2_X1 MEM_stage_inst_dmem_U10171 ( .A1(MEM_stage_inst_dmem_ram_37), .A2(MEM_stage_inst_dmem_n13690), .ZN(MEM_stage_inst_dmem_n13681) );
NAND2_X1 MEM_stage_inst_dmem_U10170 ( .A1(MEM_stage_inst_dmem_n13679), .A2(MEM_stage_inst_dmem_n13678), .ZN(MEM_stage_inst_dmem_n12385) );
NAND2_X1 MEM_stage_inst_dmem_U10169 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n13691), .ZN(MEM_stage_inst_dmem_n13678) );
NAND2_X1 MEM_stage_inst_dmem_U10168 ( .A1(MEM_stage_inst_dmem_ram_38), .A2(MEM_stage_inst_dmem_n13690), .ZN(MEM_stage_inst_dmem_n13679) );
NAND2_X1 MEM_stage_inst_dmem_U10167 ( .A1(MEM_stage_inst_dmem_n13677), .A2(MEM_stage_inst_dmem_n13676), .ZN(MEM_stage_inst_dmem_n12386) );
NAND2_X1 MEM_stage_inst_dmem_U10166 ( .A1(MEM_stage_inst_dmem_n13886), .A2(MEM_stage_inst_dmem_n13691), .ZN(MEM_stage_inst_dmem_n13676) );
NAND2_X1 MEM_stage_inst_dmem_U10165 ( .A1(MEM_stage_inst_dmem_ram_39), .A2(MEM_stage_inst_dmem_n13690), .ZN(MEM_stage_inst_dmem_n13677) );
NAND2_X1 MEM_stage_inst_dmem_U10164 ( .A1(MEM_stage_inst_dmem_n13675), .A2(MEM_stage_inst_dmem_n13674), .ZN(MEM_stage_inst_dmem_n12387) );
NAND2_X1 MEM_stage_inst_dmem_U10163 ( .A1(MEM_stage_inst_dmem_n13883), .A2(MEM_stage_inst_dmem_n13691), .ZN(MEM_stage_inst_dmem_n13674) );
NAND2_X1 MEM_stage_inst_dmem_U10162 ( .A1(MEM_stage_inst_dmem_ram_40), .A2(MEM_stage_inst_dmem_n13690), .ZN(MEM_stage_inst_dmem_n13675) );
NAND2_X1 MEM_stage_inst_dmem_U10161 ( .A1(MEM_stage_inst_dmem_n13673), .A2(MEM_stage_inst_dmem_n13672), .ZN(MEM_stage_inst_dmem_n12388) );
NAND2_X1 MEM_stage_inst_dmem_U10160 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n13691), .ZN(MEM_stage_inst_dmem_n13672) );
NAND2_X1 MEM_stage_inst_dmem_U10159 ( .A1(MEM_stage_inst_dmem_ram_41), .A2(MEM_stage_inst_dmem_n13690), .ZN(MEM_stage_inst_dmem_n13673) );
NAND2_X1 MEM_stage_inst_dmem_U10158 ( .A1(MEM_stage_inst_dmem_n13671), .A2(MEM_stage_inst_dmem_n13670), .ZN(MEM_stage_inst_dmem_n12389) );
NAND2_X1 MEM_stage_inst_dmem_U10157 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n13691), .ZN(MEM_stage_inst_dmem_n13670) );
NAND2_X1 MEM_stage_inst_dmem_U10156 ( .A1(MEM_stage_inst_dmem_ram_42), .A2(MEM_stage_inst_dmem_n13690), .ZN(MEM_stage_inst_dmem_n13671) );
NAND2_X1 MEM_stage_inst_dmem_U10155 ( .A1(MEM_stage_inst_dmem_n13669), .A2(MEM_stage_inst_dmem_n13668), .ZN(MEM_stage_inst_dmem_n12390) );
NAND2_X1 MEM_stage_inst_dmem_U10154 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n13691), .ZN(MEM_stage_inst_dmem_n13668) );
NAND2_X1 MEM_stage_inst_dmem_U10153 ( .A1(MEM_stage_inst_dmem_ram_43), .A2(MEM_stage_inst_dmem_n13690), .ZN(MEM_stage_inst_dmem_n13669) );
NAND2_X1 MEM_stage_inst_dmem_U10152 ( .A1(MEM_stage_inst_dmem_n13667), .A2(MEM_stage_inst_dmem_n13666), .ZN(MEM_stage_inst_dmem_n12391) );
NAND2_X1 MEM_stage_inst_dmem_U10151 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n13691), .ZN(MEM_stage_inst_dmem_n13666) );
NAND2_X1 MEM_stage_inst_dmem_U10150 ( .A1(MEM_stage_inst_dmem_ram_44), .A2(MEM_stage_inst_dmem_n13690), .ZN(MEM_stage_inst_dmem_n13667) );
NAND2_X1 MEM_stage_inst_dmem_U10149 ( .A1(MEM_stage_inst_dmem_n13665), .A2(MEM_stage_inst_dmem_n13664), .ZN(MEM_stage_inst_dmem_n12392) );
NAND2_X1 MEM_stage_inst_dmem_U10148 ( .A1(MEM_stage_inst_dmem_n19242), .A2(MEM_stage_inst_dmem_n13691), .ZN(MEM_stage_inst_dmem_n13664) );
NAND2_X1 MEM_stage_inst_dmem_U10147 ( .A1(MEM_stage_inst_dmem_ram_45), .A2(MEM_stage_inst_dmem_n13690), .ZN(MEM_stage_inst_dmem_n13665) );
NAND2_X1 MEM_stage_inst_dmem_U10146 ( .A1(MEM_stage_inst_dmem_n13663), .A2(MEM_stage_inst_dmem_n13662), .ZN(MEM_stage_inst_dmem_n12393) );
NAND2_X1 MEM_stage_inst_dmem_U10145 ( .A1(MEM_stage_inst_dmem_n115), .A2(MEM_stage_inst_dmem_n13691), .ZN(MEM_stage_inst_dmem_n13662) );
NAND2_X1 MEM_stage_inst_dmem_U10144 ( .A1(MEM_stage_inst_dmem_ram_46), .A2(MEM_stage_inst_dmem_n13690), .ZN(MEM_stage_inst_dmem_n13663) );
NAND2_X1 MEM_stage_inst_dmem_U10143 ( .A1(MEM_stage_inst_dmem_n13661), .A2(MEM_stage_inst_dmem_n13660), .ZN(MEM_stage_inst_dmem_n12394) );
NAND2_X1 MEM_stage_inst_dmem_U10142 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n13691), .ZN(MEM_stage_inst_dmem_n13660) );
NAND2_X1 MEM_stage_inst_dmem_U10141 ( .A1(MEM_stage_inst_dmem_ram_47), .A2(MEM_stage_inst_dmem_n13690), .ZN(MEM_stage_inst_dmem_n13661) );
NAND2_X1 MEM_stage_inst_dmem_U10140 ( .A1(MEM_stage_inst_dmem_n21394), .A2(MEM_stage_inst_dmem_n13728), .ZN(MEM_stage_inst_dmem_n13690) );
NAND2_X1 MEM_stage_inst_dmem_U10139 ( .A1(MEM_stage_inst_dmem_n13659), .A2(MEM_stage_inst_dmem_n13658), .ZN(MEM_stage_inst_dmem_n12395) );
NAND2_X1 MEM_stage_inst_dmem_U10138 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n13657), .ZN(MEM_stage_inst_dmem_n13658) );
NAND2_X1 MEM_stage_inst_dmem_U10137 ( .A1(MEM_stage_inst_dmem_ram_48), .A2(MEM_stage_inst_dmem_n13656), .ZN(MEM_stage_inst_dmem_n13659) );
NAND2_X1 MEM_stage_inst_dmem_U10136 ( .A1(MEM_stage_inst_dmem_n13655), .A2(MEM_stage_inst_dmem_n13654), .ZN(MEM_stage_inst_dmem_n12396) );
NAND2_X1 MEM_stage_inst_dmem_U10135 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n13657), .ZN(MEM_stage_inst_dmem_n13654) );
NAND2_X1 MEM_stage_inst_dmem_U10134 ( .A1(MEM_stage_inst_dmem_ram_49), .A2(MEM_stage_inst_dmem_n13656), .ZN(MEM_stage_inst_dmem_n13655) );
NAND2_X1 MEM_stage_inst_dmem_U10133 ( .A1(MEM_stage_inst_dmem_n13653), .A2(MEM_stage_inst_dmem_n13652), .ZN(MEM_stage_inst_dmem_n12397) );
NAND2_X1 MEM_stage_inst_dmem_U10132 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n13657), .ZN(MEM_stage_inst_dmem_n13652) );
NAND2_X1 MEM_stage_inst_dmem_U10131 ( .A1(MEM_stage_inst_dmem_ram_50), .A2(MEM_stage_inst_dmem_n13656), .ZN(MEM_stage_inst_dmem_n13653) );
NAND2_X1 MEM_stage_inst_dmem_U10130 ( .A1(MEM_stage_inst_dmem_n13651), .A2(MEM_stage_inst_dmem_n13650), .ZN(MEM_stage_inst_dmem_n12398) );
NAND2_X1 MEM_stage_inst_dmem_U10129 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n13657), .ZN(MEM_stage_inst_dmem_n13650) );
NAND2_X1 MEM_stage_inst_dmem_U10128 ( .A1(MEM_stage_inst_dmem_ram_51), .A2(MEM_stage_inst_dmem_n13656), .ZN(MEM_stage_inst_dmem_n13651) );
NAND2_X1 MEM_stage_inst_dmem_U10127 ( .A1(MEM_stage_inst_dmem_n13649), .A2(MEM_stage_inst_dmem_n13648), .ZN(MEM_stage_inst_dmem_n12399) );
NAND2_X1 MEM_stage_inst_dmem_U10126 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n13657), .ZN(MEM_stage_inst_dmem_n13648) );
NAND2_X1 MEM_stage_inst_dmem_U10125 ( .A1(MEM_stage_inst_dmem_ram_52), .A2(MEM_stage_inst_dmem_n13656), .ZN(MEM_stage_inst_dmem_n13649) );
NAND2_X1 MEM_stage_inst_dmem_U10124 ( .A1(MEM_stage_inst_dmem_n13647), .A2(MEM_stage_inst_dmem_n13646), .ZN(MEM_stage_inst_dmem_n12400) );
NAND2_X1 MEM_stage_inst_dmem_U10123 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n13657), .ZN(MEM_stage_inst_dmem_n13646) );
NAND2_X1 MEM_stage_inst_dmem_U10122 ( .A1(MEM_stage_inst_dmem_ram_53), .A2(MEM_stage_inst_dmem_n13656), .ZN(MEM_stage_inst_dmem_n13647) );
NAND2_X1 MEM_stage_inst_dmem_U10121 ( .A1(MEM_stage_inst_dmem_n13645), .A2(MEM_stage_inst_dmem_n13644), .ZN(MEM_stage_inst_dmem_n12401) );
NAND2_X1 MEM_stage_inst_dmem_U10120 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n13657), .ZN(MEM_stage_inst_dmem_n13644) );
NAND2_X1 MEM_stage_inst_dmem_U10119 ( .A1(MEM_stage_inst_dmem_ram_54), .A2(MEM_stage_inst_dmem_n13656), .ZN(MEM_stage_inst_dmem_n13645) );
NAND2_X1 MEM_stage_inst_dmem_U10118 ( .A1(MEM_stage_inst_dmem_n13643), .A2(MEM_stage_inst_dmem_n13642), .ZN(MEM_stage_inst_dmem_n12402) );
NAND2_X1 MEM_stage_inst_dmem_U10117 ( .A1(MEM_stage_inst_dmem_n13886), .A2(MEM_stage_inst_dmem_n13657), .ZN(MEM_stage_inst_dmem_n13642) );
NAND2_X1 MEM_stage_inst_dmem_U10116 ( .A1(MEM_stage_inst_dmem_ram_55), .A2(MEM_stage_inst_dmem_n13656), .ZN(MEM_stage_inst_dmem_n13643) );
NAND2_X1 MEM_stage_inst_dmem_U10115 ( .A1(MEM_stage_inst_dmem_n13641), .A2(MEM_stage_inst_dmem_n13640), .ZN(MEM_stage_inst_dmem_n12403) );
NAND2_X1 MEM_stage_inst_dmem_U10114 ( .A1(MEM_stage_inst_dmem_n13883), .A2(MEM_stage_inst_dmem_n13657), .ZN(MEM_stage_inst_dmem_n13640) );
NAND2_X1 MEM_stage_inst_dmem_U10113 ( .A1(MEM_stage_inst_dmem_ram_56), .A2(MEM_stage_inst_dmem_n13656), .ZN(MEM_stage_inst_dmem_n13641) );
NAND2_X1 MEM_stage_inst_dmem_U10112 ( .A1(MEM_stage_inst_dmem_n13639), .A2(MEM_stage_inst_dmem_n13638), .ZN(MEM_stage_inst_dmem_n12404) );
NAND2_X1 MEM_stage_inst_dmem_U10111 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n13657), .ZN(MEM_stage_inst_dmem_n13638) );
NAND2_X1 MEM_stage_inst_dmem_U10110 ( .A1(MEM_stage_inst_dmem_ram_57), .A2(MEM_stage_inst_dmem_n13656), .ZN(MEM_stage_inst_dmem_n13639) );
NAND2_X1 MEM_stage_inst_dmem_U10109 ( .A1(MEM_stage_inst_dmem_n13637), .A2(MEM_stage_inst_dmem_n13636), .ZN(MEM_stage_inst_dmem_n12405) );
NAND2_X1 MEM_stage_inst_dmem_U10108 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n13657), .ZN(MEM_stage_inst_dmem_n13636) );
NAND2_X1 MEM_stage_inst_dmem_U10107 ( .A1(MEM_stage_inst_dmem_ram_58), .A2(MEM_stage_inst_dmem_n13656), .ZN(MEM_stage_inst_dmem_n13637) );
NAND2_X1 MEM_stage_inst_dmem_U10106 ( .A1(MEM_stage_inst_dmem_n13635), .A2(MEM_stage_inst_dmem_n13634), .ZN(MEM_stage_inst_dmem_n12406) );
NAND2_X1 MEM_stage_inst_dmem_U10105 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n13657), .ZN(MEM_stage_inst_dmem_n13634) );
NAND2_X1 MEM_stage_inst_dmem_U10104 ( .A1(MEM_stage_inst_dmem_ram_59), .A2(MEM_stage_inst_dmem_n13656), .ZN(MEM_stage_inst_dmem_n13635) );
NAND2_X1 MEM_stage_inst_dmem_U10103 ( .A1(MEM_stage_inst_dmem_n13633), .A2(MEM_stage_inst_dmem_n13632), .ZN(MEM_stage_inst_dmem_n12407) );
NAND2_X1 MEM_stage_inst_dmem_U10102 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n13657), .ZN(MEM_stage_inst_dmem_n13632) );
NAND2_X1 MEM_stage_inst_dmem_U10101 ( .A1(MEM_stage_inst_dmem_ram_60), .A2(MEM_stage_inst_dmem_n13656), .ZN(MEM_stage_inst_dmem_n13633) );
NAND2_X1 MEM_stage_inst_dmem_U10100 ( .A1(MEM_stage_inst_dmem_n13631), .A2(MEM_stage_inst_dmem_n13630), .ZN(MEM_stage_inst_dmem_n12408) );
NAND2_X1 MEM_stage_inst_dmem_U10099 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n13657), .ZN(MEM_stage_inst_dmem_n13630) );
NAND2_X1 MEM_stage_inst_dmem_U10098 ( .A1(MEM_stage_inst_dmem_ram_61), .A2(MEM_stage_inst_dmem_n13656), .ZN(MEM_stage_inst_dmem_n13631) );
NAND2_X1 MEM_stage_inst_dmem_U10097 ( .A1(MEM_stage_inst_dmem_n13629), .A2(MEM_stage_inst_dmem_n13628), .ZN(MEM_stage_inst_dmem_n12409) );
NAND2_X1 MEM_stage_inst_dmem_U10096 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n13657), .ZN(MEM_stage_inst_dmem_n13628) );
NAND2_X1 MEM_stage_inst_dmem_U10095 ( .A1(MEM_stage_inst_dmem_ram_62), .A2(MEM_stage_inst_dmem_n13656), .ZN(MEM_stage_inst_dmem_n13629) );
NAND2_X1 MEM_stage_inst_dmem_U10094 ( .A1(MEM_stage_inst_dmem_n13627), .A2(MEM_stage_inst_dmem_n13626), .ZN(MEM_stage_inst_dmem_n12410) );
NAND2_X1 MEM_stage_inst_dmem_U10093 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n13657), .ZN(MEM_stage_inst_dmem_n13626) );
INV_X1 MEM_stage_inst_dmem_U10092 ( .A(MEM_stage_inst_dmem_n13656), .ZN(MEM_stage_inst_dmem_n13657) );
NAND2_X1 MEM_stage_inst_dmem_U10091 ( .A1(MEM_stage_inst_dmem_ram_63), .A2(MEM_stage_inst_dmem_n13656), .ZN(MEM_stage_inst_dmem_n13627) );
NAND2_X1 MEM_stage_inst_dmem_U10090 ( .A1(MEM_stage_inst_dmem_n21359), .A2(MEM_stage_inst_dmem_n13728), .ZN(MEM_stage_inst_dmem_n13656) );
NAND2_X1 MEM_stage_inst_dmem_U10089 ( .A1(MEM_stage_inst_dmem_n13625), .A2(MEM_stage_inst_dmem_n13624), .ZN(MEM_stage_inst_dmem_n12411) );
NAND2_X1 MEM_stage_inst_dmem_U10088 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n13623), .ZN(MEM_stage_inst_dmem_n13624) );
NAND2_X1 MEM_stage_inst_dmem_U10087 ( .A1(MEM_stage_inst_dmem_ram_64), .A2(MEM_stage_inst_dmem_n13622), .ZN(MEM_stage_inst_dmem_n13625) );
NAND2_X1 MEM_stage_inst_dmem_U10086 ( .A1(MEM_stage_inst_dmem_n13621), .A2(MEM_stage_inst_dmem_n13620), .ZN(MEM_stage_inst_dmem_n12412) );
NAND2_X1 MEM_stage_inst_dmem_U10085 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n13623), .ZN(MEM_stage_inst_dmem_n13620) );
NAND2_X1 MEM_stage_inst_dmem_U10084 ( .A1(MEM_stage_inst_dmem_ram_65), .A2(MEM_stage_inst_dmem_n13622), .ZN(MEM_stage_inst_dmem_n13621) );
NAND2_X1 MEM_stage_inst_dmem_U10083 ( .A1(MEM_stage_inst_dmem_n13619), .A2(MEM_stage_inst_dmem_n13618), .ZN(MEM_stage_inst_dmem_n12413) );
NAND2_X1 MEM_stage_inst_dmem_U10082 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n13623), .ZN(MEM_stage_inst_dmem_n13618) );
NAND2_X1 MEM_stage_inst_dmem_U10081 ( .A1(MEM_stage_inst_dmem_ram_66), .A2(MEM_stage_inst_dmem_n13622), .ZN(MEM_stage_inst_dmem_n13619) );
NAND2_X1 MEM_stage_inst_dmem_U10080 ( .A1(MEM_stage_inst_dmem_n13617), .A2(MEM_stage_inst_dmem_n13616), .ZN(MEM_stage_inst_dmem_n12414) );
NAND2_X1 MEM_stage_inst_dmem_U10079 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n13623), .ZN(MEM_stage_inst_dmem_n13616) );
NAND2_X1 MEM_stage_inst_dmem_U10078 ( .A1(MEM_stage_inst_dmem_ram_67), .A2(MEM_stage_inst_dmem_n13622), .ZN(MEM_stage_inst_dmem_n13617) );
NAND2_X1 MEM_stage_inst_dmem_U10077 ( .A1(MEM_stage_inst_dmem_n13615), .A2(MEM_stage_inst_dmem_n13614), .ZN(MEM_stage_inst_dmem_n12415) );
NAND2_X1 MEM_stage_inst_dmem_U10076 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n13623), .ZN(MEM_stage_inst_dmem_n13614) );
NAND2_X1 MEM_stage_inst_dmem_U10075 ( .A1(MEM_stage_inst_dmem_ram_68), .A2(MEM_stage_inst_dmem_n13622), .ZN(MEM_stage_inst_dmem_n13615) );
NAND2_X1 MEM_stage_inst_dmem_U10074 ( .A1(MEM_stage_inst_dmem_n13613), .A2(MEM_stage_inst_dmem_n13612), .ZN(MEM_stage_inst_dmem_n12416) );
NAND2_X1 MEM_stage_inst_dmem_U10073 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n13623), .ZN(MEM_stage_inst_dmem_n13612) );
NAND2_X1 MEM_stage_inst_dmem_U10072 ( .A1(MEM_stage_inst_dmem_ram_69), .A2(MEM_stage_inst_dmem_n13622), .ZN(MEM_stage_inst_dmem_n13613) );
NAND2_X1 MEM_stage_inst_dmem_U10071 ( .A1(MEM_stage_inst_dmem_n13611), .A2(MEM_stage_inst_dmem_n13610), .ZN(MEM_stage_inst_dmem_n12417) );
NAND2_X1 MEM_stage_inst_dmem_U10070 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n13623), .ZN(MEM_stage_inst_dmem_n13610) );
NAND2_X1 MEM_stage_inst_dmem_U10069 ( .A1(MEM_stage_inst_dmem_ram_70), .A2(MEM_stage_inst_dmem_n13622), .ZN(MEM_stage_inst_dmem_n13611) );
NAND2_X1 MEM_stage_inst_dmem_U10068 ( .A1(MEM_stage_inst_dmem_n13609), .A2(MEM_stage_inst_dmem_n13608), .ZN(MEM_stage_inst_dmem_n12418) );
NAND2_X1 MEM_stage_inst_dmem_U10067 ( .A1(MEM_stage_inst_dmem_n13886), .A2(MEM_stage_inst_dmem_n13623), .ZN(MEM_stage_inst_dmem_n13608) );
NAND2_X1 MEM_stage_inst_dmem_U10066 ( .A1(MEM_stage_inst_dmem_ram_71), .A2(MEM_stage_inst_dmem_n13622), .ZN(MEM_stage_inst_dmem_n13609) );
NAND2_X1 MEM_stage_inst_dmem_U10065 ( .A1(MEM_stage_inst_dmem_n13607), .A2(MEM_stage_inst_dmem_n13606), .ZN(MEM_stage_inst_dmem_n12419) );
NAND2_X1 MEM_stage_inst_dmem_U10064 ( .A1(MEM_stage_inst_dmem_n13883), .A2(MEM_stage_inst_dmem_n13623), .ZN(MEM_stage_inst_dmem_n13606) );
NAND2_X1 MEM_stage_inst_dmem_U10063 ( .A1(MEM_stage_inst_dmem_ram_72), .A2(MEM_stage_inst_dmem_n13622), .ZN(MEM_stage_inst_dmem_n13607) );
NAND2_X1 MEM_stage_inst_dmem_U10062 ( .A1(MEM_stage_inst_dmem_n13605), .A2(MEM_stage_inst_dmem_n13604), .ZN(MEM_stage_inst_dmem_n12420) );
NAND2_X1 MEM_stage_inst_dmem_U10061 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n13623), .ZN(MEM_stage_inst_dmem_n13604) );
NAND2_X1 MEM_stage_inst_dmem_U10060 ( .A1(MEM_stage_inst_dmem_ram_73), .A2(MEM_stage_inst_dmem_n13622), .ZN(MEM_stage_inst_dmem_n13605) );
NAND2_X1 MEM_stage_inst_dmem_U10059 ( .A1(MEM_stage_inst_dmem_n13603), .A2(MEM_stage_inst_dmem_n13602), .ZN(MEM_stage_inst_dmem_n12421) );
NAND2_X1 MEM_stage_inst_dmem_U10058 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n13623), .ZN(MEM_stage_inst_dmem_n13602) );
NAND2_X1 MEM_stage_inst_dmem_U10057 ( .A1(MEM_stage_inst_dmem_ram_74), .A2(MEM_stage_inst_dmem_n13622), .ZN(MEM_stage_inst_dmem_n13603) );
NAND2_X1 MEM_stage_inst_dmem_U10056 ( .A1(MEM_stage_inst_dmem_n13601), .A2(MEM_stage_inst_dmem_n13600), .ZN(MEM_stage_inst_dmem_n12422) );
NAND2_X1 MEM_stage_inst_dmem_U10055 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n13623), .ZN(MEM_stage_inst_dmem_n13600) );
NAND2_X1 MEM_stage_inst_dmem_U10054 ( .A1(MEM_stage_inst_dmem_ram_75), .A2(MEM_stage_inst_dmem_n13622), .ZN(MEM_stage_inst_dmem_n13601) );
NAND2_X1 MEM_stage_inst_dmem_U10053 ( .A1(MEM_stage_inst_dmem_n13599), .A2(MEM_stage_inst_dmem_n13598), .ZN(MEM_stage_inst_dmem_n12423) );
NAND2_X1 MEM_stage_inst_dmem_U10052 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n13623), .ZN(MEM_stage_inst_dmem_n13598) );
NAND2_X1 MEM_stage_inst_dmem_U10051 ( .A1(MEM_stage_inst_dmem_ram_76), .A2(MEM_stage_inst_dmem_n13622), .ZN(MEM_stage_inst_dmem_n13599) );
NAND2_X1 MEM_stage_inst_dmem_U10050 ( .A1(MEM_stage_inst_dmem_n13597), .A2(MEM_stage_inst_dmem_n13596), .ZN(MEM_stage_inst_dmem_n12424) );
NAND2_X1 MEM_stage_inst_dmem_U10049 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n13623), .ZN(MEM_stage_inst_dmem_n13596) );
NAND2_X1 MEM_stage_inst_dmem_U10048 ( .A1(MEM_stage_inst_dmem_ram_77), .A2(MEM_stage_inst_dmem_n13622), .ZN(MEM_stage_inst_dmem_n13597) );
NAND2_X1 MEM_stage_inst_dmem_U10047 ( .A1(MEM_stage_inst_dmem_n13595), .A2(MEM_stage_inst_dmem_n13594), .ZN(MEM_stage_inst_dmem_n12425) );
NAND2_X1 MEM_stage_inst_dmem_U10046 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n13623), .ZN(MEM_stage_inst_dmem_n13594) );
NAND2_X1 MEM_stage_inst_dmem_U10045 ( .A1(MEM_stage_inst_dmem_ram_78), .A2(MEM_stage_inst_dmem_n13622), .ZN(MEM_stage_inst_dmem_n13595) );
NAND2_X1 MEM_stage_inst_dmem_U10044 ( .A1(MEM_stage_inst_dmem_n13593), .A2(MEM_stage_inst_dmem_n13592), .ZN(MEM_stage_inst_dmem_n12426) );
NAND2_X1 MEM_stage_inst_dmem_U10043 ( .A1(MEM_stage_inst_dmem_n16758), .A2(MEM_stage_inst_dmem_n13623), .ZN(MEM_stage_inst_dmem_n13592) );
INV_X1 MEM_stage_inst_dmem_U10042 ( .A(MEM_stage_inst_dmem_n13622), .ZN(MEM_stage_inst_dmem_n13623) );
NAND2_X1 MEM_stage_inst_dmem_U10041 ( .A1(MEM_stage_inst_dmem_ram_79), .A2(MEM_stage_inst_dmem_n13622), .ZN(MEM_stage_inst_dmem_n13593) );
NAND2_X1 MEM_stage_inst_dmem_U10040 ( .A1(MEM_stage_inst_dmem_n21319), .A2(MEM_stage_inst_dmem_n13728), .ZN(MEM_stage_inst_dmem_n13622) );
NAND2_X1 MEM_stage_inst_dmem_U10039 ( .A1(MEM_stage_inst_dmem_n13591), .A2(MEM_stage_inst_dmem_n13590), .ZN(MEM_stage_inst_dmem_n12427) );
NAND2_X1 MEM_stage_inst_dmem_U10038 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n13589), .ZN(MEM_stage_inst_dmem_n13590) );
NAND2_X1 MEM_stage_inst_dmem_U10037 ( .A1(MEM_stage_inst_dmem_ram_80), .A2(MEM_stage_inst_dmem_n13588), .ZN(MEM_stage_inst_dmem_n13591) );
NAND2_X1 MEM_stage_inst_dmem_U10036 ( .A1(MEM_stage_inst_dmem_n13587), .A2(MEM_stage_inst_dmem_n13586), .ZN(MEM_stage_inst_dmem_n12428) );
NAND2_X1 MEM_stage_inst_dmem_U10035 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n13589), .ZN(MEM_stage_inst_dmem_n13586) );
NAND2_X1 MEM_stage_inst_dmem_U10034 ( .A1(MEM_stage_inst_dmem_ram_81), .A2(MEM_stage_inst_dmem_n13588), .ZN(MEM_stage_inst_dmem_n13587) );
NAND2_X1 MEM_stage_inst_dmem_U10033 ( .A1(MEM_stage_inst_dmem_n13585), .A2(MEM_stage_inst_dmem_n13584), .ZN(MEM_stage_inst_dmem_n12429) );
NAND2_X1 MEM_stage_inst_dmem_U10032 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n13589), .ZN(MEM_stage_inst_dmem_n13584) );
NAND2_X1 MEM_stage_inst_dmem_U10031 ( .A1(MEM_stage_inst_dmem_ram_82), .A2(MEM_stage_inst_dmem_n13588), .ZN(MEM_stage_inst_dmem_n13585) );
NAND2_X1 MEM_stage_inst_dmem_U10030 ( .A1(MEM_stage_inst_dmem_n13583), .A2(MEM_stage_inst_dmem_n13582), .ZN(MEM_stage_inst_dmem_n12430) );
NAND2_X1 MEM_stage_inst_dmem_U10029 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n13589), .ZN(MEM_stage_inst_dmem_n13582) );
NAND2_X1 MEM_stage_inst_dmem_U10028 ( .A1(MEM_stage_inst_dmem_ram_83), .A2(MEM_stage_inst_dmem_n13588), .ZN(MEM_stage_inst_dmem_n13583) );
NAND2_X1 MEM_stage_inst_dmem_U10027 ( .A1(MEM_stage_inst_dmem_n13581), .A2(MEM_stage_inst_dmem_n13580), .ZN(MEM_stage_inst_dmem_n12431) );
NAND2_X1 MEM_stage_inst_dmem_U10026 ( .A1(MEM_stage_inst_dmem_n16368), .A2(MEM_stage_inst_dmem_n13589), .ZN(MEM_stage_inst_dmem_n13580) );
NAND2_X1 MEM_stage_inst_dmem_U10025 ( .A1(MEM_stage_inst_dmem_ram_84), .A2(MEM_stage_inst_dmem_n13588), .ZN(MEM_stage_inst_dmem_n13581) );
NAND2_X1 MEM_stage_inst_dmem_U10024 ( .A1(MEM_stage_inst_dmem_n13579), .A2(MEM_stage_inst_dmem_n13578), .ZN(MEM_stage_inst_dmem_n12432) );
NAND2_X1 MEM_stage_inst_dmem_U10023 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n13589), .ZN(MEM_stage_inst_dmem_n13578) );
NAND2_X1 MEM_stage_inst_dmem_U10022 ( .A1(MEM_stage_inst_dmem_ram_85), .A2(MEM_stage_inst_dmem_n13588), .ZN(MEM_stage_inst_dmem_n13579) );
NAND2_X1 MEM_stage_inst_dmem_U10021 ( .A1(MEM_stage_inst_dmem_n13577), .A2(MEM_stage_inst_dmem_n13576), .ZN(MEM_stage_inst_dmem_n12433) );
NAND2_X1 MEM_stage_inst_dmem_U10020 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n13589), .ZN(MEM_stage_inst_dmem_n13576) );
NAND2_X1 MEM_stage_inst_dmem_U10019 ( .A1(MEM_stage_inst_dmem_ram_86), .A2(MEM_stage_inst_dmem_n13588), .ZN(MEM_stage_inst_dmem_n13577) );
NAND2_X1 MEM_stage_inst_dmem_U10018 ( .A1(MEM_stage_inst_dmem_n13575), .A2(MEM_stage_inst_dmem_n13574), .ZN(MEM_stage_inst_dmem_n12434) );
NAND2_X1 MEM_stage_inst_dmem_U10017 ( .A1(MEM_stage_inst_dmem_n13886), .A2(MEM_stage_inst_dmem_n13589), .ZN(MEM_stage_inst_dmem_n13574) );
NAND2_X1 MEM_stage_inst_dmem_U10016 ( .A1(MEM_stage_inst_dmem_ram_87), .A2(MEM_stage_inst_dmem_n13588), .ZN(MEM_stage_inst_dmem_n13575) );
NAND2_X1 MEM_stage_inst_dmem_U10015 ( .A1(MEM_stage_inst_dmem_n13573), .A2(MEM_stage_inst_dmem_n13572), .ZN(MEM_stage_inst_dmem_n12435) );
NAND2_X1 MEM_stage_inst_dmem_U10014 ( .A1(MEM_stage_inst_dmem_n13883), .A2(MEM_stage_inst_dmem_n13589), .ZN(MEM_stage_inst_dmem_n13572) );
NAND2_X1 MEM_stage_inst_dmem_U10013 ( .A1(MEM_stage_inst_dmem_ram_88), .A2(MEM_stage_inst_dmem_n13588), .ZN(MEM_stage_inst_dmem_n13573) );
NAND2_X1 MEM_stage_inst_dmem_U10012 ( .A1(MEM_stage_inst_dmem_n13571), .A2(MEM_stage_inst_dmem_n13570), .ZN(MEM_stage_inst_dmem_n12436) );
NAND2_X1 MEM_stage_inst_dmem_U10011 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n13589), .ZN(MEM_stage_inst_dmem_n13570) );
NAND2_X1 MEM_stage_inst_dmem_U10010 ( .A1(MEM_stage_inst_dmem_ram_89), .A2(MEM_stage_inst_dmem_n13588), .ZN(MEM_stage_inst_dmem_n13571) );
NAND2_X1 MEM_stage_inst_dmem_U10009 ( .A1(MEM_stage_inst_dmem_n13569), .A2(MEM_stage_inst_dmem_n13568), .ZN(MEM_stage_inst_dmem_n12437) );
NAND2_X1 MEM_stage_inst_dmem_U10008 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n13589), .ZN(MEM_stage_inst_dmem_n13568) );
NAND2_X1 MEM_stage_inst_dmem_U10007 ( .A1(MEM_stage_inst_dmem_ram_90), .A2(MEM_stage_inst_dmem_n13588), .ZN(MEM_stage_inst_dmem_n13569) );
NAND2_X1 MEM_stage_inst_dmem_U10006 ( .A1(MEM_stage_inst_dmem_n13567), .A2(MEM_stage_inst_dmem_n13566), .ZN(MEM_stage_inst_dmem_n12438) );
NAND2_X1 MEM_stage_inst_dmem_U10005 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n13589), .ZN(MEM_stage_inst_dmem_n13566) );
NAND2_X1 MEM_stage_inst_dmem_U10004 ( .A1(MEM_stage_inst_dmem_ram_91), .A2(MEM_stage_inst_dmem_n13588), .ZN(MEM_stage_inst_dmem_n13567) );
NAND2_X1 MEM_stage_inst_dmem_U10003 ( .A1(MEM_stage_inst_dmem_n13565), .A2(MEM_stage_inst_dmem_n13564), .ZN(MEM_stage_inst_dmem_n12439) );
NAND2_X1 MEM_stage_inst_dmem_U10002 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n13589), .ZN(MEM_stage_inst_dmem_n13564) );
NAND2_X1 MEM_stage_inst_dmem_U10001 ( .A1(MEM_stage_inst_dmem_ram_92), .A2(MEM_stage_inst_dmem_n13588), .ZN(MEM_stage_inst_dmem_n13565) );
NAND2_X1 MEM_stage_inst_dmem_U10000 ( .A1(MEM_stage_inst_dmem_n13563), .A2(MEM_stage_inst_dmem_n13562), .ZN(MEM_stage_inst_dmem_n12440) );
NAND2_X1 MEM_stage_inst_dmem_U9999 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n13589), .ZN(MEM_stage_inst_dmem_n13562) );
NAND2_X1 MEM_stage_inst_dmem_U9998 ( .A1(MEM_stage_inst_dmem_ram_93), .A2(MEM_stage_inst_dmem_n13588), .ZN(MEM_stage_inst_dmem_n13563) );
NAND2_X1 MEM_stage_inst_dmem_U9997 ( .A1(MEM_stage_inst_dmem_n13561), .A2(MEM_stage_inst_dmem_n13560), .ZN(MEM_stage_inst_dmem_n12441) );
NAND2_X1 MEM_stage_inst_dmem_U9996 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n13589), .ZN(MEM_stage_inst_dmem_n13560) );
NAND2_X1 MEM_stage_inst_dmem_U9995 ( .A1(MEM_stage_inst_dmem_ram_94), .A2(MEM_stage_inst_dmem_n13588), .ZN(MEM_stage_inst_dmem_n13561) );
NAND2_X1 MEM_stage_inst_dmem_U9994 ( .A1(MEM_stage_inst_dmem_n13559), .A2(MEM_stage_inst_dmem_n13558), .ZN(MEM_stage_inst_dmem_n12442) );
NAND2_X1 MEM_stage_inst_dmem_U9993 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n13589), .ZN(MEM_stage_inst_dmem_n13558) );
INV_X1 MEM_stage_inst_dmem_U9992 ( .A(MEM_stage_inst_dmem_n13588), .ZN(MEM_stage_inst_dmem_n13589) );
NAND2_X1 MEM_stage_inst_dmem_U9991 ( .A1(MEM_stage_inst_dmem_ram_95), .A2(MEM_stage_inst_dmem_n13588), .ZN(MEM_stage_inst_dmem_n13559) );
NAND2_X1 MEM_stage_inst_dmem_U9990 ( .A1(MEM_stage_inst_dmem_n21284), .A2(MEM_stage_inst_dmem_n13728), .ZN(MEM_stage_inst_dmem_n13588) );
NAND2_X1 MEM_stage_inst_dmem_U9989 ( .A1(MEM_stage_inst_dmem_n13557), .A2(MEM_stage_inst_dmem_n13556), .ZN(MEM_stage_inst_dmem_n12443) );
NAND2_X1 MEM_stage_inst_dmem_U9988 ( .A1(MEM_stage_inst_dmem_n15145), .A2(MEM_stage_inst_dmem_n13555), .ZN(MEM_stage_inst_dmem_n13556) );
NAND2_X1 MEM_stage_inst_dmem_U9987 ( .A1(MEM_stage_inst_dmem_ram_96), .A2(MEM_stage_inst_dmem_n13554), .ZN(MEM_stage_inst_dmem_n13557) );
NAND2_X1 MEM_stage_inst_dmem_U9986 ( .A1(MEM_stage_inst_dmem_n13553), .A2(MEM_stage_inst_dmem_n13552), .ZN(MEM_stage_inst_dmem_n12444) );
NAND2_X1 MEM_stage_inst_dmem_U9985 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n13555), .ZN(MEM_stage_inst_dmem_n13552) );
NAND2_X1 MEM_stage_inst_dmem_U9984 ( .A1(MEM_stage_inst_dmem_ram_97), .A2(MEM_stage_inst_dmem_n13554), .ZN(MEM_stage_inst_dmem_n13553) );
NAND2_X1 MEM_stage_inst_dmem_U9983 ( .A1(MEM_stage_inst_dmem_n13551), .A2(MEM_stage_inst_dmem_n13550), .ZN(MEM_stage_inst_dmem_n12445) );
NAND2_X1 MEM_stage_inst_dmem_U9982 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n13555), .ZN(MEM_stage_inst_dmem_n13550) );
NAND2_X1 MEM_stage_inst_dmem_U9981 ( .A1(MEM_stage_inst_dmem_ram_98), .A2(MEM_stage_inst_dmem_n13554), .ZN(MEM_stage_inst_dmem_n13551) );
NAND2_X1 MEM_stage_inst_dmem_U9980 ( .A1(MEM_stage_inst_dmem_n13549), .A2(MEM_stage_inst_dmem_n13548), .ZN(MEM_stage_inst_dmem_n12446) );
NAND2_X1 MEM_stage_inst_dmem_U9979 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n13555), .ZN(MEM_stage_inst_dmem_n13548) );
NAND2_X1 MEM_stage_inst_dmem_U9978 ( .A1(MEM_stage_inst_dmem_ram_99), .A2(MEM_stage_inst_dmem_n13554), .ZN(MEM_stage_inst_dmem_n13549) );
NAND2_X1 MEM_stage_inst_dmem_U9977 ( .A1(MEM_stage_inst_dmem_n13547), .A2(MEM_stage_inst_dmem_n13546), .ZN(MEM_stage_inst_dmem_n12447) );
NAND2_X1 MEM_stage_inst_dmem_U9976 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n13555), .ZN(MEM_stage_inst_dmem_n13546) );
NAND2_X1 MEM_stage_inst_dmem_U9975 ( .A1(MEM_stage_inst_dmem_ram_100), .A2(MEM_stage_inst_dmem_n13554), .ZN(MEM_stage_inst_dmem_n13547) );
NAND2_X1 MEM_stage_inst_dmem_U9974 ( .A1(MEM_stage_inst_dmem_n13545), .A2(MEM_stage_inst_dmem_n13544), .ZN(MEM_stage_inst_dmem_n12448) );
NAND2_X1 MEM_stage_inst_dmem_U9973 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n13555), .ZN(MEM_stage_inst_dmem_n13544) );
NAND2_X1 MEM_stage_inst_dmem_U9972 ( .A1(MEM_stage_inst_dmem_ram_101), .A2(MEM_stage_inst_dmem_n13554), .ZN(MEM_stage_inst_dmem_n13545) );
NAND2_X1 MEM_stage_inst_dmem_U9971 ( .A1(MEM_stage_inst_dmem_n13543), .A2(MEM_stage_inst_dmem_n13542), .ZN(MEM_stage_inst_dmem_n12449) );
NAND2_X1 MEM_stage_inst_dmem_U9970 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n13555), .ZN(MEM_stage_inst_dmem_n13542) );
NAND2_X1 MEM_stage_inst_dmem_U9969 ( .A1(MEM_stage_inst_dmem_ram_102), .A2(MEM_stage_inst_dmem_n13554), .ZN(MEM_stage_inst_dmem_n13543) );
NAND2_X1 MEM_stage_inst_dmem_U9968 ( .A1(MEM_stage_inst_dmem_n13541), .A2(MEM_stage_inst_dmem_n13540), .ZN(MEM_stage_inst_dmem_n12450) );
NAND2_X1 MEM_stage_inst_dmem_U9967 ( .A1(MEM_stage_inst_dmem_n13886), .A2(MEM_stage_inst_dmem_n13555), .ZN(MEM_stage_inst_dmem_n13540) );
NAND2_X1 MEM_stage_inst_dmem_U9966 ( .A1(MEM_stage_inst_dmem_ram_103), .A2(MEM_stage_inst_dmem_n13554), .ZN(MEM_stage_inst_dmem_n13541) );
NAND2_X1 MEM_stage_inst_dmem_U9965 ( .A1(MEM_stage_inst_dmem_n13539), .A2(MEM_stage_inst_dmem_n13538), .ZN(MEM_stage_inst_dmem_n12451) );
NAND2_X1 MEM_stage_inst_dmem_U9964 ( .A1(MEM_stage_inst_dmem_n13883), .A2(MEM_stage_inst_dmem_n13555), .ZN(MEM_stage_inst_dmem_n13538) );
NAND2_X1 MEM_stage_inst_dmem_U9963 ( .A1(MEM_stage_inst_dmem_ram_104), .A2(MEM_stage_inst_dmem_n13554), .ZN(MEM_stage_inst_dmem_n13539) );
NAND2_X1 MEM_stage_inst_dmem_U9962 ( .A1(MEM_stage_inst_dmem_n13537), .A2(MEM_stage_inst_dmem_n13536), .ZN(MEM_stage_inst_dmem_n12452) );
NAND2_X1 MEM_stage_inst_dmem_U9961 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n13555), .ZN(MEM_stage_inst_dmem_n13536) );
NAND2_X1 MEM_stage_inst_dmem_U9960 ( .A1(MEM_stage_inst_dmem_ram_105), .A2(MEM_stage_inst_dmem_n13554), .ZN(MEM_stage_inst_dmem_n13537) );
NAND2_X1 MEM_stage_inst_dmem_U9959 ( .A1(MEM_stage_inst_dmem_n13535), .A2(MEM_stage_inst_dmem_n13534), .ZN(MEM_stage_inst_dmem_n12453) );
NAND2_X1 MEM_stage_inst_dmem_U9958 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n13555), .ZN(MEM_stage_inst_dmem_n13534) );
NAND2_X1 MEM_stage_inst_dmem_U9957 ( .A1(MEM_stage_inst_dmem_ram_106), .A2(MEM_stage_inst_dmem_n13554), .ZN(MEM_stage_inst_dmem_n13535) );
NAND2_X1 MEM_stage_inst_dmem_U9956 ( .A1(MEM_stage_inst_dmem_n13533), .A2(MEM_stage_inst_dmem_n13532), .ZN(MEM_stage_inst_dmem_n12454) );
NAND2_X1 MEM_stage_inst_dmem_U9955 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n13555), .ZN(MEM_stage_inst_dmem_n13532) );
NAND2_X1 MEM_stage_inst_dmem_U9954 ( .A1(MEM_stage_inst_dmem_ram_107), .A2(MEM_stage_inst_dmem_n13554), .ZN(MEM_stage_inst_dmem_n13533) );
NAND2_X1 MEM_stage_inst_dmem_U9953 ( .A1(MEM_stage_inst_dmem_n13531), .A2(MEM_stage_inst_dmem_n13530), .ZN(MEM_stage_inst_dmem_n12455) );
NAND2_X1 MEM_stage_inst_dmem_U9952 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n13555), .ZN(MEM_stage_inst_dmem_n13530) );
NAND2_X1 MEM_stage_inst_dmem_U9951 ( .A1(MEM_stage_inst_dmem_ram_108), .A2(MEM_stage_inst_dmem_n13554), .ZN(MEM_stage_inst_dmem_n13531) );
NAND2_X1 MEM_stage_inst_dmem_U9950 ( .A1(MEM_stage_inst_dmem_n13529), .A2(MEM_stage_inst_dmem_n13528), .ZN(MEM_stage_inst_dmem_n12456) );
NAND2_X1 MEM_stage_inst_dmem_U9949 ( .A1(MEM_stage_inst_dmem_n15116), .A2(MEM_stage_inst_dmem_n13555), .ZN(MEM_stage_inst_dmem_n13528) );
NAND2_X1 MEM_stage_inst_dmem_U9948 ( .A1(MEM_stage_inst_dmem_ram_109), .A2(MEM_stage_inst_dmem_n13554), .ZN(MEM_stage_inst_dmem_n13529) );
NAND2_X1 MEM_stage_inst_dmem_U9947 ( .A1(MEM_stage_inst_dmem_n13527), .A2(MEM_stage_inst_dmem_n13526), .ZN(MEM_stage_inst_dmem_n12457) );
NAND2_X1 MEM_stage_inst_dmem_U9946 ( .A1(MEM_stage_inst_dmem_n15113), .A2(MEM_stage_inst_dmem_n13555), .ZN(MEM_stage_inst_dmem_n13526) );
NAND2_X1 MEM_stage_inst_dmem_U9945 ( .A1(MEM_stage_inst_dmem_ram_110), .A2(MEM_stage_inst_dmem_n13554), .ZN(MEM_stage_inst_dmem_n13527) );
NAND2_X1 MEM_stage_inst_dmem_U9944 ( .A1(MEM_stage_inst_dmem_n13525), .A2(MEM_stage_inst_dmem_n13524), .ZN(MEM_stage_inst_dmem_n12458) );
NAND2_X1 MEM_stage_inst_dmem_U9943 ( .A1(MEM_stage_inst_dmem_n16343), .A2(MEM_stage_inst_dmem_n13555), .ZN(MEM_stage_inst_dmem_n13524) );
INV_X1 MEM_stage_inst_dmem_U9942 ( .A(MEM_stage_inst_dmem_n13554), .ZN(MEM_stage_inst_dmem_n13555) );
NAND2_X1 MEM_stage_inst_dmem_U9941 ( .A1(MEM_stage_inst_dmem_ram_111), .A2(MEM_stage_inst_dmem_n13554), .ZN(MEM_stage_inst_dmem_n13525) );
NAND2_X1 MEM_stage_inst_dmem_U9940 ( .A1(MEM_stage_inst_dmem_n21249), .A2(MEM_stage_inst_dmem_n13728), .ZN(MEM_stage_inst_dmem_n13554) );
NAND2_X1 MEM_stage_inst_dmem_U9939 ( .A1(MEM_stage_inst_dmem_n13523), .A2(MEM_stage_inst_dmem_n13522), .ZN(MEM_stage_inst_dmem_n12459) );
NAND2_X1 MEM_stage_inst_dmem_U9938 ( .A1(MEM_stage_inst_dmem_n19275), .A2(MEM_stage_inst_dmem_n13521), .ZN(MEM_stage_inst_dmem_n13522) );
NAND2_X1 MEM_stage_inst_dmem_U9937 ( .A1(MEM_stage_inst_dmem_ram_112), .A2(MEM_stage_inst_dmem_n13520), .ZN(MEM_stage_inst_dmem_n13523) );
NAND2_X1 MEM_stage_inst_dmem_U9936 ( .A1(MEM_stage_inst_dmem_n13519), .A2(MEM_stage_inst_dmem_n13518), .ZN(MEM_stage_inst_dmem_n12460) );
NAND2_X1 MEM_stage_inst_dmem_U9935 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n13521), .ZN(MEM_stage_inst_dmem_n13518) );
NAND2_X1 MEM_stage_inst_dmem_U9934 ( .A1(MEM_stage_inst_dmem_ram_113), .A2(MEM_stage_inst_dmem_n13520), .ZN(MEM_stage_inst_dmem_n13519) );
NAND2_X1 MEM_stage_inst_dmem_U9933 ( .A1(MEM_stage_inst_dmem_n13517), .A2(MEM_stage_inst_dmem_n13516), .ZN(MEM_stage_inst_dmem_n12461) );
NAND2_X1 MEM_stage_inst_dmem_U9932 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n13521), .ZN(MEM_stage_inst_dmem_n13516) );
NAND2_X1 MEM_stage_inst_dmem_U9931 ( .A1(MEM_stage_inst_dmem_ram_114), .A2(MEM_stage_inst_dmem_n13520), .ZN(MEM_stage_inst_dmem_n13517) );
NAND2_X1 MEM_stage_inst_dmem_U9930 ( .A1(MEM_stage_inst_dmem_n13515), .A2(MEM_stage_inst_dmem_n13514), .ZN(MEM_stage_inst_dmem_n12462) );
NAND2_X1 MEM_stage_inst_dmem_U9929 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n13521), .ZN(MEM_stage_inst_dmem_n13514) );
NAND2_X1 MEM_stage_inst_dmem_U9928 ( .A1(MEM_stage_inst_dmem_ram_115), .A2(MEM_stage_inst_dmem_n13520), .ZN(MEM_stage_inst_dmem_n13515) );
NAND2_X1 MEM_stage_inst_dmem_U9927 ( .A1(MEM_stage_inst_dmem_n13513), .A2(MEM_stage_inst_dmem_n13512), .ZN(MEM_stage_inst_dmem_n12463) );
NAND2_X1 MEM_stage_inst_dmem_U9926 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n13521), .ZN(MEM_stage_inst_dmem_n13512) );
NAND2_X1 MEM_stage_inst_dmem_U9925 ( .A1(MEM_stage_inst_dmem_ram_116), .A2(MEM_stage_inst_dmem_n13520), .ZN(MEM_stage_inst_dmem_n13513) );
NAND2_X1 MEM_stage_inst_dmem_U9924 ( .A1(MEM_stage_inst_dmem_n13511), .A2(MEM_stage_inst_dmem_n13510), .ZN(MEM_stage_inst_dmem_n12464) );
NAND2_X1 MEM_stage_inst_dmem_U9923 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n13521), .ZN(MEM_stage_inst_dmem_n13510) );
NAND2_X1 MEM_stage_inst_dmem_U9922 ( .A1(MEM_stage_inst_dmem_ram_117), .A2(MEM_stage_inst_dmem_n13520), .ZN(MEM_stage_inst_dmem_n13511) );
NAND2_X1 MEM_stage_inst_dmem_U9921 ( .A1(MEM_stage_inst_dmem_n13509), .A2(MEM_stage_inst_dmem_n13508), .ZN(MEM_stage_inst_dmem_n12465) );
NAND2_X1 MEM_stage_inst_dmem_U9920 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n13521), .ZN(MEM_stage_inst_dmem_n13508) );
NAND2_X1 MEM_stage_inst_dmem_U9919 ( .A1(MEM_stage_inst_dmem_ram_118), .A2(MEM_stage_inst_dmem_n13520), .ZN(MEM_stage_inst_dmem_n13509) );
NAND2_X1 MEM_stage_inst_dmem_U9918 ( .A1(MEM_stage_inst_dmem_n13507), .A2(MEM_stage_inst_dmem_n13506), .ZN(MEM_stage_inst_dmem_n12466) );
NAND2_X1 MEM_stage_inst_dmem_U9917 ( .A1(MEM_stage_inst_dmem_n17), .A2(MEM_stage_inst_dmem_n13521), .ZN(MEM_stage_inst_dmem_n13506) );
NAND2_X1 MEM_stage_inst_dmem_U9916 ( .A1(MEM_stage_inst_dmem_ram_119), .A2(MEM_stage_inst_dmem_n13520), .ZN(MEM_stage_inst_dmem_n13507) );
NAND2_X1 MEM_stage_inst_dmem_U9915 ( .A1(MEM_stage_inst_dmem_n13505), .A2(MEM_stage_inst_dmem_n13504), .ZN(MEM_stage_inst_dmem_n12467) );
NAND2_X1 MEM_stage_inst_dmem_U9914 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n13521), .ZN(MEM_stage_inst_dmem_n13504) );
NAND2_X1 MEM_stage_inst_dmem_U9913 ( .A1(MEM_stage_inst_dmem_ram_120), .A2(MEM_stage_inst_dmem_n13520), .ZN(MEM_stage_inst_dmem_n13505) );
NAND2_X1 MEM_stage_inst_dmem_U9912 ( .A1(MEM_stage_inst_dmem_n13503), .A2(MEM_stage_inst_dmem_n13502), .ZN(MEM_stage_inst_dmem_n12468) );
NAND2_X1 MEM_stage_inst_dmem_U9911 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n13521), .ZN(MEM_stage_inst_dmem_n13502) );
NAND2_X1 MEM_stage_inst_dmem_U9910 ( .A1(MEM_stage_inst_dmem_ram_121), .A2(MEM_stage_inst_dmem_n13520), .ZN(MEM_stage_inst_dmem_n13503) );
NAND2_X1 MEM_stage_inst_dmem_U9909 ( .A1(MEM_stage_inst_dmem_n13501), .A2(MEM_stage_inst_dmem_n13500), .ZN(MEM_stage_inst_dmem_n12469) );
NAND2_X1 MEM_stage_inst_dmem_U9908 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n13521), .ZN(MEM_stage_inst_dmem_n13500) );
NAND2_X1 MEM_stage_inst_dmem_U9907 ( .A1(MEM_stage_inst_dmem_ram_122), .A2(MEM_stage_inst_dmem_n13520), .ZN(MEM_stage_inst_dmem_n13501) );
NAND2_X1 MEM_stage_inst_dmem_U9906 ( .A1(MEM_stage_inst_dmem_n13499), .A2(MEM_stage_inst_dmem_n13498), .ZN(MEM_stage_inst_dmem_n12470) );
NAND2_X1 MEM_stage_inst_dmem_U9905 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n13521), .ZN(MEM_stage_inst_dmem_n13498) );
NAND2_X1 MEM_stage_inst_dmem_U9904 ( .A1(MEM_stage_inst_dmem_ram_123), .A2(MEM_stage_inst_dmem_n13520), .ZN(MEM_stage_inst_dmem_n13499) );
NAND2_X1 MEM_stage_inst_dmem_U9903 ( .A1(MEM_stage_inst_dmem_n13497), .A2(MEM_stage_inst_dmem_n13496), .ZN(MEM_stage_inst_dmem_n12471) );
NAND2_X1 MEM_stage_inst_dmem_U9902 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n13521), .ZN(MEM_stage_inst_dmem_n13496) );
NAND2_X1 MEM_stage_inst_dmem_U9901 ( .A1(MEM_stage_inst_dmem_ram_124), .A2(MEM_stage_inst_dmem_n13520), .ZN(MEM_stage_inst_dmem_n13497) );
NAND2_X1 MEM_stage_inst_dmem_U9900 ( .A1(MEM_stage_inst_dmem_n13495), .A2(MEM_stage_inst_dmem_n13494), .ZN(MEM_stage_inst_dmem_n12472) );
NAND2_X1 MEM_stage_inst_dmem_U9899 ( .A1(MEM_stage_inst_dmem_n19242), .A2(MEM_stage_inst_dmem_n13521), .ZN(MEM_stage_inst_dmem_n13494) );
NAND2_X1 MEM_stage_inst_dmem_U9898 ( .A1(MEM_stage_inst_dmem_ram_125), .A2(MEM_stage_inst_dmem_n13520), .ZN(MEM_stage_inst_dmem_n13495) );
NAND2_X1 MEM_stage_inst_dmem_U9897 ( .A1(MEM_stage_inst_dmem_n13493), .A2(MEM_stage_inst_dmem_n13492), .ZN(MEM_stage_inst_dmem_n12473) );
NAND2_X1 MEM_stage_inst_dmem_U9896 ( .A1(MEM_stage_inst_dmem_n115), .A2(MEM_stage_inst_dmem_n13521), .ZN(MEM_stage_inst_dmem_n13492) );
NAND2_X1 MEM_stage_inst_dmem_U9895 ( .A1(MEM_stage_inst_dmem_ram_126), .A2(MEM_stage_inst_dmem_n13520), .ZN(MEM_stage_inst_dmem_n13493) );
NAND2_X1 MEM_stage_inst_dmem_U9894 ( .A1(MEM_stage_inst_dmem_n13491), .A2(MEM_stage_inst_dmem_n13490), .ZN(MEM_stage_inst_dmem_n12474) );
NAND2_X1 MEM_stage_inst_dmem_U9893 ( .A1(MEM_stage_inst_dmem_n16758), .A2(MEM_stage_inst_dmem_n13521), .ZN(MEM_stage_inst_dmem_n13490) );
INV_X1 MEM_stage_inst_dmem_U9892 ( .A(MEM_stage_inst_dmem_n13520), .ZN(MEM_stage_inst_dmem_n13521) );
NAND2_X1 MEM_stage_inst_dmem_U9891 ( .A1(MEM_stage_inst_dmem_ram_127), .A2(MEM_stage_inst_dmem_n13520), .ZN(MEM_stage_inst_dmem_n13491) );
NAND2_X1 MEM_stage_inst_dmem_U9890 ( .A1(MEM_stage_inst_dmem_n21214), .A2(MEM_stage_inst_dmem_n13728), .ZN(MEM_stage_inst_dmem_n13520) );
NAND2_X1 MEM_stage_inst_dmem_U9889 ( .A1(MEM_stage_inst_dmem_n13489), .A2(MEM_stage_inst_dmem_n13488), .ZN(MEM_stage_inst_dmem_n12475) );
NAND2_X1 MEM_stage_inst_dmem_U9888 ( .A1(MEM_stage_inst_dmem_n14732), .A2(MEM_stage_inst_dmem_n13487), .ZN(MEM_stage_inst_dmem_n13488) );
NAND2_X1 MEM_stage_inst_dmem_U9887 ( .A1(MEM_stage_inst_dmem_ram_128), .A2(MEM_stage_inst_dmem_n13486), .ZN(MEM_stage_inst_dmem_n13489) );
NAND2_X1 MEM_stage_inst_dmem_U9886 ( .A1(MEM_stage_inst_dmem_n13485), .A2(MEM_stage_inst_dmem_n13484), .ZN(MEM_stage_inst_dmem_n12476) );
NAND2_X1 MEM_stage_inst_dmem_U9885 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n13487), .ZN(MEM_stage_inst_dmem_n13484) );
NAND2_X1 MEM_stage_inst_dmem_U9884 ( .A1(MEM_stage_inst_dmem_ram_129), .A2(MEM_stage_inst_dmem_n13486), .ZN(MEM_stage_inst_dmem_n13485) );
NAND2_X1 MEM_stage_inst_dmem_U9883 ( .A1(MEM_stage_inst_dmem_n13483), .A2(MEM_stage_inst_dmem_n13482), .ZN(MEM_stage_inst_dmem_n12477) );
NAND2_X1 MEM_stage_inst_dmem_U9882 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n13487), .ZN(MEM_stage_inst_dmem_n13482) );
NAND2_X1 MEM_stage_inst_dmem_U9881 ( .A1(MEM_stage_inst_dmem_ram_130), .A2(MEM_stage_inst_dmem_n13486), .ZN(MEM_stage_inst_dmem_n13483) );
NAND2_X1 MEM_stage_inst_dmem_U9880 ( .A1(MEM_stage_inst_dmem_n13481), .A2(MEM_stage_inst_dmem_n13480), .ZN(MEM_stage_inst_dmem_n12478) );
NAND2_X1 MEM_stage_inst_dmem_U9879 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n13487), .ZN(MEM_stage_inst_dmem_n13480) );
NAND2_X1 MEM_stage_inst_dmem_U9878 ( .A1(MEM_stage_inst_dmem_ram_131), .A2(MEM_stage_inst_dmem_n13486), .ZN(MEM_stage_inst_dmem_n13481) );
NAND2_X1 MEM_stage_inst_dmem_U9877 ( .A1(MEM_stage_inst_dmem_n13479), .A2(MEM_stage_inst_dmem_n13478), .ZN(MEM_stage_inst_dmem_n12479) );
NAND2_X1 MEM_stage_inst_dmem_U9876 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n13487), .ZN(MEM_stage_inst_dmem_n13478) );
NAND2_X1 MEM_stage_inst_dmem_U9875 ( .A1(MEM_stage_inst_dmem_ram_132), .A2(MEM_stage_inst_dmem_n13486), .ZN(MEM_stage_inst_dmem_n13479) );
NAND2_X1 MEM_stage_inst_dmem_U9874 ( .A1(MEM_stage_inst_dmem_n13477), .A2(MEM_stage_inst_dmem_n13476), .ZN(MEM_stage_inst_dmem_n12480) );
NAND2_X1 MEM_stage_inst_dmem_U9873 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n13487), .ZN(MEM_stage_inst_dmem_n13476) );
NAND2_X1 MEM_stage_inst_dmem_U9872 ( .A1(MEM_stage_inst_dmem_ram_133), .A2(MEM_stage_inst_dmem_n13486), .ZN(MEM_stage_inst_dmem_n13477) );
NAND2_X1 MEM_stage_inst_dmem_U9871 ( .A1(MEM_stage_inst_dmem_n13475), .A2(MEM_stage_inst_dmem_n13474), .ZN(MEM_stage_inst_dmem_n12481) );
NAND2_X1 MEM_stage_inst_dmem_U9870 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n13487), .ZN(MEM_stage_inst_dmem_n13474) );
NAND2_X1 MEM_stage_inst_dmem_U9869 ( .A1(MEM_stage_inst_dmem_ram_134), .A2(MEM_stage_inst_dmem_n13486), .ZN(MEM_stage_inst_dmem_n13475) );
NAND2_X1 MEM_stage_inst_dmem_U9868 ( .A1(MEM_stage_inst_dmem_n13473), .A2(MEM_stage_inst_dmem_n13472), .ZN(MEM_stage_inst_dmem_n12482) );
NAND2_X1 MEM_stage_inst_dmem_U9867 ( .A1(MEM_stage_inst_dmem_n13886), .A2(MEM_stage_inst_dmem_n13487), .ZN(MEM_stage_inst_dmem_n13472) );
NAND2_X1 MEM_stage_inst_dmem_U9866 ( .A1(MEM_stage_inst_dmem_ram_135), .A2(MEM_stage_inst_dmem_n13486), .ZN(MEM_stage_inst_dmem_n13473) );
NAND2_X1 MEM_stage_inst_dmem_U9865 ( .A1(MEM_stage_inst_dmem_n13471), .A2(MEM_stage_inst_dmem_n13470), .ZN(MEM_stage_inst_dmem_n12483) );
NAND2_X1 MEM_stage_inst_dmem_U9864 ( .A1(MEM_stage_inst_dmem_n13883), .A2(MEM_stage_inst_dmem_n13487), .ZN(MEM_stage_inst_dmem_n13470) );
NAND2_X1 MEM_stage_inst_dmem_U9863 ( .A1(MEM_stage_inst_dmem_ram_136), .A2(MEM_stage_inst_dmem_n13486), .ZN(MEM_stage_inst_dmem_n13471) );
NAND2_X1 MEM_stage_inst_dmem_U9862 ( .A1(MEM_stage_inst_dmem_n13469), .A2(MEM_stage_inst_dmem_n13468), .ZN(MEM_stage_inst_dmem_n12484) );
NAND2_X1 MEM_stage_inst_dmem_U9861 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n13487), .ZN(MEM_stage_inst_dmem_n13468) );
NAND2_X1 MEM_stage_inst_dmem_U9860 ( .A1(MEM_stage_inst_dmem_ram_137), .A2(MEM_stage_inst_dmem_n13486), .ZN(MEM_stage_inst_dmem_n13469) );
NAND2_X1 MEM_stage_inst_dmem_U9859 ( .A1(MEM_stage_inst_dmem_n13467), .A2(MEM_stage_inst_dmem_n13466), .ZN(MEM_stage_inst_dmem_n12485) );
NAND2_X1 MEM_stage_inst_dmem_U9858 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n13487), .ZN(MEM_stage_inst_dmem_n13466) );
NAND2_X1 MEM_stage_inst_dmem_U9857 ( .A1(MEM_stage_inst_dmem_ram_138), .A2(MEM_stage_inst_dmem_n13486), .ZN(MEM_stage_inst_dmem_n13467) );
NAND2_X1 MEM_stage_inst_dmem_U9856 ( .A1(MEM_stage_inst_dmem_n13465), .A2(MEM_stage_inst_dmem_n13464), .ZN(MEM_stage_inst_dmem_n12486) );
NAND2_X1 MEM_stage_inst_dmem_U9855 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n13487), .ZN(MEM_stage_inst_dmem_n13464) );
NAND2_X1 MEM_stage_inst_dmem_U9854 ( .A1(MEM_stage_inst_dmem_ram_139), .A2(MEM_stage_inst_dmem_n13486), .ZN(MEM_stage_inst_dmem_n13465) );
NAND2_X1 MEM_stage_inst_dmem_U9853 ( .A1(MEM_stage_inst_dmem_n13463), .A2(MEM_stage_inst_dmem_n13462), .ZN(MEM_stage_inst_dmem_n12487) );
NAND2_X1 MEM_stage_inst_dmem_U9852 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n13487), .ZN(MEM_stage_inst_dmem_n13462) );
NAND2_X1 MEM_stage_inst_dmem_U9851 ( .A1(MEM_stage_inst_dmem_ram_140), .A2(MEM_stage_inst_dmem_n13486), .ZN(MEM_stage_inst_dmem_n13463) );
NAND2_X1 MEM_stage_inst_dmem_U9850 ( .A1(MEM_stage_inst_dmem_n13461), .A2(MEM_stage_inst_dmem_n13460), .ZN(MEM_stage_inst_dmem_n12488) );
NAND2_X1 MEM_stage_inst_dmem_U9849 ( .A1(MEM_stage_inst_dmem_n116), .A2(MEM_stage_inst_dmem_n13487), .ZN(MEM_stage_inst_dmem_n13460) );
NAND2_X1 MEM_stage_inst_dmem_U9848 ( .A1(MEM_stage_inst_dmem_ram_141), .A2(MEM_stage_inst_dmem_n13486), .ZN(MEM_stage_inst_dmem_n13461) );
NAND2_X1 MEM_stage_inst_dmem_U9847 ( .A1(MEM_stage_inst_dmem_n13459), .A2(MEM_stage_inst_dmem_n13458), .ZN(MEM_stage_inst_dmem_n12489) );
NAND2_X1 MEM_stage_inst_dmem_U9846 ( .A1(MEM_stage_inst_dmem_n14696), .A2(MEM_stage_inst_dmem_n13487), .ZN(MEM_stage_inst_dmem_n13458) );
NAND2_X1 MEM_stage_inst_dmem_U9845 ( .A1(MEM_stage_inst_dmem_ram_142), .A2(MEM_stage_inst_dmem_n13486), .ZN(MEM_stage_inst_dmem_n13459) );
NAND2_X1 MEM_stage_inst_dmem_U9844 ( .A1(MEM_stage_inst_dmem_n13457), .A2(MEM_stage_inst_dmem_n13456), .ZN(MEM_stage_inst_dmem_n12490) );
NAND2_X1 MEM_stage_inst_dmem_U9843 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n13487), .ZN(MEM_stage_inst_dmem_n13456) );
INV_X1 MEM_stage_inst_dmem_U9842 ( .A(MEM_stage_inst_dmem_n13486), .ZN(MEM_stage_inst_dmem_n13487) );
NAND2_X1 MEM_stage_inst_dmem_U9841 ( .A1(MEM_stage_inst_dmem_ram_143), .A2(MEM_stage_inst_dmem_n13486), .ZN(MEM_stage_inst_dmem_n13457) );
NAND2_X1 MEM_stage_inst_dmem_U9840 ( .A1(MEM_stage_inst_dmem_n21179), .A2(MEM_stage_inst_dmem_n13728), .ZN(MEM_stage_inst_dmem_n13486) );
NAND2_X1 MEM_stage_inst_dmem_U9839 ( .A1(MEM_stage_inst_dmem_n13455), .A2(MEM_stage_inst_dmem_n13454), .ZN(MEM_stage_inst_dmem_n12491) );
NAND2_X1 MEM_stage_inst_dmem_U9838 ( .A1(EX_pipeline_reg_out_5), .A2(MEM_stage_inst_dmem_n13453), .ZN(MEM_stage_inst_dmem_n13454) );
NAND2_X1 MEM_stage_inst_dmem_U9837 ( .A1(MEM_stage_inst_dmem_ram_144), .A2(MEM_stage_inst_dmem_n13452), .ZN(MEM_stage_inst_dmem_n13455) );
NAND2_X1 MEM_stage_inst_dmem_U9836 ( .A1(MEM_stage_inst_dmem_n13451), .A2(MEM_stage_inst_dmem_n13450), .ZN(MEM_stage_inst_dmem_n12492) );
NAND2_X1 MEM_stage_inst_dmem_U9835 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n13453), .ZN(MEM_stage_inst_dmem_n13450) );
NAND2_X1 MEM_stage_inst_dmem_U9834 ( .A1(MEM_stage_inst_dmem_ram_145), .A2(MEM_stage_inst_dmem_n13452), .ZN(MEM_stage_inst_dmem_n13451) );
NAND2_X1 MEM_stage_inst_dmem_U9833 ( .A1(MEM_stage_inst_dmem_n13449), .A2(MEM_stage_inst_dmem_n13448), .ZN(MEM_stage_inst_dmem_n12493) );
NAND2_X1 MEM_stage_inst_dmem_U9832 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n13453), .ZN(MEM_stage_inst_dmem_n13448) );
NAND2_X1 MEM_stage_inst_dmem_U9831 ( .A1(MEM_stage_inst_dmem_ram_146), .A2(MEM_stage_inst_dmem_n13452), .ZN(MEM_stage_inst_dmem_n13449) );
NAND2_X1 MEM_stage_inst_dmem_U9830 ( .A1(MEM_stage_inst_dmem_n13447), .A2(MEM_stage_inst_dmem_n13446), .ZN(MEM_stage_inst_dmem_n12494) );
NAND2_X1 MEM_stage_inst_dmem_U9829 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n13453), .ZN(MEM_stage_inst_dmem_n13446) );
NAND2_X1 MEM_stage_inst_dmem_U9828 ( .A1(MEM_stage_inst_dmem_ram_147), .A2(MEM_stage_inst_dmem_n13452), .ZN(MEM_stage_inst_dmem_n13447) );
NAND2_X1 MEM_stage_inst_dmem_U9827 ( .A1(MEM_stage_inst_dmem_n13445), .A2(MEM_stage_inst_dmem_n13444), .ZN(MEM_stage_inst_dmem_n12495) );
NAND2_X1 MEM_stage_inst_dmem_U9826 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n13453), .ZN(MEM_stage_inst_dmem_n13444) );
NAND2_X1 MEM_stage_inst_dmem_U9825 ( .A1(MEM_stage_inst_dmem_ram_148), .A2(MEM_stage_inst_dmem_n13452), .ZN(MEM_stage_inst_dmem_n13445) );
NAND2_X1 MEM_stage_inst_dmem_U9824 ( .A1(MEM_stage_inst_dmem_n13443), .A2(MEM_stage_inst_dmem_n13442), .ZN(MEM_stage_inst_dmem_n12496) );
NAND2_X1 MEM_stage_inst_dmem_U9823 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n13453), .ZN(MEM_stage_inst_dmem_n13442) );
NAND2_X1 MEM_stage_inst_dmem_U9822 ( .A1(MEM_stage_inst_dmem_ram_149), .A2(MEM_stage_inst_dmem_n13452), .ZN(MEM_stage_inst_dmem_n13443) );
NAND2_X1 MEM_stage_inst_dmem_U9821 ( .A1(MEM_stage_inst_dmem_n13441), .A2(MEM_stage_inst_dmem_n13440), .ZN(MEM_stage_inst_dmem_n12497) );
NAND2_X1 MEM_stage_inst_dmem_U9820 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n13453), .ZN(MEM_stage_inst_dmem_n13440) );
NAND2_X1 MEM_stage_inst_dmem_U9819 ( .A1(MEM_stage_inst_dmem_ram_150), .A2(MEM_stage_inst_dmem_n13452), .ZN(MEM_stage_inst_dmem_n13441) );
NAND2_X1 MEM_stage_inst_dmem_U9818 ( .A1(MEM_stage_inst_dmem_n13439), .A2(MEM_stage_inst_dmem_n13438), .ZN(MEM_stage_inst_dmem_n12498) );
NAND2_X1 MEM_stage_inst_dmem_U9817 ( .A1(MEM_stage_inst_dmem_n13886), .A2(MEM_stage_inst_dmem_n13453), .ZN(MEM_stage_inst_dmem_n13438) );
NAND2_X1 MEM_stage_inst_dmem_U9816 ( .A1(MEM_stage_inst_dmem_ram_151), .A2(MEM_stage_inst_dmem_n13452), .ZN(MEM_stage_inst_dmem_n13439) );
NAND2_X1 MEM_stage_inst_dmem_U9815 ( .A1(MEM_stage_inst_dmem_n13437), .A2(MEM_stage_inst_dmem_n13436), .ZN(MEM_stage_inst_dmem_n12499) );
NAND2_X1 MEM_stage_inst_dmem_U9814 ( .A1(MEM_stage_inst_dmem_n13883), .A2(MEM_stage_inst_dmem_n13453), .ZN(MEM_stage_inst_dmem_n13436) );
NAND2_X1 MEM_stage_inst_dmem_U9813 ( .A1(MEM_stage_inst_dmem_ram_152), .A2(MEM_stage_inst_dmem_n13452), .ZN(MEM_stage_inst_dmem_n13437) );
NAND2_X1 MEM_stage_inst_dmem_U9812 ( .A1(MEM_stage_inst_dmem_n13435), .A2(MEM_stage_inst_dmem_n13434), .ZN(MEM_stage_inst_dmem_n12500) );
NAND2_X1 MEM_stage_inst_dmem_U9811 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n13453), .ZN(MEM_stage_inst_dmem_n13434) );
NAND2_X1 MEM_stage_inst_dmem_U9810 ( .A1(MEM_stage_inst_dmem_ram_153), .A2(MEM_stage_inst_dmem_n13452), .ZN(MEM_stage_inst_dmem_n13435) );
NAND2_X1 MEM_stage_inst_dmem_U9809 ( .A1(MEM_stage_inst_dmem_n13433), .A2(MEM_stage_inst_dmem_n13432), .ZN(MEM_stage_inst_dmem_n12501) );
NAND2_X1 MEM_stage_inst_dmem_U9808 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n13453), .ZN(MEM_stage_inst_dmem_n13432) );
NAND2_X1 MEM_stage_inst_dmem_U9807 ( .A1(MEM_stage_inst_dmem_ram_154), .A2(MEM_stage_inst_dmem_n13452), .ZN(MEM_stage_inst_dmem_n13433) );
NAND2_X1 MEM_stage_inst_dmem_U9806 ( .A1(MEM_stage_inst_dmem_n13431), .A2(MEM_stage_inst_dmem_n13430), .ZN(MEM_stage_inst_dmem_n12502) );
NAND2_X1 MEM_stage_inst_dmem_U9805 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n13453), .ZN(MEM_stage_inst_dmem_n13430) );
NAND2_X1 MEM_stage_inst_dmem_U9804 ( .A1(MEM_stage_inst_dmem_ram_155), .A2(MEM_stage_inst_dmem_n13452), .ZN(MEM_stage_inst_dmem_n13431) );
NAND2_X1 MEM_stage_inst_dmem_U9803 ( .A1(MEM_stage_inst_dmem_n13429), .A2(MEM_stage_inst_dmem_n13428), .ZN(MEM_stage_inst_dmem_n12503) );
NAND2_X1 MEM_stage_inst_dmem_U9802 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n13453), .ZN(MEM_stage_inst_dmem_n13428) );
NAND2_X1 MEM_stage_inst_dmem_U9801 ( .A1(MEM_stage_inst_dmem_ram_156), .A2(MEM_stage_inst_dmem_n13452), .ZN(MEM_stage_inst_dmem_n13429) );
NAND2_X1 MEM_stage_inst_dmem_U9800 ( .A1(MEM_stage_inst_dmem_n13427), .A2(MEM_stage_inst_dmem_n13426), .ZN(MEM_stage_inst_dmem_n12504) );
NAND2_X1 MEM_stage_inst_dmem_U9799 ( .A1(EX_pipeline_reg_out_18), .A2(MEM_stage_inst_dmem_n13453), .ZN(MEM_stage_inst_dmem_n13426) );
NAND2_X1 MEM_stage_inst_dmem_U9798 ( .A1(MEM_stage_inst_dmem_ram_157), .A2(MEM_stage_inst_dmem_n13452), .ZN(MEM_stage_inst_dmem_n13427) );
NAND2_X1 MEM_stage_inst_dmem_U9797 ( .A1(MEM_stage_inst_dmem_n13425), .A2(MEM_stage_inst_dmem_n13424), .ZN(MEM_stage_inst_dmem_n12505) );
NAND2_X1 MEM_stage_inst_dmem_U9796 ( .A1(EX_pipeline_reg_out_19), .A2(MEM_stage_inst_dmem_n13453), .ZN(MEM_stage_inst_dmem_n13424) );
NAND2_X1 MEM_stage_inst_dmem_U9795 ( .A1(MEM_stage_inst_dmem_ram_158), .A2(MEM_stage_inst_dmem_n13452), .ZN(MEM_stage_inst_dmem_n13425) );
NAND2_X1 MEM_stage_inst_dmem_U9794 ( .A1(MEM_stage_inst_dmem_n13423), .A2(MEM_stage_inst_dmem_n13422), .ZN(MEM_stage_inst_dmem_n12506) );
NAND2_X1 MEM_stage_inst_dmem_U9793 ( .A1(EX_pipeline_reg_out_20), .A2(MEM_stage_inst_dmem_n13453), .ZN(MEM_stage_inst_dmem_n13422) );
INV_X1 MEM_stage_inst_dmem_U9792 ( .A(MEM_stage_inst_dmem_n13452), .ZN(MEM_stage_inst_dmem_n13453) );
NAND2_X1 MEM_stage_inst_dmem_U9791 ( .A1(MEM_stage_inst_dmem_ram_159), .A2(MEM_stage_inst_dmem_n13452), .ZN(MEM_stage_inst_dmem_n13423) );
NAND2_X1 MEM_stage_inst_dmem_U9790 ( .A1(MEM_stage_inst_dmem_n21144), .A2(MEM_stage_inst_dmem_n13728), .ZN(MEM_stage_inst_dmem_n13452) );
NAND2_X1 MEM_stage_inst_dmem_U9789 ( .A1(MEM_stage_inst_dmem_n13421), .A2(MEM_stage_inst_dmem_n13420), .ZN(MEM_stage_inst_dmem_n12507) );
NAND2_X1 MEM_stage_inst_dmem_U9788 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n13419), .ZN(MEM_stage_inst_dmem_n13420) );
NAND2_X1 MEM_stage_inst_dmem_U9787 ( .A1(MEM_stage_inst_dmem_ram_160), .A2(MEM_stage_inst_dmem_n13418), .ZN(MEM_stage_inst_dmem_n13421) );
NAND2_X1 MEM_stage_inst_dmem_U9786 ( .A1(MEM_stage_inst_dmem_n13417), .A2(MEM_stage_inst_dmem_n13416), .ZN(MEM_stage_inst_dmem_n12508) );
NAND2_X1 MEM_stage_inst_dmem_U9785 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n13419), .ZN(MEM_stage_inst_dmem_n13416) );
NAND2_X1 MEM_stage_inst_dmem_U9784 ( .A1(MEM_stage_inst_dmem_ram_161), .A2(MEM_stage_inst_dmem_n13418), .ZN(MEM_stage_inst_dmem_n13417) );
NAND2_X1 MEM_stage_inst_dmem_U9783 ( .A1(MEM_stage_inst_dmem_n13415), .A2(MEM_stage_inst_dmem_n13414), .ZN(MEM_stage_inst_dmem_n12509) );
NAND2_X1 MEM_stage_inst_dmem_U9782 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n13419), .ZN(MEM_stage_inst_dmem_n13414) );
NAND2_X1 MEM_stage_inst_dmem_U9781 ( .A1(MEM_stage_inst_dmem_ram_162), .A2(MEM_stage_inst_dmem_n13418), .ZN(MEM_stage_inst_dmem_n13415) );
NAND2_X1 MEM_stage_inst_dmem_U9780 ( .A1(MEM_stage_inst_dmem_n13413), .A2(MEM_stage_inst_dmem_n13412), .ZN(MEM_stage_inst_dmem_n12510) );
NAND2_X1 MEM_stage_inst_dmem_U9779 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n13419), .ZN(MEM_stage_inst_dmem_n13412) );
NAND2_X1 MEM_stage_inst_dmem_U9778 ( .A1(MEM_stage_inst_dmem_ram_163), .A2(MEM_stage_inst_dmem_n13418), .ZN(MEM_stage_inst_dmem_n13413) );
NAND2_X1 MEM_stage_inst_dmem_U9777 ( .A1(MEM_stage_inst_dmem_n13411), .A2(MEM_stage_inst_dmem_n13410), .ZN(MEM_stage_inst_dmem_n12511) );
NAND2_X1 MEM_stage_inst_dmem_U9776 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n13419), .ZN(MEM_stage_inst_dmem_n13410) );
NAND2_X1 MEM_stage_inst_dmem_U9775 ( .A1(MEM_stage_inst_dmem_ram_164), .A2(MEM_stage_inst_dmem_n13418), .ZN(MEM_stage_inst_dmem_n13411) );
NAND2_X1 MEM_stage_inst_dmem_U9774 ( .A1(MEM_stage_inst_dmem_n13409), .A2(MEM_stage_inst_dmem_n13408), .ZN(MEM_stage_inst_dmem_n12512) );
NAND2_X1 MEM_stage_inst_dmem_U9773 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n13419), .ZN(MEM_stage_inst_dmem_n13408) );
NAND2_X1 MEM_stage_inst_dmem_U9772 ( .A1(MEM_stage_inst_dmem_ram_165), .A2(MEM_stage_inst_dmem_n13418), .ZN(MEM_stage_inst_dmem_n13409) );
NAND2_X1 MEM_stage_inst_dmem_U9771 ( .A1(MEM_stage_inst_dmem_n13407), .A2(MEM_stage_inst_dmem_n13406), .ZN(MEM_stage_inst_dmem_n12513) );
NAND2_X1 MEM_stage_inst_dmem_U9770 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n13419), .ZN(MEM_stage_inst_dmem_n13406) );
NAND2_X1 MEM_stage_inst_dmem_U9769 ( .A1(MEM_stage_inst_dmem_ram_166), .A2(MEM_stage_inst_dmem_n13418), .ZN(MEM_stage_inst_dmem_n13407) );
NAND2_X1 MEM_stage_inst_dmem_U9768 ( .A1(MEM_stage_inst_dmem_n13405), .A2(MEM_stage_inst_dmem_n13404), .ZN(MEM_stage_inst_dmem_n12514) );
NAND2_X1 MEM_stage_inst_dmem_U9767 ( .A1(MEM_stage_inst_dmem_n18), .A2(MEM_stage_inst_dmem_n13419), .ZN(MEM_stage_inst_dmem_n13404) );
NAND2_X1 MEM_stage_inst_dmem_U9766 ( .A1(MEM_stage_inst_dmem_ram_167), .A2(MEM_stage_inst_dmem_n13418), .ZN(MEM_stage_inst_dmem_n13405) );
NAND2_X1 MEM_stage_inst_dmem_U9765 ( .A1(MEM_stage_inst_dmem_n13403), .A2(MEM_stage_inst_dmem_n13402), .ZN(MEM_stage_inst_dmem_n12515) );
NAND2_X1 MEM_stage_inst_dmem_U9764 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n13419), .ZN(MEM_stage_inst_dmem_n13402) );
NAND2_X1 MEM_stage_inst_dmem_U9763 ( .A1(MEM_stage_inst_dmem_ram_168), .A2(MEM_stage_inst_dmem_n13418), .ZN(MEM_stage_inst_dmem_n13403) );
NAND2_X1 MEM_stage_inst_dmem_U9762 ( .A1(MEM_stage_inst_dmem_n13401), .A2(MEM_stage_inst_dmem_n13400), .ZN(MEM_stage_inst_dmem_n12516) );
NAND2_X1 MEM_stage_inst_dmem_U9761 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n13419), .ZN(MEM_stage_inst_dmem_n13400) );
NAND2_X1 MEM_stage_inst_dmem_U9760 ( .A1(MEM_stage_inst_dmem_ram_169), .A2(MEM_stage_inst_dmem_n13418), .ZN(MEM_stage_inst_dmem_n13401) );
NAND2_X1 MEM_stage_inst_dmem_U9759 ( .A1(MEM_stage_inst_dmem_n13399), .A2(MEM_stage_inst_dmem_n13398), .ZN(MEM_stage_inst_dmem_n12517) );
NAND2_X1 MEM_stage_inst_dmem_U9758 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n13419), .ZN(MEM_stage_inst_dmem_n13398) );
NAND2_X1 MEM_stage_inst_dmem_U9757 ( .A1(MEM_stage_inst_dmem_ram_170), .A2(MEM_stage_inst_dmem_n13418), .ZN(MEM_stage_inst_dmem_n13399) );
NAND2_X1 MEM_stage_inst_dmem_U9756 ( .A1(MEM_stage_inst_dmem_n13397), .A2(MEM_stage_inst_dmem_n13396), .ZN(MEM_stage_inst_dmem_n12518) );
NAND2_X1 MEM_stage_inst_dmem_U9755 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n13419), .ZN(MEM_stage_inst_dmem_n13396) );
NAND2_X1 MEM_stage_inst_dmem_U9754 ( .A1(MEM_stage_inst_dmem_ram_171), .A2(MEM_stage_inst_dmem_n13418), .ZN(MEM_stage_inst_dmem_n13397) );
NAND2_X1 MEM_stage_inst_dmem_U9753 ( .A1(MEM_stage_inst_dmem_n13395), .A2(MEM_stage_inst_dmem_n13394), .ZN(MEM_stage_inst_dmem_n12519) );
NAND2_X1 MEM_stage_inst_dmem_U9752 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n13419), .ZN(MEM_stage_inst_dmem_n13394) );
NAND2_X1 MEM_stage_inst_dmem_U9751 ( .A1(MEM_stage_inst_dmem_ram_172), .A2(MEM_stage_inst_dmem_n13418), .ZN(MEM_stage_inst_dmem_n13395) );
NAND2_X1 MEM_stage_inst_dmem_U9750 ( .A1(MEM_stage_inst_dmem_n13393), .A2(MEM_stage_inst_dmem_n13392), .ZN(MEM_stage_inst_dmem_n12520) );
NAND2_X1 MEM_stage_inst_dmem_U9749 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n13419), .ZN(MEM_stage_inst_dmem_n13392) );
NAND2_X1 MEM_stage_inst_dmem_U9748 ( .A1(MEM_stage_inst_dmem_ram_173), .A2(MEM_stage_inst_dmem_n13418), .ZN(MEM_stage_inst_dmem_n13393) );
NAND2_X1 MEM_stage_inst_dmem_U9747 ( .A1(MEM_stage_inst_dmem_n13391), .A2(MEM_stage_inst_dmem_n13390), .ZN(MEM_stage_inst_dmem_n12521) );
NAND2_X1 MEM_stage_inst_dmem_U9746 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n13419), .ZN(MEM_stage_inst_dmem_n13390) );
NAND2_X1 MEM_stage_inst_dmem_U9745 ( .A1(MEM_stage_inst_dmem_ram_174), .A2(MEM_stage_inst_dmem_n13418), .ZN(MEM_stage_inst_dmem_n13391) );
NAND2_X1 MEM_stage_inst_dmem_U9744 ( .A1(MEM_stage_inst_dmem_n13389), .A2(MEM_stage_inst_dmem_n13388), .ZN(MEM_stage_inst_dmem_n12522) );
NAND2_X1 MEM_stage_inst_dmem_U9743 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n13419), .ZN(MEM_stage_inst_dmem_n13388) );
NAND2_X1 MEM_stage_inst_dmem_U9742 ( .A1(MEM_stage_inst_dmem_ram_175), .A2(MEM_stage_inst_dmem_n13418), .ZN(MEM_stage_inst_dmem_n13389) );
NAND2_X1 MEM_stage_inst_dmem_U9741 ( .A1(MEM_stage_inst_dmem_n21109), .A2(MEM_stage_inst_dmem_n13728), .ZN(MEM_stage_inst_dmem_n13418) );
NAND2_X1 MEM_stage_inst_dmem_U9740 ( .A1(MEM_stage_inst_dmem_n13387), .A2(MEM_stage_inst_dmem_n13386), .ZN(MEM_stage_inst_dmem_n12523) );
NAND2_X1 MEM_stage_inst_dmem_U9739 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n13385), .ZN(MEM_stage_inst_dmem_n13386) );
NAND2_X1 MEM_stage_inst_dmem_U9738 ( .A1(MEM_stage_inst_dmem_ram_176), .A2(MEM_stage_inst_dmem_n13384), .ZN(MEM_stage_inst_dmem_n13387) );
NAND2_X1 MEM_stage_inst_dmem_U9737 ( .A1(MEM_stage_inst_dmem_n13383), .A2(MEM_stage_inst_dmem_n13382), .ZN(MEM_stage_inst_dmem_n12524) );
NAND2_X1 MEM_stage_inst_dmem_U9736 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n13385), .ZN(MEM_stage_inst_dmem_n13382) );
NAND2_X1 MEM_stage_inst_dmem_U9735 ( .A1(MEM_stage_inst_dmem_ram_177), .A2(MEM_stage_inst_dmem_n13384), .ZN(MEM_stage_inst_dmem_n13383) );
NAND2_X1 MEM_stage_inst_dmem_U9734 ( .A1(MEM_stage_inst_dmem_n13381), .A2(MEM_stage_inst_dmem_n13380), .ZN(MEM_stage_inst_dmem_n12525) );
NAND2_X1 MEM_stage_inst_dmem_U9733 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n13385), .ZN(MEM_stage_inst_dmem_n13380) );
NAND2_X1 MEM_stage_inst_dmem_U9732 ( .A1(MEM_stage_inst_dmem_ram_178), .A2(MEM_stage_inst_dmem_n13384), .ZN(MEM_stage_inst_dmem_n13381) );
NAND2_X1 MEM_stage_inst_dmem_U9731 ( .A1(MEM_stage_inst_dmem_n13379), .A2(MEM_stage_inst_dmem_n13378), .ZN(MEM_stage_inst_dmem_n12526) );
NAND2_X1 MEM_stage_inst_dmem_U9730 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n13385), .ZN(MEM_stage_inst_dmem_n13378) );
NAND2_X1 MEM_stage_inst_dmem_U9729 ( .A1(MEM_stage_inst_dmem_ram_179), .A2(MEM_stage_inst_dmem_n13384), .ZN(MEM_stage_inst_dmem_n13379) );
NAND2_X1 MEM_stage_inst_dmem_U9728 ( .A1(MEM_stage_inst_dmem_n13377), .A2(MEM_stage_inst_dmem_n13376), .ZN(MEM_stage_inst_dmem_n12527) );
NAND2_X1 MEM_stage_inst_dmem_U9727 ( .A1(MEM_stage_inst_dmem_n16368), .A2(MEM_stage_inst_dmem_n13385), .ZN(MEM_stage_inst_dmem_n13376) );
NAND2_X1 MEM_stage_inst_dmem_U9726 ( .A1(MEM_stage_inst_dmem_ram_180), .A2(MEM_stage_inst_dmem_n13384), .ZN(MEM_stage_inst_dmem_n13377) );
NAND2_X1 MEM_stage_inst_dmem_U9725 ( .A1(MEM_stage_inst_dmem_n13375), .A2(MEM_stage_inst_dmem_n13374), .ZN(MEM_stage_inst_dmem_n12528) );
NAND2_X1 MEM_stage_inst_dmem_U9724 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n13385), .ZN(MEM_stage_inst_dmem_n13374) );
NAND2_X1 MEM_stage_inst_dmem_U9723 ( .A1(MEM_stage_inst_dmem_ram_181), .A2(MEM_stage_inst_dmem_n13384), .ZN(MEM_stage_inst_dmem_n13375) );
NAND2_X1 MEM_stage_inst_dmem_U9722 ( .A1(MEM_stage_inst_dmem_n13373), .A2(MEM_stage_inst_dmem_n13372), .ZN(MEM_stage_inst_dmem_n12529) );
NAND2_X1 MEM_stage_inst_dmem_U9721 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n13385), .ZN(MEM_stage_inst_dmem_n13372) );
NAND2_X1 MEM_stage_inst_dmem_U9720 ( .A1(MEM_stage_inst_dmem_ram_182), .A2(MEM_stage_inst_dmem_n13384), .ZN(MEM_stage_inst_dmem_n13373) );
NAND2_X1 MEM_stage_inst_dmem_U9719 ( .A1(MEM_stage_inst_dmem_n13371), .A2(MEM_stage_inst_dmem_n13370), .ZN(MEM_stage_inst_dmem_n12530) );
NAND2_X1 MEM_stage_inst_dmem_U9718 ( .A1(MEM_stage_inst_dmem_n13886), .A2(MEM_stage_inst_dmem_n13385), .ZN(MEM_stage_inst_dmem_n13370) );
NAND2_X1 MEM_stage_inst_dmem_U9717 ( .A1(MEM_stage_inst_dmem_ram_183), .A2(MEM_stage_inst_dmem_n13384), .ZN(MEM_stage_inst_dmem_n13371) );
NAND2_X1 MEM_stage_inst_dmem_U9716 ( .A1(MEM_stage_inst_dmem_n13369), .A2(MEM_stage_inst_dmem_n13368), .ZN(MEM_stage_inst_dmem_n12531) );
NAND2_X1 MEM_stage_inst_dmem_U9715 ( .A1(MEM_stage_inst_dmem_n13883), .A2(MEM_stage_inst_dmem_n13385), .ZN(MEM_stage_inst_dmem_n13368) );
NAND2_X1 MEM_stage_inst_dmem_U9714 ( .A1(MEM_stage_inst_dmem_ram_184), .A2(MEM_stage_inst_dmem_n13384), .ZN(MEM_stage_inst_dmem_n13369) );
NAND2_X1 MEM_stage_inst_dmem_U9713 ( .A1(MEM_stage_inst_dmem_n13367), .A2(MEM_stage_inst_dmem_n13366), .ZN(MEM_stage_inst_dmem_n12532) );
NAND2_X1 MEM_stage_inst_dmem_U9712 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n13385), .ZN(MEM_stage_inst_dmem_n13366) );
NAND2_X1 MEM_stage_inst_dmem_U9711 ( .A1(MEM_stage_inst_dmem_ram_185), .A2(MEM_stage_inst_dmem_n13384), .ZN(MEM_stage_inst_dmem_n13367) );
NAND2_X1 MEM_stage_inst_dmem_U9710 ( .A1(MEM_stage_inst_dmem_n13365), .A2(MEM_stage_inst_dmem_n13364), .ZN(MEM_stage_inst_dmem_n12533) );
NAND2_X1 MEM_stage_inst_dmem_U9709 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n13385), .ZN(MEM_stage_inst_dmem_n13364) );
NAND2_X1 MEM_stage_inst_dmem_U9708 ( .A1(MEM_stage_inst_dmem_ram_186), .A2(MEM_stage_inst_dmem_n13384), .ZN(MEM_stage_inst_dmem_n13365) );
NAND2_X1 MEM_stage_inst_dmem_U9707 ( .A1(MEM_stage_inst_dmem_n13363), .A2(MEM_stage_inst_dmem_n13362), .ZN(MEM_stage_inst_dmem_n12534) );
NAND2_X1 MEM_stage_inst_dmem_U9706 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n13385), .ZN(MEM_stage_inst_dmem_n13362) );
NAND2_X1 MEM_stage_inst_dmem_U9705 ( .A1(MEM_stage_inst_dmem_ram_187), .A2(MEM_stage_inst_dmem_n13384), .ZN(MEM_stage_inst_dmem_n13363) );
NAND2_X1 MEM_stage_inst_dmem_U9704 ( .A1(MEM_stage_inst_dmem_n13361), .A2(MEM_stage_inst_dmem_n13360), .ZN(MEM_stage_inst_dmem_n12535) );
NAND2_X1 MEM_stage_inst_dmem_U9703 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n13385), .ZN(MEM_stage_inst_dmem_n13360) );
NAND2_X1 MEM_stage_inst_dmem_U9702 ( .A1(MEM_stage_inst_dmem_ram_188), .A2(MEM_stage_inst_dmem_n13384), .ZN(MEM_stage_inst_dmem_n13361) );
NAND2_X1 MEM_stage_inst_dmem_U9701 ( .A1(MEM_stage_inst_dmem_n13359), .A2(MEM_stage_inst_dmem_n13358), .ZN(MEM_stage_inst_dmem_n12536) );
NAND2_X1 MEM_stage_inst_dmem_U9700 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n13385), .ZN(MEM_stage_inst_dmem_n13358) );
NAND2_X1 MEM_stage_inst_dmem_U9699 ( .A1(MEM_stage_inst_dmem_ram_189), .A2(MEM_stage_inst_dmem_n13384), .ZN(MEM_stage_inst_dmem_n13359) );
NAND2_X1 MEM_stage_inst_dmem_U9698 ( .A1(MEM_stage_inst_dmem_n13357), .A2(MEM_stage_inst_dmem_n13356), .ZN(MEM_stage_inst_dmem_n12537) );
NAND2_X1 MEM_stage_inst_dmem_U9697 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n13385), .ZN(MEM_stage_inst_dmem_n13356) );
NAND2_X1 MEM_stage_inst_dmem_U9696 ( .A1(MEM_stage_inst_dmem_ram_190), .A2(MEM_stage_inst_dmem_n13384), .ZN(MEM_stage_inst_dmem_n13357) );
NAND2_X1 MEM_stage_inst_dmem_U9695 ( .A1(MEM_stage_inst_dmem_n13355), .A2(MEM_stage_inst_dmem_n13354), .ZN(MEM_stage_inst_dmem_n12538) );
NAND2_X1 MEM_stage_inst_dmem_U9694 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n13385), .ZN(MEM_stage_inst_dmem_n13354) );
INV_X1 MEM_stage_inst_dmem_U9693 ( .A(MEM_stage_inst_dmem_n13384), .ZN(MEM_stage_inst_dmem_n13385) );
NAND2_X1 MEM_stage_inst_dmem_U9692 ( .A1(MEM_stage_inst_dmem_ram_191), .A2(MEM_stage_inst_dmem_n13384), .ZN(MEM_stage_inst_dmem_n13355) );
NAND2_X1 MEM_stage_inst_dmem_U9691 ( .A1(MEM_stage_inst_dmem_n21074), .A2(MEM_stage_inst_dmem_n13728), .ZN(MEM_stage_inst_dmem_n13384) );
NAND2_X1 MEM_stage_inst_dmem_U9690 ( .A1(MEM_stage_inst_dmem_n13353), .A2(MEM_stage_inst_dmem_n13352), .ZN(MEM_stage_inst_dmem_n12539) );
NAND2_X1 MEM_stage_inst_dmem_U9689 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n13351), .ZN(MEM_stage_inst_dmem_n13352) );
NAND2_X1 MEM_stage_inst_dmem_U9688 ( .A1(MEM_stage_inst_dmem_ram_192), .A2(MEM_stage_inst_dmem_n13350), .ZN(MEM_stage_inst_dmem_n13353) );
NAND2_X1 MEM_stage_inst_dmem_U9687 ( .A1(MEM_stage_inst_dmem_n13349), .A2(MEM_stage_inst_dmem_n13348), .ZN(MEM_stage_inst_dmem_n12540) );
NAND2_X1 MEM_stage_inst_dmem_U9686 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n13351), .ZN(MEM_stage_inst_dmem_n13348) );
NAND2_X1 MEM_stage_inst_dmem_U9685 ( .A1(MEM_stage_inst_dmem_ram_193), .A2(MEM_stage_inst_dmem_n13350), .ZN(MEM_stage_inst_dmem_n13349) );
NAND2_X1 MEM_stage_inst_dmem_U9684 ( .A1(MEM_stage_inst_dmem_n13347), .A2(MEM_stage_inst_dmem_n13346), .ZN(MEM_stage_inst_dmem_n12541) );
NAND2_X1 MEM_stage_inst_dmem_U9683 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n13351), .ZN(MEM_stage_inst_dmem_n13346) );
NAND2_X1 MEM_stage_inst_dmem_U9682 ( .A1(MEM_stage_inst_dmem_ram_194), .A2(MEM_stage_inst_dmem_n13350), .ZN(MEM_stage_inst_dmem_n13347) );
NAND2_X1 MEM_stage_inst_dmem_U9681 ( .A1(MEM_stage_inst_dmem_n13345), .A2(MEM_stage_inst_dmem_n13344), .ZN(MEM_stage_inst_dmem_n12542) );
NAND2_X1 MEM_stage_inst_dmem_U9680 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n13351), .ZN(MEM_stage_inst_dmem_n13344) );
NAND2_X1 MEM_stage_inst_dmem_U9679 ( .A1(MEM_stage_inst_dmem_ram_195), .A2(MEM_stage_inst_dmem_n13350), .ZN(MEM_stage_inst_dmem_n13345) );
NAND2_X1 MEM_stage_inst_dmem_U9678 ( .A1(MEM_stage_inst_dmem_n13343), .A2(MEM_stage_inst_dmem_n13342), .ZN(MEM_stage_inst_dmem_n12543) );
NAND2_X1 MEM_stage_inst_dmem_U9677 ( .A1(MEM_stage_inst_dmem_n16784), .A2(MEM_stage_inst_dmem_n13351), .ZN(MEM_stage_inst_dmem_n13342) );
NAND2_X1 MEM_stage_inst_dmem_U9676 ( .A1(MEM_stage_inst_dmem_ram_196), .A2(MEM_stage_inst_dmem_n13350), .ZN(MEM_stage_inst_dmem_n13343) );
NAND2_X1 MEM_stage_inst_dmem_U9675 ( .A1(MEM_stage_inst_dmem_n13341), .A2(MEM_stage_inst_dmem_n13340), .ZN(MEM_stage_inst_dmem_n12544) );
NAND2_X1 MEM_stage_inst_dmem_U9674 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n13351), .ZN(MEM_stage_inst_dmem_n13340) );
NAND2_X1 MEM_stage_inst_dmem_U9673 ( .A1(MEM_stage_inst_dmem_ram_197), .A2(MEM_stage_inst_dmem_n13350), .ZN(MEM_stage_inst_dmem_n13341) );
NAND2_X1 MEM_stage_inst_dmem_U9672 ( .A1(MEM_stage_inst_dmem_n13339), .A2(MEM_stage_inst_dmem_n13338), .ZN(MEM_stage_inst_dmem_n12545) );
NAND2_X1 MEM_stage_inst_dmem_U9671 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n13351), .ZN(MEM_stage_inst_dmem_n13338) );
NAND2_X1 MEM_stage_inst_dmem_U9670 ( .A1(MEM_stage_inst_dmem_ram_198), .A2(MEM_stage_inst_dmem_n13350), .ZN(MEM_stage_inst_dmem_n13339) );
NAND2_X1 MEM_stage_inst_dmem_U9669 ( .A1(MEM_stage_inst_dmem_n13337), .A2(MEM_stage_inst_dmem_n13336), .ZN(MEM_stage_inst_dmem_n12546) );
NAND2_X1 MEM_stage_inst_dmem_U9668 ( .A1(MEM_stage_inst_dmem_n17), .A2(MEM_stage_inst_dmem_n13351), .ZN(MEM_stage_inst_dmem_n13336) );
NAND2_X1 MEM_stage_inst_dmem_U9667 ( .A1(MEM_stage_inst_dmem_ram_199), .A2(MEM_stage_inst_dmem_n13350), .ZN(MEM_stage_inst_dmem_n13337) );
NAND2_X1 MEM_stage_inst_dmem_U9666 ( .A1(MEM_stage_inst_dmem_n13335), .A2(MEM_stage_inst_dmem_n13334), .ZN(MEM_stage_inst_dmem_n12547) );
NAND2_X1 MEM_stage_inst_dmem_U9665 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n13351), .ZN(MEM_stage_inst_dmem_n13334) );
NAND2_X1 MEM_stage_inst_dmem_U9664 ( .A1(MEM_stage_inst_dmem_ram_200), .A2(MEM_stage_inst_dmem_n13350), .ZN(MEM_stage_inst_dmem_n13335) );
NAND2_X1 MEM_stage_inst_dmem_U9663 ( .A1(MEM_stage_inst_dmem_n13333), .A2(MEM_stage_inst_dmem_n13332), .ZN(MEM_stage_inst_dmem_n12548) );
NAND2_X1 MEM_stage_inst_dmem_U9662 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n13351), .ZN(MEM_stage_inst_dmem_n13332) );
NAND2_X1 MEM_stage_inst_dmem_U9661 ( .A1(MEM_stage_inst_dmem_ram_201), .A2(MEM_stage_inst_dmem_n13350), .ZN(MEM_stage_inst_dmem_n13333) );
NAND2_X1 MEM_stage_inst_dmem_U9660 ( .A1(MEM_stage_inst_dmem_n13331), .A2(MEM_stage_inst_dmem_n13330), .ZN(MEM_stage_inst_dmem_n12549) );
NAND2_X1 MEM_stage_inst_dmem_U9659 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n13351), .ZN(MEM_stage_inst_dmem_n13330) );
NAND2_X1 MEM_stage_inst_dmem_U9658 ( .A1(MEM_stage_inst_dmem_ram_202), .A2(MEM_stage_inst_dmem_n13350), .ZN(MEM_stage_inst_dmem_n13331) );
NAND2_X1 MEM_stage_inst_dmem_U9657 ( .A1(MEM_stage_inst_dmem_n13329), .A2(MEM_stage_inst_dmem_n13328), .ZN(MEM_stage_inst_dmem_n12550) );
NAND2_X1 MEM_stage_inst_dmem_U9656 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n13351), .ZN(MEM_stage_inst_dmem_n13328) );
NAND2_X1 MEM_stage_inst_dmem_U9655 ( .A1(MEM_stage_inst_dmem_ram_203), .A2(MEM_stage_inst_dmem_n13350), .ZN(MEM_stage_inst_dmem_n13329) );
NAND2_X1 MEM_stage_inst_dmem_U9654 ( .A1(MEM_stage_inst_dmem_n13327), .A2(MEM_stage_inst_dmem_n13326), .ZN(MEM_stage_inst_dmem_n12551) );
NAND2_X1 MEM_stage_inst_dmem_U9653 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n13351), .ZN(MEM_stage_inst_dmem_n13326) );
NAND2_X1 MEM_stage_inst_dmem_U9652 ( .A1(MEM_stage_inst_dmem_ram_204), .A2(MEM_stage_inst_dmem_n13350), .ZN(MEM_stage_inst_dmem_n13327) );
NAND2_X1 MEM_stage_inst_dmem_U9651 ( .A1(MEM_stage_inst_dmem_n13325), .A2(MEM_stage_inst_dmem_n13324), .ZN(MEM_stage_inst_dmem_n12552) );
NAND2_X1 MEM_stage_inst_dmem_U9650 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n13351), .ZN(MEM_stage_inst_dmem_n13324) );
NAND2_X1 MEM_stage_inst_dmem_U9649 ( .A1(MEM_stage_inst_dmem_ram_205), .A2(MEM_stage_inst_dmem_n13350), .ZN(MEM_stage_inst_dmem_n13325) );
NAND2_X1 MEM_stage_inst_dmem_U9648 ( .A1(MEM_stage_inst_dmem_n13323), .A2(MEM_stage_inst_dmem_n13322), .ZN(MEM_stage_inst_dmem_n12553) );
NAND2_X1 MEM_stage_inst_dmem_U9647 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n13351), .ZN(MEM_stage_inst_dmem_n13322) );
NAND2_X1 MEM_stage_inst_dmem_U9646 ( .A1(MEM_stage_inst_dmem_ram_206), .A2(MEM_stage_inst_dmem_n13350), .ZN(MEM_stage_inst_dmem_n13323) );
NAND2_X1 MEM_stage_inst_dmem_U9645 ( .A1(MEM_stage_inst_dmem_n13321), .A2(MEM_stage_inst_dmem_n13320), .ZN(MEM_stage_inst_dmem_n12554) );
NAND2_X1 MEM_stage_inst_dmem_U9644 ( .A1(MEM_stage_inst_dmem_n14693), .A2(MEM_stage_inst_dmem_n13351), .ZN(MEM_stage_inst_dmem_n13320) );
INV_X1 MEM_stage_inst_dmem_U9643 ( .A(MEM_stage_inst_dmem_n13350), .ZN(MEM_stage_inst_dmem_n13351) );
NAND2_X1 MEM_stage_inst_dmem_U9642 ( .A1(MEM_stage_inst_dmem_ram_207), .A2(MEM_stage_inst_dmem_n13350), .ZN(MEM_stage_inst_dmem_n13321) );
NAND2_X1 MEM_stage_inst_dmem_U9641 ( .A1(MEM_stage_inst_dmem_n21039), .A2(MEM_stage_inst_dmem_n13728), .ZN(MEM_stage_inst_dmem_n13350) );
NAND2_X1 MEM_stage_inst_dmem_U9640 ( .A1(MEM_stage_inst_dmem_n13319), .A2(MEM_stage_inst_dmem_n13318), .ZN(MEM_stage_inst_dmem_n12555) );
NAND2_X1 MEM_stage_inst_dmem_U9639 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n13317), .ZN(MEM_stage_inst_dmem_n13318) );
NAND2_X1 MEM_stage_inst_dmem_U9638 ( .A1(MEM_stage_inst_dmem_ram_208), .A2(MEM_stage_inst_dmem_n13316), .ZN(MEM_stage_inst_dmem_n13319) );
NAND2_X1 MEM_stage_inst_dmem_U9637 ( .A1(MEM_stage_inst_dmem_n13315), .A2(MEM_stage_inst_dmem_n13314), .ZN(MEM_stage_inst_dmem_n12556) );
NAND2_X1 MEM_stage_inst_dmem_U9636 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n13317), .ZN(MEM_stage_inst_dmem_n13314) );
NAND2_X1 MEM_stage_inst_dmem_U9635 ( .A1(MEM_stage_inst_dmem_ram_209), .A2(MEM_stage_inst_dmem_n13316), .ZN(MEM_stage_inst_dmem_n13315) );
NAND2_X1 MEM_stage_inst_dmem_U9634 ( .A1(MEM_stage_inst_dmem_n13313), .A2(MEM_stage_inst_dmem_n13312), .ZN(MEM_stage_inst_dmem_n12557) );
NAND2_X1 MEM_stage_inst_dmem_U9633 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n13317), .ZN(MEM_stage_inst_dmem_n13312) );
NAND2_X1 MEM_stage_inst_dmem_U9632 ( .A1(MEM_stage_inst_dmem_ram_210), .A2(MEM_stage_inst_dmem_n13316), .ZN(MEM_stage_inst_dmem_n13313) );
NAND2_X1 MEM_stage_inst_dmem_U9631 ( .A1(MEM_stage_inst_dmem_n13311), .A2(MEM_stage_inst_dmem_n13310), .ZN(MEM_stage_inst_dmem_n12558) );
NAND2_X1 MEM_stage_inst_dmem_U9630 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n13317), .ZN(MEM_stage_inst_dmem_n13310) );
NAND2_X1 MEM_stage_inst_dmem_U9629 ( .A1(MEM_stage_inst_dmem_ram_211), .A2(MEM_stage_inst_dmem_n13316), .ZN(MEM_stage_inst_dmem_n13311) );
NAND2_X1 MEM_stage_inst_dmem_U9628 ( .A1(MEM_stage_inst_dmem_n13309), .A2(MEM_stage_inst_dmem_n13308), .ZN(MEM_stage_inst_dmem_n12559) );
NAND2_X1 MEM_stage_inst_dmem_U9627 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n13317), .ZN(MEM_stage_inst_dmem_n13308) );
NAND2_X1 MEM_stage_inst_dmem_U9626 ( .A1(MEM_stage_inst_dmem_ram_212), .A2(MEM_stage_inst_dmem_n13316), .ZN(MEM_stage_inst_dmem_n13309) );
NAND2_X1 MEM_stage_inst_dmem_U9625 ( .A1(MEM_stage_inst_dmem_n13307), .A2(MEM_stage_inst_dmem_n13306), .ZN(MEM_stage_inst_dmem_n12560) );
NAND2_X1 MEM_stage_inst_dmem_U9624 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n13317), .ZN(MEM_stage_inst_dmem_n13306) );
NAND2_X1 MEM_stage_inst_dmem_U9623 ( .A1(MEM_stage_inst_dmem_ram_213), .A2(MEM_stage_inst_dmem_n13316), .ZN(MEM_stage_inst_dmem_n13307) );
NAND2_X1 MEM_stage_inst_dmem_U9622 ( .A1(MEM_stage_inst_dmem_n13305), .A2(MEM_stage_inst_dmem_n13304), .ZN(MEM_stage_inst_dmem_n12561) );
NAND2_X1 MEM_stage_inst_dmem_U9621 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n13317), .ZN(MEM_stage_inst_dmem_n13304) );
NAND2_X1 MEM_stage_inst_dmem_U9620 ( .A1(MEM_stage_inst_dmem_ram_214), .A2(MEM_stage_inst_dmem_n13316), .ZN(MEM_stage_inst_dmem_n13305) );
NAND2_X1 MEM_stage_inst_dmem_U9619 ( .A1(MEM_stage_inst_dmem_n13303), .A2(MEM_stage_inst_dmem_n13302), .ZN(MEM_stage_inst_dmem_n12562) );
NAND2_X1 MEM_stage_inst_dmem_U9618 ( .A1(MEM_stage_inst_dmem_n13886), .A2(MEM_stage_inst_dmem_n13317), .ZN(MEM_stage_inst_dmem_n13302) );
NAND2_X1 MEM_stage_inst_dmem_U9617 ( .A1(MEM_stage_inst_dmem_ram_215), .A2(MEM_stage_inst_dmem_n13316), .ZN(MEM_stage_inst_dmem_n13303) );
NAND2_X1 MEM_stage_inst_dmem_U9616 ( .A1(MEM_stage_inst_dmem_n13301), .A2(MEM_stage_inst_dmem_n13300), .ZN(MEM_stage_inst_dmem_n12563) );
NAND2_X1 MEM_stage_inst_dmem_U9615 ( .A1(MEM_stage_inst_dmem_n13883), .A2(MEM_stage_inst_dmem_n13317), .ZN(MEM_stage_inst_dmem_n13300) );
NAND2_X1 MEM_stage_inst_dmem_U9614 ( .A1(MEM_stage_inst_dmem_ram_216), .A2(MEM_stage_inst_dmem_n13316), .ZN(MEM_stage_inst_dmem_n13301) );
NAND2_X1 MEM_stage_inst_dmem_U9613 ( .A1(MEM_stage_inst_dmem_n13299), .A2(MEM_stage_inst_dmem_n13298), .ZN(MEM_stage_inst_dmem_n12564) );
NAND2_X1 MEM_stage_inst_dmem_U9612 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n13317), .ZN(MEM_stage_inst_dmem_n13298) );
NAND2_X1 MEM_stage_inst_dmem_U9611 ( .A1(MEM_stage_inst_dmem_ram_217), .A2(MEM_stage_inst_dmem_n13316), .ZN(MEM_stage_inst_dmem_n13299) );
NAND2_X1 MEM_stage_inst_dmem_U9610 ( .A1(MEM_stage_inst_dmem_n13297), .A2(MEM_stage_inst_dmem_n13296), .ZN(MEM_stage_inst_dmem_n12565) );
NAND2_X1 MEM_stage_inst_dmem_U9609 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n13317), .ZN(MEM_stage_inst_dmem_n13296) );
NAND2_X1 MEM_stage_inst_dmem_U9608 ( .A1(MEM_stage_inst_dmem_ram_218), .A2(MEM_stage_inst_dmem_n13316), .ZN(MEM_stage_inst_dmem_n13297) );
NAND2_X1 MEM_stage_inst_dmem_U9607 ( .A1(MEM_stage_inst_dmem_n13295), .A2(MEM_stage_inst_dmem_n13294), .ZN(MEM_stage_inst_dmem_n12566) );
NAND2_X1 MEM_stage_inst_dmem_U9606 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n13317), .ZN(MEM_stage_inst_dmem_n13294) );
NAND2_X1 MEM_stage_inst_dmem_U9605 ( .A1(MEM_stage_inst_dmem_ram_219), .A2(MEM_stage_inst_dmem_n13316), .ZN(MEM_stage_inst_dmem_n13295) );
NAND2_X1 MEM_stage_inst_dmem_U9604 ( .A1(MEM_stage_inst_dmem_n13293), .A2(MEM_stage_inst_dmem_n13292), .ZN(MEM_stage_inst_dmem_n12567) );
NAND2_X1 MEM_stage_inst_dmem_U9603 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n13317), .ZN(MEM_stage_inst_dmem_n13292) );
NAND2_X1 MEM_stage_inst_dmem_U9602 ( .A1(MEM_stage_inst_dmem_ram_220), .A2(MEM_stage_inst_dmem_n13316), .ZN(MEM_stage_inst_dmem_n13293) );
NAND2_X1 MEM_stage_inst_dmem_U9601 ( .A1(MEM_stage_inst_dmem_n13291), .A2(MEM_stage_inst_dmem_n13290), .ZN(MEM_stage_inst_dmem_n12568) );
NAND2_X1 MEM_stage_inst_dmem_U9600 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n13317), .ZN(MEM_stage_inst_dmem_n13290) );
NAND2_X1 MEM_stage_inst_dmem_U9599 ( .A1(MEM_stage_inst_dmem_ram_221), .A2(MEM_stage_inst_dmem_n13316), .ZN(MEM_stage_inst_dmem_n13291) );
NAND2_X1 MEM_stage_inst_dmem_U9598 ( .A1(MEM_stage_inst_dmem_n13289), .A2(MEM_stage_inst_dmem_n13288), .ZN(MEM_stage_inst_dmem_n12569) );
NAND2_X1 MEM_stage_inst_dmem_U9597 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n13317), .ZN(MEM_stage_inst_dmem_n13288) );
NAND2_X1 MEM_stage_inst_dmem_U9596 ( .A1(MEM_stage_inst_dmem_ram_222), .A2(MEM_stage_inst_dmem_n13316), .ZN(MEM_stage_inst_dmem_n13289) );
NAND2_X1 MEM_stage_inst_dmem_U9595 ( .A1(MEM_stage_inst_dmem_n13287), .A2(MEM_stage_inst_dmem_n13286), .ZN(MEM_stage_inst_dmem_n12570) );
NAND2_X1 MEM_stage_inst_dmem_U9594 ( .A1(MEM_stage_inst_dmem_n21320), .A2(MEM_stage_inst_dmem_n13317), .ZN(MEM_stage_inst_dmem_n13286) );
INV_X1 MEM_stage_inst_dmem_U9593 ( .A(MEM_stage_inst_dmem_n13316), .ZN(MEM_stage_inst_dmem_n13317) );
NAND2_X1 MEM_stage_inst_dmem_U9592 ( .A1(MEM_stage_inst_dmem_ram_223), .A2(MEM_stage_inst_dmem_n13316), .ZN(MEM_stage_inst_dmem_n13287) );
NAND2_X1 MEM_stage_inst_dmem_U9591 ( .A1(MEM_stage_inst_dmem_n21004), .A2(MEM_stage_inst_dmem_n13728), .ZN(MEM_stage_inst_dmem_n13316) );
NAND2_X1 MEM_stage_inst_dmem_U9590 ( .A1(MEM_stage_inst_dmem_n13285), .A2(MEM_stage_inst_dmem_n13284), .ZN(MEM_stage_inst_dmem_n12571) );
NAND2_X1 MEM_stage_inst_dmem_U9589 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n13283), .ZN(MEM_stage_inst_dmem_n13284) );
NAND2_X1 MEM_stage_inst_dmem_U9588 ( .A1(MEM_stage_inst_dmem_ram_224), .A2(MEM_stage_inst_dmem_n13282), .ZN(MEM_stage_inst_dmem_n13285) );
NAND2_X1 MEM_stage_inst_dmem_U9587 ( .A1(MEM_stage_inst_dmem_n13281), .A2(MEM_stage_inst_dmem_n13280), .ZN(MEM_stage_inst_dmem_n12572) );
NAND2_X1 MEM_stage_inst_dmem_U9586 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n13283), .ZN(MEM_stage_inst_dmem_n13280) );
NAND2_X1 MEM_stage_inst_dmem_U9585 ( .A1(MEM_stage_inst_dmem_ram_225), .A2(MEM_stage_inst_dmem_n13282), .ZN(MEM_stage_inst_dmem_n13281) );
NAND2_X1 MEM_stage_inst_dmem_U9584 ( .A1(MEM_stage_inst_dmem_n13279), .A2(MEM_stage_inst_dmem_n13278), .ZN(MEM_stage_inst_dmem_n12573) );
NAND2_X1 MEM_stage_inst_dmem_U9583 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n13283), .ZN(MEM_stage_inst_dmem_n13278) );
NAND2_X1 MEM_stage_inst_dmem_U9582 ( .A1(MEM_stage_inst_dmem_ram_226), .A2(MEM_stage_inst_dmem_n13282), .ZN(MEM_stage_inst_dmem_n13279) );
NAND2_X1 MEM_stage_inst_dmem_U9581 ( .A1(MEM_stage_inst_dmem_n13277), .A2(MEM_stage_inst_dmem_n13276), .ZN(MEM_stage_inst_dmem_n12574) );
NAND2_X1 MEM_stage_inst_dmem_U9580 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n13283), .ZN(MEM_stage_inst_dmem_n13276) );
NAND2_X1 MEM_stage_inst_dmem_U9579 ( .A1(MEM_stage_inst_dmem_ram_227), .A2(MEM_stage_inst_dmem_n13282), .ZN(MEM_stage_inst_dmem_n13277) );
NAND2_X1 MEM_stage_inst_dmem_U9578 ( .A1(MEM_stage_inst_dmem_n13275), .A2(MEM_stage_inst_dmem_n13274), .ZN(MEM_stage_inst_dmem_n12575) );
NAND2_X1 MEM_stage_inst_dmem_U9577 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n13283), .ZN(MEM_stage_inst_dmem_n13274) );
NAND2_X1 MEM_stage_inst_dmem_U9576 ( .A1(MEM_stage_inst_dmem_ram_228), .A2(MEM_stage_inst_dmem_n13282), .ZN(MEM_stage_inst_dmem_n13275) );
NAND2_X1 MEM_stage_inst_dmem_U9575 ( .A1(MEM_stage_inst_dmem_n13273), .A2(MEM_stage_inst_dmem_n13272), .ZN(MEM_stage_inst_dmem_n12576) );
NAND2_X1 MEM_stage_inst_dmem_U9574 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n13283), .ZN(MEM_stage_inst_dmem_n13272) );
NAND2_X1 MEM_stage_inst_dmem_U9573 ( .A1(MEM_stage_inst_dmem_ram_229), .A2(MEM_stage_inst_dmem_n13282), .ZN(MEM_stage_inst_dmem_n13273) );
NAND2_X1 MEM_stage_inst_dmem_U9572 ( .A1(MEM_stage_inst_dmem_n13271), .A2(MEM_stage_inst_dmem_n13270), .ZN(MEM_stage_inst_dmem_n12577) );
NAND2_X1 MEM_stage_inst_dmem_U9571 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n13283), .ZN(MEM_stage_inst_dmem_n13270) );
NAND2_X1 MEM_stage_inst_dmem_U9570 ( .A1(MEM_stage_inst_dmem_ram_230), .A2(MEM_stage_inst_dmem_n13282), .ZN(MEM_stage_inst_dmem_n13271) );
NAND2_X1 MEM_stage_inst_dmem_U9569 ( .A1(MEM_stage_inst_dmem_n13269), .A2(MEM_stage_inst_dmem_n13268), .ZN(MEM_stage_inst_dmem_n12578) );
NAND2_X1 MEM_stage_inst_dmem_U9568 ( .A1(MEM_stage_inst_dmem_n18), .A2(MEM_stage_inst_dmem_n13283), .ZN(MEM_stage_inst_dmem_n13268) );
NAND2_X1 MEM_stage_inst_dmem_U9567 ( .A1(MEM_stage_inst_dmem_ram_231), .A2(MEM_stage_inst_dmem_n13282), .ZN(MEM_stage_inst_dmem_n13269) );
NAND2_X1 MEM_stage_inst_dmem_U9566 ( .A1(MEM_stage_inst_dmem_n13267), .A2(MEM_stage_inst_dmem_n13266), .ZN(MEM_stage_inst_dmem_n12579) );
NAND2_X1 MEM_stage_inst_dmem_U9565 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n13283), .ZN(MEM_stage_inst_dmem_n13266) );
NAND2_X1 MEM_stage_inst_dmem_U9564 ( .A1(MEM_stage_inst_dmem_ram_232), .A2(MEM_stage_inst_dmem_n13282), .ZN(MEM_stage_inst_dmem_n13267) );
NAND2_X1 MEM_stage_inst_dmem_U9563 ( .A1(MEM_stage_inst_dmem_n13265), .A2(MEM_stage_inst_dmem_n13264), .ZN(MEM_stage_inst_dmem_n12580) );
NAND2_X1 MEM_stage_inst_dmem_U9562 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n13283), .ZN(MEM_stage_inst_dmem_n13264) );
NAND2_X1 MEM_stage_inst_dmem_U9561 ( .A1(MEM_stage_inst_dmem_ram_233), .A2(MEM_stage_inst_dmem_n13282), .ZN(MEM_stage_inst_dmem_n13265) );
NAND2_X1 MEM_stage_inst_dmem_U9560 ( .A1(MEM_stage_inst_dmem_n13263), .A2(MEM_stage_inst_dmem_n13262), .ZN(MEM_stage_inst_dmem_n12581) );
NAND2_X1 MEM_stage_inst_dmem_U9559 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n13283), .ZN(MEM_stage_inst_dmem_n13262) );
NAND2_X1 MEM_stage_inst_dmem_U9558 ( .A1(MEM_stage_inst_dmem_ram_234), .A2(MEM_stage_inst_dmem_n13282), .ZN(MEM_stage_inst_dmem_n13263) );
NAND2_X1 MEM_stage_inst_dmem_U9557 ( .A1(MEM_stage_inst_dmem_n13261), .A2(MEM_stage_inst_dmem_n13260), .ZN(MEM_stage_inst_dmem_n12582) );
NAND2_X1 MEM_stage_inst_dmem_U9556 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n13283), .ZN(MEM_stage_inst_dmem_n13260) );
NAND2_X1 MEM_stage_inst_dmem_U9555 ( .A1(MEM_stage_inst_dmem_ram_235), .A2(MEM_stage_inst_dmem_n13282), .ZN(MEM_stage_inst_dmem_n13261) );
NAND2_X1 MEM_stage_inst_dmem_U9554 ( .A1(MEM_stage_inst_dmem_n13259), .A2(MEM_stage_inst_dmem_n13258), .ZN(MEM_stage_inst_dmem_n12583) );
NAND2_X1 MEM_stage_inst_dmem_U9553 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n13283), .ZN(MEM_stage_inst_dmem_n13258) );
NAND2_X1 MEM_stage_inst_dmem_U9552 ( .A1(MEM_stage_inst_dmem_ram_236), .A2(MEM_stage_inst_dmem_n13282), .ZN(MEM_stage_inst_dmem_n13259) );
NAND2_X1 MEM_stage_inst_dmem_U9551 ( .A1(MEM_stage_inst_dmem_n13257), .A2(MEM_stage_inst_dmem_n13256), .ZN(MEM_stage_inst_dmem_n12584) );
NAND2_X1 MEM_stage_inst_dmem_U9550 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n13283), .ZN(MEM_stage_inst_dmem_n13256) );
NAND2_X1 MEM_stage_inst_dmem_U9549 ( .A1(MEM_stage_inst_dmem_ram_237), .A2(MEM_stage_inst_dmem_n13282), .ZN(MEM_stage_inst_dmem_n13257) );
NAND2_X1 MEM_stage_inst_dmem_U9548 ( .A1(MEM_stage_inst_dmem_n13255), .A2(MEM_stage_inst_dmem_n13254), .ZN(MEM_stage_inst_dmem_n12585) );
NAND2_X1 MEM_stage_inst_dmem_U9547 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n13283), .ZN(MEM_stage_inst_dmem_n13254) );
NAND2_X1 MEM_stage_inst_dmem_U9546 ( .A1(MEM_stage_inst_dmem_ram_238), .A2(MEM_stage_inst_dmem_n13282), .ZN(MEM_stage_inst_dmem_n13255) );
NAND2_X1 MEM_stage_inst_dmem_U9545 ( .A1(MEM_stage_inst_dmem_n13253), .A2(MEM_stage_inst_dmem_n13252), .ZN(MEM_stage_inst_dmem_n12586) );
NAND2_X1 MEM_stage_inst_dmem_U9544 ( .A1(MEM_stage_inst_dmem_n14693), .A2(MEM_stage_inst_dmem_n13283), .ZN(MEM_stage_inst_dmem_n13252) );
INV_X1 MEM_stage_inst_dmem_U9543 ( .A(MEM_stage_inst_dmem_n13282), .ZN(MEM_stage_inst_dmem_n13283) );
NAND2_X1 MEM_stage_inst_dmem_U9542 ( .A1(MEM_stage_inst_dmem_ram_239), .A2(MEM_stage_inst_dmem_n13282), .ZN(MEM_stage_inst_dmem_n13253) );
NAND2_X1 MEM_stage_inst_dmem_U9541 ( .A1(MEM_stage_inst_dmem_n20969), .A2(MEM_stage_inst_dmem_n13728), .ZN(MEM_stage_inst_dmem_n13282) );
NAND2_X1 MEM_stage_inst_dmem_U9540 ( .A1(MEM_stage_inst_dmem_n13251), .A2(MEM_stage_inst_dmem_n13250), .ZN(MEM_stage_inst_dmem_n12587) );
NAND2_X1 MEM_stage_inst_dmem_U9539 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n13249), .ZN(MEM_stage_inst_dmem_n13250) );
NAND2_X1 MEM_stage_inst_dmem_U9538 ( .A1(MEM_stage_inst_dmem_ram_240), .A2(MEM_stage_inst_dmem_n13248), .ZN(MEM_stage_inst_dmem_n13251) );
NAND2_X1 MEM_stage_inst_dmem_U9537 ( .A1(MEM_stage_inst_dmem_n13247), .A2(MEM_stage_inst_dmem_n13246), .ZN(MEM_stage_inst_dmem_n12588) );
NAND2_X1 MEM_stage_inst_dmem_U9536 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n13249), .ZN(MEM_stage_inst_dmem_n13246) );
NAND2_X1 MEM_stage_inst_dmem_U9535 ( .A1(MEM_stage_inst_dmem_ram_241), .A2(MEM_stage_inst_dmem_n13248), .ZN(MEM_stage_inst_dmem_n13247) );
NAND2_X1 MEM_stage_inst_dmem_U9534 ( .A1(MEM_stage_inst_dmem_n13245), .A2(MEM_stage_inst_dmem_n13244), .ZN(MEM_stage_inst_dmem_n12589) );
NAND2_X1 MEM_stage_inst_dmem_U9533 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n13249), .ZN(MEM_stage_inst_dmem_n13244) );
NAND2_X1 MEM_stage_inst_dmem_U9532 ( .A1(MEM_stage_inst_dmem_ram_242), .A2(MEM_stage_inst_dmem_n13248), .ZN(MEM_stage_inst_dmem_n13245) );
NAND2_X1 MEM_stage_inst_dmem_U9531 ( .A1(MEM_stage_inst_dmem_n13243), .A2(MEM_stage_inst_dmem_n13242), .ZN(MEM_stage_inst_dmem_n12590) );
NAND2_X1 MEM_stage_inst_dmem_U9530 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n13249), .ZN(MEM_stage_inst_dmem_n13242) );
NAND2_X1 MEM_stage_inst_dmem_U9529 ( .A1(MEM_stage_inst_dmem_ram_243), .A2(MEM_stage_inst_dmem_n13248), .ZN(MEM_stage_inst_dmem_n13243) );
NAND2_X1 MEM_stage_inst_dmem_U9528 ( .A1(MEM_stage_inst_dmem_n13241), .A2(MEM_stage_inst_dmem_n13240), .ZN(MEM_stage_inst_dmem_n12591) );
NAND2_X1 MEM_stage_inst_dmem_U9527 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n13249), .ZN(MEM_stage_inst_dmem_n13240) );
NAND2_X1 MEM_stage_inst_dmem_U9526 ( .A1(MEM_stage_inst_dmem_ram_244), .A2(MEM_stage_inst_dmem_n13248), .ZN(MEM_stage_inst_dmem_n13241) );
NAND2_X1 MEM_stage_inst_dmem_U9525 ( .A1(MEM_stage_inst_dmem_n13239), .A2(MEM_stage_inst_dmem_n13238), .ZN(MEM_stage_inst_dmem_n12592) );
NAND2_X1 MEM_stage_inst_dmem_U9524 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n13249), .ZN(MEM_stage_inst_dmem_n13238) );
NAND2_X1 MEM_stage_inst_dmem_U9523 ( .A1(MEM_stage_inst_dmem_ram_245), .A2(MEM_stage_inst_dmem_n13248), .ZN(MEM_stage_inst_dmem_n13239) );
NAND2_X1 MEM_stage_inst_dmem_U9522 ( .A1(MEM_stage_inst_dmem_n13237), .A2(MEM_stage_inst_dmem_n13236), .ZN(MEM_stage_inst_dmem_n12593) );
NAND2_X1 MEM_stage_inst_dmem_U9521 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n13249), .ZN(MEM_stage_inst_dmem_n13236) );
NAND2_X1 MEM_stage_inst_dmem_U9520 ( .A1(MEM_stage_inst_dmem_ram_246), .A2(MEM_stage_inst_dmem_n13248), .ZN(MEM_stage_inst_dmem_n13237) );
NAND2_X1 MEM_stage_inst_dmem_U9519 ( .A1(MEM_stage_inst_dmem_n13235), .A2(MEM_stage_inst_dmem_n13234), .ZN(MEM_stage_inst_dmem_n12594) );
NAND2_X1 MEM_stage_inst_dmem_U9518 ( .A1(MEM_stage_inst_dmem_n13886), .A2(MEM_stage_inst_dmem_n13249), .ZN(MEM_stage_inst_dmem_n13234) );
NAND2_X1 MEM_stage_inst_dmem_U9517 ( .A1(MEM_stage_inst_dmem_ram_247), .A2(MEM_stage_inst_dmem_n13248), .ZN(MEM_stage_inst_dmem_n13235) );
NAND2_X1 MEM_stage_inst_dmem_U9516 ( .A1(MEM_stage_inst_dmem_n13233), .A2(MEM_stage_inst_dmem_n13232), .ZN(MEM_stage_inst_dmem_n12595) );
NAND2_X1 MEM_stage_inst_dmem_U9515 ( .A1(MEM_stage_inst_dmem_n13883), .A2(MEM_stage_inst_dmem_n13249), .ZN(MEM_stage_inst_dmem_n13232) );
NAND2_X1 MEM_stage_inst_dmem_U9514 ( .A1(MEM_stage_inst_dmem_ram_248), .A2(MEM_stage_inst_dmem_n13248), .ZN(MEM_stage_inst_dmem_n13233) );
NAND2_X1 MEM_stage_inst_dmem_U9513 ( .A1(MEM_stage_inst_dmem_n13231), .A2(MEM_stage_inst_dmem_n13230), .ZN(MEM_stage_inst_dmem_n12596) );
NAND2_X1 MEM_stage_inst_dmem_U9512 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n13249), .ZN(MEM_stage_inst_dmem_n13230) );
NAND2_X1 MEM_stage_inst_dmem_U9511 ( .A1(MEM_stage_inst_dmem_ram_249), .A2(MEM_stage_inst_dmem_n13248), .ZN(MEM_stage_inst_dmem_n13231) );
NAND2_X1 MEM_stage_inst_dmem_U9510 ( .A1(MEM_stage_inst_dmem_n13229), .A2(MEM_stage_inst_dmem_n13228), .ZN(MEM_stage_inst_dmem_n12597) );
NAND2_X1 MEM_stage_inst_dmem_U9509 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n13249), .ZN(MEM_stage_inst_dmem_n13228) );
NAND2_X1 MEM_stage_inst_dmem_U9508 ( .A1(MEM_stage_inst_dmem_ram_250), .A2(MEM_stage_inst_dmem_n13248), .ZN(MEM_stage_inst_dmem_n13229) );
NAND2_X1 MEM_stage_inst_dmem_U9507 ( .A1(MEM_stage_inst_dmem_n13227), .A2(MEM_stage_inst_dmem_n13226), .ZN(MEM_stage_inst_dmem_n12598) );
NAND2_X1 MEM_stage_inst_dmem_U9506 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n13249), .ZN(MEM_stage_inst_dmem_n13226) );
NAND2_X1 MEM_stage_inst_dmem_U9505 ( .A1(MEM_stage_inst_dmem_ram_251), .A2(MEM_stage_inst_dmem_n13248), .ZN(MEM_stage_inst_dmem_n13227) );
NAND2_X1 MEM_stage_inst_dmem_U9504 ( .A1(MEM_stage_inst_dmem_n13225), .A2(MEM_stage_inst_dmem_n13224), .ZN(MEM_stage_inst_dmem_n12599) );
NAND2_X1 MEM_stage_inst_dmem_U9503 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n13249), .ZN(MEM_stage_inst_dmem_n13224) );
NAND2_X1 MEM_stage_inst_dmem_U9502 ( .A1(MEM_stage_inst_dmem_ram_252), .A2(MEM_stage_inst_dmem_n13248), .ZN(MEM_stage_inst_dmem_n13225) );
NAND2_X1 MEM_stage_inst_dmem_U9501 ( .A1(MEM_stage_inst_dmem_n13223), .A2(MEM_stage_inst_dmem_n13222), .ZN(MEM_stage_inst_dmem_n12600) );
NAND2_X1 MEM_stage_inst_dmem_U9500 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n13249), .ZN(MEM_stage_inst_dmem_n13222) );
NAND2_X1 MEM_stage_inst_dmem_U9499 ( .A1(MEM_stage_inst_dmem_ram_253), .A2(MEM_stage_inst_dmem_n13248), .ZN(MEM_stage_inst_dmem_n13223) );
NAND2_X1 MEM_stage_inst_dmem_U9498 ( .A1(MEM_stage_inst_dmem_n13221), .A2(MEM_stage_inst_dmem_n13220), .ZN(MEM_stage_inst_dmem_n12601) );
NAND2_X1 MEM_stage_inst_dmem_U9497 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n13249), .ZN(MEM_stage_inst_dmem_n13220) );
NAND2_X1 MEM_stage_inst_dmem_U9496 ( .A1(MEM_stage_inst_dmem_ram_254), .A2(MEM_stage_inst_dmem_n13248), .ZN(MEM_stage_inst_dmem_n13221) );
NAND2_X1 MEM_stage_inst_dmem_U9495 ( .A1(MEM_stage_inst_dmem_n13219), .A2(MEM_stage_inst_dmem_n13218), .ZN(MEM_stage_inst_dmem_n12602) );
NAND2_X1 MEM_stage_inst_dmem_U9494 ( .A1(MEM_stage_inst_dmem_n15110), .A2(MEM_stage_inst_dmem_n13249), .ZN(MEM_stage_inst_dmem_n13218) );
INV_X1 MEM_stage_inst_dmem_U9493 ( .A(MEM_stage_inst_dmem_n13248), .ZN(MEM_stage_inst_dmem_n13249) );
NAND2_X1 MEM_stage_inst_dmem_U9492 ( .A1(MEM_stage_inst_dmem_ram_255), .A2(MEM_stage_inst_dmem_n13248), .ZN(MEM_stage_inst_dmem_n13219) );
NAND2_X1 MEM_stage_inst_dmem_U9491 ( .A1(MEM_stage_inst_dmem_n20934), .A2(MEM_stage_inst_dmem_n13728), .ZN(MEM_stage_inst_dmem_n13248) );
NOR2_X2 MEM_stage_inst_dmem_U9490 ( .A1(MEM_stage_inst_dmem_n17619), .A2(MEM_stage_inst_dmem_n16519), .ZN(MEM_stage_inst_dmem_n13728) );
NAND2_X1 MEM_stage_inst_dmem_U9489 ( .A1(MEM_stage_inst_dmem_n13217), .A2(MEM_stage_inst_dmem_n17617), .ZN(MEM_stage_inst_dmem_n16519) );
INV_X1 MEM_stage_inst_dmem_U9488 ( .A(EX_pipeline_reg_out_26), .ZN(MEM_stage_inst_dmem_n17617) );
NAND2_X1 MEM_stage_inst_dmem_U9487 ( .A1(MEM_stage_inst_dmem_n13216), .A2(MEM_stage_inst_dmem_n13215), .ZN(MEM_stage_inst_dmem_n12603) );
NAND2_X1 MEM_stage_inst_dmem_U9486 ( .A1(MEM_stage_inst_dmem_n15145), .A2(MEM_stage_inst_dmem_n13214), .ZN(MEM_stage_inst_dmem_n13215) );
NAND2_X1 MEM_stage_inst_dmem_U9485 ( .A1(MEM_stage_inst_dmem_ram_256), .A2(MEM_stage_inst_dmem_n13213), .ZN(MEM_stage_inst_dmem_n13216) );
NAND2_X1 MEM_stage_inst_dmem_U9484 ( .A1(MEM_stage_inst_dmem_n13212), .A2(MEM_stage_inst_dmem_n13211), .ZN(MEM_stage_inst_dmem_n12604) );
NAND2_X1 MEM_stage_inst_dmem_U9483 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n13214), .ZN(MEM_stage_inst_dmem_n13211) );
NAND2_X1 MEM_stage_inst_dmem_U9482 ( .A1(MEM_stage_inst_dmem_ram_257), .A2(MEM_stage_inst_dmem_n13213), .ZN(MEM_stage_inst_dmem_n13212) );
NAND2_X1 MEM_stage_inst_dmem_U9481 ( .A1(MEM_stage_inst_dmem_n13210), .A2(MEM_stage_inst_dmem_n13209), .ZN(MEM_stage_inst_dmem_n12605) );
NAND2_X1 MEM_stage_inst_dmem_U9480 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n13214), .ZN(MEM_stage_inst_dmem_n13209) );
NAND2_X1 MEM_stage_inst_dmem_U9479 ( .A1(MEM_stage_inst_dmem_ram_258), .A2(MEM_stage_inst_dmem_n13213), .ZN(MEM_stage_inst_dmem_n13210) );
NAND2_X1 MEM_stage_inst_dmem_U9478 ( .A1(MEM_stage_inst_dmem_n13208), .A2(MEM_stage_inst_dmem_n13207), .ZN(MEM_stage_inst_dmem_n12606) );
NAND2_X1 MEM_stage_inst_dmem_U9477 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n13214), .ZN(MEM_stage_inst_dmem_n13207) );
NAND2_X1 MEM_stage_inst_dmem_U9476 ( .A1(MEM_stage_inst_dmem_ram_259), .A2(MEM_stage_inst_dmem_n13213), .ZN(MEM_stage_inst_dmem_n13208) );
NAND2_X1 MEM_stage_inst_dmem_U9475 ( .A1(MEM_stage_inst_dmem_n13206), .A2(MEM_stage_inst_dmem_n13205), .ZN(MEM_stage_inst_dmem_n12607) );
NAND2_X1 MEM_stage_inst_dmem_U9474 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n13214), .ZN(MEM_stage_inst_dmem_n13205) );
NAND2_X1 MEM_stage_inst_dmem_U9473 ( .A1(MEM_stage_inst_dmem_ram_260), .A2(MEM_stage_inst_dmem_n13213), .ZN(MEM_stage_inst_dmem_n13206) );
NAND2_X1 MEM_stage_inst_dmem_U9472 ( .A1(MEM_stage_inst_dmem_n13204), .A2(MEM_stage_inst_dmem_n13203), .ZN(MEM_stage_inst_dmem_n12608) );
NAND2_X1 MEM_stage_inst_dmem_U9471 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n13214), .ZN(MEM_stage_inst_dmem_n13203) );
NAND2_X1 MEM_stage_inst_dmem_U9470 ( .A1(MEM_stage_inst_dmem_ram_261), .A2(MEM_stage_inst_dmem_n13213), .ZN(MEM_stage_inst_dmem_n13204) );
NAND2_X1 MEM_stage_inst_dmem_U9469 ( .A1(MEM_stage_inst_dmem_n13202), .A2(MEM_stage_inst_dmem_n13201), .ZN(MEM_stage_inst_dmem_n12609) );
NAND2_X1 MEM_stage_inst_dmem_U9468 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n13214), .ZN(MEM_stage_inst_dmem_n13201) );
NAND2_X1 MEM_stage_inst_dmem_U9467 ( .A1(MEM_stage_inst_dmem_ram_262), .A2(MEM_stage_inst_dmem_n13213), .ZN(MEM_stage_inst_dmem_n13202) );
NAND2_X1 MEM_stage_inst_dmem_U9466 ( .A1(MEM_stage_inst_dmem_n13200), .A2(MEM_stage_inst_dmem_n13199), .ZN(MEM_stage_inst_dmem_n12610) );
NAND2_X1 MEM_stage_inst_dmem_U9465 ( .A1(MEM_stage_inst_dmem_n17), .A2(MEM_stage_inst_dmem_n13214), .ZN(MEM_stage_inst_dmem_n13199) );
NAND2_X1 MEM_stage_inst_dmem_U9464 ( .A1(MEM_stage_inst_dmem_ram_263), .A2(MEM_stage_inst_dmem_n13213), .ZN(MEM_stage_inst_dmem_n13200) );
NAND2_X1 MEM_stage_inst_dmem_U9463 ( .A1(MEM_stage_inst_dmem_n13198), .A2(MEM_stage_inst_dmem_n13197), .ZN(MEM_stage_inst_dmem_n12611) );
NAND2_X1 MEM_stage_inst_dmem_U9462 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n13214), .ZN(MEM_stage_inst_dmem_n13197) );
NAND2_X1 MEM_stage_inst_dmem_U9461 ( .A1(MEM_stage_inst_dmem_ram_264), .A2(MEM_stage_inst_dmem_n13213), .ZN(MEM_stage_inst_dmem_n13198) );
NAND2_X1 MEM_stage_inst_dmem_U9460 ( .A1(MEM_stage_inst_dmem_n13196), .A2(MEM_stage_inst_dmem_n13195), .ZN(MEM_stage_inst_dmem_n12612) );
NAND2_X1 MEM_stage_inst_dmem_U9459 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n13214), .ZN(MEM_stage_inst_dmem_n13195) );
NAND2_X1 MEM_stage_inst_dmem_U9458 ( .A1(MEM_stage_inst_dmem_ram_265), .A2(MEM_stage_inst_dmem_n13213), .ZN(MEM_stage_inst_dmem_n13196) );
NAND2_X1 MEM_stage_inst_dmem_U9457 ( .A1(MEM_stage_inst_dmem_n13194), .A2(MEM_stage_inst_dmem_n13193), .ZN(MEM_stage_inst_dmem_n12613) );
NAND2_X1 MEM_stage_inst_dmem_U9456 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n13214), .ZN(MEM_stage_inst_dmem_n13193) );
NAND2_X1 MEM_stage_inst_dmem_U9455 ( .A1(MEM_stage_inst_dmem_ram_266), .A2(MEM_stage_inst_dmem_n13213), .ZN(MEM_stage_inst_dmem_n13194) );
NAND2_X1 MEM_stage_inst_dmem_U9454 ( .A1(MEM_stage_inst_dmem_n13192), .A2(MEM_stage_inst_dmem_n13191), .ZN(MEM_stage_inst_dmem_n12614) );
NAND2_X1 MEM_stage_inst_dmem_U9453 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n13214), .ZN(MEM_stage_inst_dmem_n13191) );
NAND2_X1 MEM_stage_inst_dmem_U9452 ( .A1(MEM_stage_inst_dmem_ram_267), .A2(MEM_stage_inst_dmem_n13213), .ZN(MEM_stage_inst_dmem_n13192) );
NAND2_X1 MEM_stage_inst_dmem_U9451 ( .A1(MEM_stage_inst_dmem_n13190), .A2(MEM_stage_inst_dmem_n13189), .ZN(MEM_stage_inst_dmem_n12615) );
NAND2_X1 MEM_stage_inst_dmem_U9450 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n13214), .ZN(MEM_stage_inst_dmem_n13189) );
NAND2_X1 MEM_stage_inst_dmem_U9449 ( .A1(MEM_stage_inst_dmem_ram_268), .A2(MEM_stage_inst_dmem_n13213), .ZN(MEM_stage_inst_dmem_n13190) );
NAND2_X1 MEM_stage_inst_dmem_U9448 ( .A1(MEM_stage_inst_dmem_n13188), .A2(MEM_stage_inst_dmem_n13187), .ZN(MEM_stage_inst_dmem_n12616) );
NAND2_X1 MEM_stage_inst_dmem_U9447 ( .A1(MEM_stage_inst_dmem_n15116), .A2(MEM_stage_inst_dmem_n13214), .ZN(MEM_stage_inst_dmem_n13187) );
NAND2_X1 MEM_stage_inst_dmem_U9446 ( .A1(MEM_stage_inst_dmem_ram_269), .A2(MEM_stage_inst_dmem_n13213), .ZN(MEM_stage_inst_dmem_n13188) );
NAND2_X1 MEM_stage_inst_dmem_U9445 ( .A1(MEM_stage_inst_dmem_n13186), .A2(MEM_stage_inst_dmem_n13185), .ZN(MEM_stage_inst_dmem_n12617) );
NAND2_X1 MEM_stage_inst_dmem_U9444 ( .A1(MEM_stage_inst_dmem_n15113), .A2(MEM_stage_inst_dmem_n13214), .ZN(MEM_stage_inst_dmem_n13185) );
NAND2_X1 MEM_stage_inst_dmem_U9443 ( .A1(MEM_stage_inst_dmem_ram_270), .A2(MEM_stage_inst_dmem_n13213), .ZN(MEM_stage_inst_dmem_n13186) );
NAND2_X1 MEM_stage_inst_dmem_U9442 ( .A1(MEM_stage_inst_dmem_n13184), .A2(MEM_stage_inst_dmem_n13183), .ZN(MEM_stage_inst_dmem_n12618) );
NAND2_X1 MEM_stage_inst_dmem_U9441 ( .A1(MEM_stage_inst_dmem_n15110), .A2(MEM_stage_inst_dmem_n13214), .ZN(MEM_stage_inst_dmem_n13183) );
INV_X1 MEM_stage_inst_dmem_U9440 ( .A(MEM_stage_inst_dmem_n13213), .ZN(MEM_stage_inst_dmem_n13214) );
NAND2_X1 MEM_stage_inst_dmem_U9439 ( .A1(MEM_stage_inst_dmem_ram_271), .A2(MEM_stage_inst_dmem_n13213), .ZN(MEM_stage_inst_dmem_n13184) );
NAND2_X1 MEM_stage_inst_dmem_U9438 ( .A1(MEM_stage_inst_dmem_n13182), .A2(MEM_stage_inst_dmem_n21465), .ZN(MEM_stage_inst_dmem_n13213) );
NOR2_X2 MEM_stage_inst_dmem_U9437 ( .A1(MEM_stage_inst_dmem_n13181), .A2(MEM_stage_inst_dmem_n13180), .ZN(MEM_stage_inst_dmem_n21465) );
NAND2_X1 MEM_stage_inst_dmem_U9436 ( .A1(MEM_stage_inst_dmem_n13179), .A2(MEM_stage_inst_dmem_n13178), .ZN(MEM_stage_inst_dmem_n12619) );
NAND2_X1 MEM_stage_inst_dmem_U9435 ( .A1(MEM_stage_inst_dmem_n15145), .A2(MEM_stage_inst_dmem_n13177), .ZN(MEM_stage_inst_dmem_n13178) );
NAND2_X1 MEM_stage_inst_dmem_U9434 ( .A1(MEM_stage_inst_dmem_ram_272), .A2(MEM_stage_inst_dmem_n13176), .ZN(MEM_stage_inst_dmem_n13179) );
NAND2_X1 MEM_stage_inst_dmem_U9433 ( .A1(MEM_stage_inst_dmem_n13175), .A2(MEM_stage_inst_dmem_n13174), .ZN(MEM_stage_inst_dmem_n12620) );
NAND2_X1 MEM_stage_inst_dmem_U9432 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n13177), .ZN(MEM_stage_inst_dmem_n13174) );
NAND2_X1 MEM_stage_inst_dmem_U9431 ( .A1(MEM_stage_inst_dmem_ram_273), .A2(MEM_stage_inst_dmem_n13176), .ZN(MEM_stage_inst_dmem_n13175) );
NAND2_X1 MEM_stage_inst_dmem_U9430 ( .A1(MEM_stage_inst_dmem_n13173), .A2(MEM_stage_inst_dmem_n13172), .ZN(MEM_stage_inst_dmem_n12621) );
NAND2_X1 MEM_stage_inst_dmem_U9429 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n13177), .ZN(MEM_stage_inst_dmem_n13172) );
NAND2_X1 MEM_stage_inst_dmem_U9428 ( .A1(MEM_stage_inst_dmem_ram_274), .A2(MEM_stage_inst_dmem_n13176), .ZN(MEM_stage_inst_dmem_n13173) );
NAND2_X1 MEM_stage_inst_dmem_U9427 ( .A1(MEM_stage_inst_dmem_n13171), .A2(MEM_stage_inst_dmem_n13170), .ZN(MEM_stage_inst_dmem_n12622) );
NAND2_X1 MEM_stage_inst_dmem_U9426 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n13177), .ZN(MEM_stage_inst_dmem_n13170) );
NAND2_X1 MEM_stage_inst_dmem_U9425 ( .A1(MEM_stage_inst_dmem_ram_275), .A2(MEM_stage_inst_dmem_n13176), .ZN(MEM_stage_inst_dmem_n13171) );
NAND2_X1 MEM_stage_inst_dmem_U9424 ( .A1(MEM_stage_inst_dmem_n13169), .A2(MEM_stage_inst_dmem_n13168), .ZN(MEM_stage_inst_dmem_n12623) );
NAND2_X1 MEM_stage_inst_dmem_U9423 ( .A1(MEM_stage_inst_dmem_n16368), .A2(MEM_stage_inst_dmem_n13177), .ZN(MEM_stage_inst_dmem_n13168) );
NAND2_X1 MEM_stage_inst_dmem_U9422 ( .A1(MEM_stage_inst_dmem_ram_276), .A2(MEM_stage_inst_dmem_n13176), .ZN(MEM_stage_inst_dmem_n13169) );
NAND2_X1 MEM_stage_inst_dmem_U9421 ( .A1(MEM_stage_inst_dmem_n13167), .A2(MEM_stage_inst_dmem_n13166), .ZN(MEM_stage_inst_dmem_n12624) );
NAND2_X1 MEM_stage_inst_dmem_U9420 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n13177), .ZN(MEM_stage_inst_dmem_n13166) );
NAND2_X1 MEM_stage_inst_dmem_U9419 ( .A1(MEM_stage_inst_dmem_ram_277), .A2(MEM_stage_inst_dmem_n13176), .ZN(MEM_stage_inst_dmem_n13167) );
NAND2_X1 MEM_stage_inst_dmem_U9418 ( .A1(MEM_stage_inst_dmem_n13165), .A2(MEM_stage_inst_dmem_n13164), .ZN(MEM_stage_inst_dmem_n12625) );
NAND2_X1 MEM_stage_inst_dmem_U9417 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n13177), .ZN(MEM_stage_inst_dmem_n13164) );
NAND2_X1 MEM_stage_inst_dmem_U9416 ( .A1(MEM_stage_inst_dmem_ram_278), .A2(MEM_stage_inst_dmem_n13176), .ZN(MEM_stage_inst_dmem_n13165) );
NAND2_X1 MEM_stage_inst_dmem_U9415 ( .A1(MEM_stage_inst_dmem_n13163), .A2(MEM_stage_inst_dmem_n13162), .ZN(MEM_stage_inst_dmem_n12626) );
NAND2_X1 MEM_stage_inst_dmem_U9414 ( .A1(MEM_stage_inst_dmem_n13886), .A2(MEM_stage_inst_dmem_n13177), .ZN(MEM_stage_inst_dmem_n13162) );
NAND2_X1 MEM_stage_inst_dmem_U9413 ( .A1(MEM_stage_inst_dmem_ram_279), .A2(MEM_stage_inst_dmem_n13176), .ZN(MEM_stage_inst_dmem_n13163) );
NAND2_X1 MEM_stage_inst_dmem_U9412 ( .A1(MEM_stage_inst_dmem_n13161), .A2(MEM_stage_inst_dmem_n13160), .ZN(MEM_stage_inst_dmem_n12627) );
NAND2_X1 MEM_stage_inst_dmem_U9411 ( .A1(MEM_stage_inst_dmem_n13883), .A2(MEM_stage_inst_dmem_n13177), .ZN(MEM_stage_inst_dmem_n13160) );
NAND2_X1 MEM_stage_inst_dmem_U9410 ( .A1(MEM_stage_inst_dmem_ram_280), .A2(MEM_stage_inst_dmem_n13176), .ZN(MEM_stage_inst_dmem_n13161) );
NAND2_X1 MEM_stage_inst_dmem_U9409 ( .A1(MEM_stage_inst_dmem_n13159), .A2(MEM_stage_inst_dmem_n13158), .ZN(MEM_stage_inst_dmem_n12628) );
NAND2_X1 MEM_stage_inst_dmem_U9408 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n13177), .ZN(MEM_stage_inst_dmem_n13158) );
NAND2_X1 MEM_stage_inst_dmem_U9407 ( .A1(MEM_stage_inst_dmem_ram_281), .A2(MEM_stage_inst_dmem_n13176), .ZN(MEM_stage_inst_dmem_n13159) );
NAND2_X1 MEM_stage_inst_dmem_U9406 ( .A1(MEM_stage_inst_dmem_n13157), .A2(MEM_stage_inst_dmem_n13156), .ZN(MEM_stage_inst_dmem_n12629) );
NAND2_X1 MEM_stage_inst_dmem_U9405 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n13177), .ZN(MEM_stage_inst_dmem_n13156) );
NAND2_X1 MEM_stage_inst_dmem_U9404 ( .A1(MEM_stage_inst_dmem_ram_282), .A2(MEM_stage_inst_dmem_n13176), .ZN(MEM_stage_inst_dmem_n13157) );
NAND2_X1 MEM_stage_inst_dmem_U9403 ( .A1(MEM_stage_inst_dmem_n13155), .A2(MEM_stage_inst_dmem_n13154), .ZN(MEM_stage_inst_dmem_n12630) );
NAND2_X1 MEM_stage_inst_dmem_U9402 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n13177), .ZN(MEM_stage_inst_dmem_n13154) );
NAND2_X1 MEM_stage_inst_dmem_U9401 ( .A1(MEM_stage_inst_dmem_ram_283), .A2(MEM_stage_inst_dmem_n13176), .ZN(MEM_stage_inst_dmem_n13155) );
NAND2_X1 MEM_stage_inst_dmem_U9400 ( .A1(MEM_stage_inst_dmem_n13153), .A2(MEM_stage_inst_dmem_n13152), .ZN(MEM_stage_inst_dmem_n12631) );
NAND2_X1 MEM_stage_inst_dmem_U9399 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n13177), .ZN(MEM_stage_inst_dmem_n13152) );
NAND2_X1 MEM_stage_inst_dmem_U9398 ( .A1(MEM_stage_inst_dmem_ram_284), .A2(MEM_stage_inst_dmem_n13176), .ZN(MEM_stage_inst_dmem_n13153) );
NAND2_X1 MEM_stage_inst_dmem_U9397 ( .A1(MEM_stage_inst_dmem_n13151), .A2(MEM_stage_inst_dmem_n13150), .ZN(MEM_stage_inst_dmem_n12632) );
NAND2_X1 MEM_stage_inst_dmem_U9396 ( .A1(MEM_stage_inst_dmem_n15116), .A2(MEM_stage_inst_dmem_n13177), .ZN(MEM_stage_inst_dmem_n13150) );
NAND2_X1 MEM_stage_inst_dmem_U9395 ( .A1(MEM_stage_inst_dmem_ram_285), .A2(MEM_stage_inst_dmem_n13176), .ZN(MEM_stage_inst_dmem_n13151) );
NAND2_X1 MEM_stage_inst_dmem_U9394 ( .A1(MEM_stage_inst_dmem_n13149), .A2(MEM_stage_inst_dmem_n13148), .ZN(MEM_stage_inst_dmem_n12633) );
NAND2_X1 MEM_stage_inst_dmem_U9393 ( .A1(MEM_stage_inst_dmem_n15113), .A2(MEM_stage_inst_dmem_n13177), .ZN(MEM_stage_inst_dmem_n13148) );
NAND2_X1 MEM_stage_inst_dmem_U9392 ( .A1(MEM_stage_inst_dmem_ram_286), .A2(MEM_stage_inst_dmem_n13176), .ZN(MEM_stage_inst_dmem_n13149) );
NAND2_X1 MEM_stage_inst_dmem_U9391 ( .A1(MEM_stage_inst_dmem_n13147), .A2(MEM_stage_inst_dmem_n13146), .ZN(MEM_stage_inst_dmem_n12634) );
NAND2_X1 MEM_stage_inst_dmem_U9390 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n13177), .ZN(MEM_stage_inst_dmem_n13146) );
NAND2_X1 MEM_stage_inst_dmem_U9389 ( .A1(MEM_stage_inst_dmem_ram_287), .A2(MEM_stage_inst_dmem_n13176), .ZN(MEM_stage_inst_dmem_n13147) );
NAND2_X1 MEM_stage_inst_dmem_U9388 ( .A1(MEM_stage_inst_dmem_n13182), .A2(MEM_stage_inst_dmem_n21429), .ZN(MEM_stage_inst_dmem_n13176) );
NOR2_X2 MEM_stage_inst_dmem_U9387 ( .A1(MEM_stage_inst_dmem_n13181), .A2(MEM_stage_inst_dmem_n13145), .ZN(MEM_stage_inst_dmem_n21429) );
NAND2_X1 MEM_stage_inst_dmem_U9386 ( .A1(MEM_stage_inst_dmem_n13144), .A2(MEM_stage_inst_dmem_n13143), .ZN(MEM_stage_inst_dmem_n12635) );
NAND2_X1 MEM_stage_inst_dmem_U9385 ( .A1(MEM_stage_inst_dmem_n14732), .A2(MEM_stage_inst_dmem_n13142), .ZN(MEM_stage_inst_dmem_n13143) );
NAND2_X1 MEM_stage_inst_dmem_U9384 ( .A1(MEM_stage_inst_dmem_ram_288), .A2(MEM_stage_inst_dmem_n13141), .ZN(MEM_stage_inst_dmem_n13144) );
NAND2_X1 MEM_stage_inst_dmem_U9383 ( .A1(MEM_stage_inst_dmem_n13140), .A2(MEM_stage_inst_dmem_n13139), .ZN(MEM_stage_inst_dmem_n12636) );
NAND2_X1 MEM_stage_inst_dmem_U9382 ( .A1(MEM_stage_inst_dmem_n15), .A2(MEM_stage_inst_dmem_n13142), .ZN(MEM_stage_inst_dmem_n13139) );
NAND2_X1 MEM_stage_inst_dmem_U9381 ( .A1(MEM_stage_inst_dmem_ram_289), .A2(MEM_stage_inst_dmem_n13141), .ZN(MEM_stage_inst_dmem_n13140) );
NAND2_X1 MEM_stage_inst_dmem_U9380 ( .A1(MEM_stage_inst_dmem_n13138), .A2(MEM_stage_inst_dmem_n13137), .ZN(MEM_stage_inst_dmem_n12637) );
NAND2_X1 MEM_stage_inst_dmem_U9379 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n13142), .ZN(MEM_stage_inst_dmem_n13137) );
NAND2_X1 MEM_stage_inst_dmem_U9378 ( .A1(MEM_stage_inst_dmem_ram_290), .A2(MEM_stage_inst_dmem_n13141), .ZN(MEM_stage_inst_dmem_n13138) );
NAND2_X1 MEM_stage_inst_dmem_U9377 ( .A1(MEM_stage_inst_dmem_n13136), .A2(MEM_stage_inst_dmem_n13135), .ZN(MEM_stage_inst_dmem_n12638) );
NAND2_X1 MEM_stage_inst_dmem_U9376 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n13142), .ZN(MEM_stage_inst_dmem_n13135) );
NAND2_X1 MEM_stage_inst_dmem_U9375 ( .A1(MEM_stage_inst_dmem_ram_291), .A2(MEM_stage_inst_dmem_n13141), .ZN(MEM_stage_inst_dmem_n13136) );
NAND2_X1 MEM_stage_inst_dmem_U9374 ( .A1(MEM_stage_inst_dmem_n13134), .A2(MEM_stage_inst_dmem_n13133), .ZN(MEM_stage_inst_dmem_n12639) );
NAND2_X1 MEM_stage_inst_dmem_U9373 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n13142), .ZN(MEM_stage_inst_dmem_n13133) );
NAND2_X1 MEM_stage_inst_dmem_U9372 ( .A1(MEM_stage_inst_dmem_ram_292), .A2(MEM_stage_inst_dmem_n13141), .ZN(MEM_stage_inst_dmem_n13134) );
NAND2_X1 MEM_stage_inst_dmem_U9371 ( .A1(MEM_stage_inst_dmem_n13132), .A2(MEM_stage_inst_dmem_n13131), .ZN(MEM_stage_inst_dmem_n12640) );
NAND2_X1 MEM_stage_inst_dmem_U9370 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n13142), .ZN(MEM_stage_inst_dmem_n13131) );
NAND2_X1 MEM_stage_inst_dmem_U9369 ( .A1(MEM_stage_inst_dmem_ram_293), .A2(MEM_stage_inst_dmem_n13141), .ZN(MEM_stage_inst_dmem_n13132) );
NAND2_X1 MEM_stage_inst_dmem_U9368 ( .A1(MEM_stage_inst_dmem_n13130), .A2(MEM_stage_inst_dmem_n13129), .ZN(MEM_stage_inst_dmem_n12641) );
NAND2_X1 MEM_stage_inst_dmem_U9367 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n13142), .ZN(MEM_stage_inst_dmem_n13129) );
NAND2_X1 MEM_stage_inst_dmem_U9366 ( .A1(MEM_stage_inst_dmem_ram_294), .A2(MEM_stage_inst_dmem_n13141), .ZN(MEM_stage_inst_dmem_n13130) );
NAND2_X1 MEM_stage_inst_dmem_U9365 ( .A1(MEM_stage_inst_dmem_n13128), .A2(MEM_stage_inst_dmem_n13127), .ZN(MEM_stage_inst_dmem_n12642) );
NAND2_X1 MEM_stage_inst_dmem_U9364 ( .A1(MEM_stage_inst_dmem_n18), .A2(MEM_stage_inst_dmem_n13142), .ZN(MEM_stage_inst_dmem_n13127) );
NAND2_X1 MEM_stage_inst_dmem_U9363 ( .A1(MEM_stage_inst_dmem_ram_295), .A2(MEM_stage_inst_dmem_n13141), .ZN(MEM_stage_inst_dmem_n13128) );
NAND2_X1 MEM_stage_inst_dmem_U9362 ( .A1(MEM_stage_inst_dmem_n13126), .A2(MEM_stage_inst_dmem_n13125), .ZN(MEM_stage_inst_dmem_n12643) );
NAND2_X1 MEM_stage_inst_dmem_U9361 ( .A1(MEM_stage_inst_dmem_n4), .A2(MEM_stage_inst_dmem_n13142), .ZN(MEM_stage_inst_dmem_n13125) );
NAND2_X1 MEM_stage_inst_dmem_U9360 ( .A1(MEM_stage_inst_dmem_ram_296), .A2(MEM_stage_inst_dmem_n13141), .ZN(MEM_stage_inst_dmem_n13126) );
NAND2_X1 MEM_stage_inst_dmem_U9359 ( .A1(MEM_stage_inst_dmem_n13124), .A2(MEM_stage_inst_dmem_n13123), .ZN(MEM_stage_inst_dmem_n12644) );
NAND2_X1 MEM_stage_inst_dmem_U9358 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n13142), .ZN(MEM_stage_inst_dmem_n13123) );
NAND2_X1 MEM_stage_inst_dmem_U9357 ( .A1(MEM_stage_inst_dmem_ram_297), .A2(MEM_stage_inst_dmem_n13141), .ZN(MEM_stage_inst_dmem_n13124) );
NAND2_X1 MEM_stage_inst_dmem_U9356 ( .A1(MEM_stage_inst_dmem_n13122), .A2(MEM_stage_inst_dmem_n13121), .ZN(MEM_stage_inst_dmem_n12645) );
NAND2_X1 MEM_stage_inst_dmem_U9355 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n13142), .ZN(MEM_stage_inst_dmem_n13121) );
NAND2_X1 MEM_stage_inst_dmem_U9354 ( .A1(MEM_stage_inst_dmem_ram_298), .A2(MEM_stage_inst_dmem_n13141), .ZN(MEM_stage_inst_dmem_n13122) );
NAND2_X1 MEM_stage_inst_dmem_U9353 ( .A1(MEM_stage_inst_dmem_n13120), .A2(MEM_stage_inst_dmem_n13119), .ZN(MEM_stage_inst_dmem_n12646) );
NAND2_X1 MEM_stage_inst_dmem_U9352 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n13142), .ZN(MEM_stage_inst_dmem_n13119) );
NAND2_X1 MEM_stage_inst_dmem_U9351 ( .A1(MEM_stage_inst_dmem_ram_299), .A2(MEM_stage_inst_dmem_n13141), .ZN(MEM_stage_inst_dmem_n13120) );
NAND2_X1 MEM_stage_inst_dmem_U9350 ( .A1(MEM_stage_inst_dmem_n13118), .A2(MEM_stage_inst_dmem_n13117), .ZN(MEM_stage_inst_dmem_n12647) );
NAND2_X1 MEM_stage_inst_dmem_U9349 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n13142), .ZN(MEM_stage_inst_dmem_n13117) );
NAND2_X1 MEM_stage_inst_dmem_U9348 ( .A1(MEM_stage_inst_dmem_ram_300), .A2(MEM_stage_inst_dmem_n13141), .ZN(MEM_stage_inst_dmem_n13118) );
NAND2_X1 MEM_stage_inst_dmem_U9347 ( .A1(MEM_stage_inst_dmem_n13116), .A2(MEM_stage_inst_dmem_n13115), .ZN(MEM_stage_inst_dmem_n12648) );
NAND2_X1 MEM_stage_inst_dmem_U9346 ( .A1(MEM_stage_inst_dmem_n116), .A2(MEM_stage_inst_dmem_n13142), .ZN(MEM_stage_inst_dmem_n13115) );
NAND2_X1 MEM_stage_inst_dmem_U9345 ( .A1(MEM_stage_inst_dmem_ram_301), .A2(MEM_stage_inst_dmem_n13141), .ZN(MEM_stage_inst_dmem_n13116) );
NAND2_X1 MEM_stage_inst_dmem_U9344 ( .A1(MEM_stage_inst_dmem_n13114), .A2(MEM_stage_inst_dmem_n13113), .ZN(MEM_stage_inst_dmem_n12649) );
NAND2_X1 MEM_stage_inst_dmem_U9343 ( .A1(MEM_stage_inst_dmem_n14696), .A2(MEM_stage_inst_dmem_n13142), .ZN(MEM_stage_inst_dmem_n13113) );
NAND2_X1 MEM_stage_inst_dmem_U9342 ( .A1(MEM_stage_inst_dmem_ram_302), .A2(MEM_stage_inst_dmem_n13141), .ZN(MEM_stage_inst_dmem_n13114) );
NAND2_X1 MEM_stage_inst_dmem_U9341 ( .A1(MEM_stage_inst_dmem_n13112), .A2(MEM_stage_inst_dmem_n13111), .ZN(MEM_stage_inst_dmem_n12650) );
NAND2_X1 MEM_stage_inst_dmem_U9340 ( .A1(MEM_stage_inst_dmem_n14693), .A2(MEM_stage_inst_dmem_n13142), .ZN(MEM_stage_inst_dmem_n13111) );
INV_X1 MEM_stage_inst_dmem_U9339 ( .A(MEM_stage_inst_dmem_n13141), .ZN(MEM_stage_inst_dmem_n13142) );
NAND2_X1 MEM_stage_inst_dmem_U9338 ( .A1(MEM_stage_inst_dmem_ram_303), .A2(MEM_stage_inst_dmem_n13141), .ZN(MEM_stage_inst_dmem_n13112) );
NAND2_X1 MEM_stage_inst_dmem_U9337 ( .A1(MEM_stage_inst_dmem_n13182), .A2(MEM_stage_inst_dmem_n21394), .ZN(MEM_stage_inst_dmem_n13141) );
NOR2_X2 MEM_stage_inst_dmem_U9336 ( .A1(MEM_stage_inst_dmem_n13110), .A2(MEM_stage_inst_dmem_n13180), .ZN(MEM_stage_inst_dmem_n21394) );
NAND2_X1 MEM_stage_inst_dmem_U9335 ( .A1(MEM_stage_inst_dmem_n13109), .A2(MEM_stage_inst_dmem_n13108), .ZN(MEM_stage_inst_dmem_n12651) );
NAND2_X1 MEM_stage_inst_dmem_U9334 ( .A1(MEM_stage_inst_dmem_n14732), .A2(MEM_stage_inst_dmem_n13107), .ZN(MEM_stage_inst_dmem_n13108) );
NAND2_X1 MEM_stage_inst_dmem_U9333 ( .A1(MEM_stage_inst_dmem_ram_304), .A2(MEM_stage_inst_dmem_n13106), .ZN(MEM_stage_inst_dmem_n13109) );
NAND2_X1 MEM_stage_inst_dmem_U9332 ( .A1(MEM_stage_inst_dmem_n13105), .A2(MEM_stage_inst_dmem_n13104), .ZN(MEM_stage_inst_dmem_n12652) );
NAND2_X1 MEM_stage_inst_dmem_U9331 ( .A1(MEM_stage_inst_dmem_n14), .A2(MEM_stage_inst_dmem_n13107), .ZN(MEM_stage_inst_dmem_n13104) );
NAND2_X1 MEM_stage_inst_dmem_U9330 ( .A1(MEM_stage_inst_dmem_ram_305), .A2(MEM_stage_inst_dmem_n13106), .ZN(MEM_stage_inst_dmem_n13105) );
NAND2_X1 MEM_stage_inst_dmem_U9329 ( .A1(MEM_stage_inst_dmem_n13103), .A2(MEM_stage_inst_dmem_n13102), .ZN(MEM_stage_inst_dmem_n12653) );
NAND2_X1 MEM_stage_inst_dmem_U9328 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n13107), .ZN(MEM_stage_inst_dmem_n13102) );
NAND2_X1 MEM_stage_inst_dmem_U9327 ( .A1(MEM_stage_inst_dmem_ram_306), .A2(MEM_stage_inst_dmem_n13106), .ZN(MEM_stage_inst_dmem_n13103) );
NAND2_X1 MEM_stage_inst_dmem_U9326 ( .A1(MEM_stage_inst_dmem_n13101), .A2(MEM_stage_inst_dmem_n13100), .ZN(MEM_stage_inst_dmem_n12654) );
NAND2_X1 MEM_stage_inst_dmem_U9325 ( .A1(MEM_stage_inst_dmem_n13897), .A2(MEM_stage_inst_dmem_n13107), .ZN(MEM_stage_inst_dmem_n13100) );
NAND2_X1 MEM_stage_inst_dmem_U9324 ( .A1(MEM_stage_inst_dmem_ram_307), .A2(MEM_stage_inst_dmem_n13106), .ZN(MEM_stage_inst_dmem_n13101) );
NAND2_X1 MEM_stage_inst_dmem_U9323 ( .A1(MEM_stage_inst_dmem_n13099), .A2(MEM_stage_inst_dmem_n13098), .ZN(MEM_stage_inst_dmem_n12655) );
NAND2_X1 MEM_stage_inst_dmem_U9322 ( .A1(MEM_stage_inst_dmem_n16368), .A2(MEM_stage_inst_dmem_n13107), .ZN(MEM_stage_inst_dmem_n13098) );
NAND2_X1 MEM_stage_inst_dmem_U9321 ( .A1(MEM_stage_inst_dmem_ram_308), .A2(MEM_stage_inst_dmem_n13106), .ZN(MEM_stage_inst_dmem_n13099) );
NAND2_X1 MEM_stage_inst_dmem_U9320 ( .A1(MEM_stage_inst_dmem_n13097), .A2(MEM_stage_inst_dmem_n13096), .ZN(MEM_stage_inst_dmem_n12656) );
NAND2_X1 MEM_stage_inst_dmem_U9319 ( .A1(MEM_stage_inst_dmem_n13892), .A2(MEM_stage_inst_dmem_n13107), .ZN(MEM_stage_inst_dmem_n13096) );
NAND2_X1 MEM_stage_inst_dmem_U9318 ( .A1(MEM_stage_inst_dmem_ram_309), .A2(MEM_stage_inst_dmem_n13106), .ZN(MEM_stage_inst_dmem_n13097) );
NAND2_X1 MEM_stage_inst_dmem_U9317 ( .A1(MEM_stage_inst_dmem_n13095), .A2(MEM_stage_inst_dmem_n13094), .ZN(MEM_stage_inst_dmem_n12657) );
NAND2_X1 MEM_stage_inst_dmem_U9316 ( .A1(MEM_stage_inst_dmem_n13889), .A2(MEM_stage_inst_dmem_n13107), .ZN(MEM_stage_inst_dmem_n13094) );
NAND2_X1 MEM_stage_inst_dmem_U9315 ( .A1(MEM_stage_inst_dmem_ram_310), .A2(MEM_stage_inst_dmem_n13106), .ZN(MEM_stage_inst_dmem_n13095) );
NAND2_X1 MEM_stage_inst_dmem_U9314 ( .A1(MEM_stage_inst_dmem_n13093), .A2(MEM_stage_inst_dmem_n13092), .ZN(MEM_stage_inst_dmem_n12658) );
NAND2_X1 MEM_stage_inst_dmem_U9313 ( .A1(MEM_stage_inst_dmem_n13886), .A2(MEM_stage_inst_dmem_n13107), .ZN(MEM_stage_inst_dmem_n13092) );
BUF_X1 MEM_stage_inst_dmem_U9312 ( .A(EX_pipeline_reg_out_12), .Z(MEM_stage_inst_dmem_n13886) );
NAND2_X1 MEM_stage_inst_dmem_U9311 ( .A1(MEM_stage_inst_dmem_ram_311), .A2(MEM_stage_inst_dmem_n13106), .ZN(MEM_stage_inst_dmem_n13093) );
NAND2_X1 MEM_stage_inst_dmem_U9310 ( .A1(MEM_stage_inst_dmem_n13091), .A2(MEM_stage_inst_dmem_n13090), .ZN(MEM_stage_inst_dmem_n12659) );
NAND2_X1 MEM_stage_inst_dmem_U9309 ( .A1(MEM_stage_inst_dmem_n13883), .A2(MEM_stage_inst_dmem_n13107), .ZN(MEM_stage_inst_dmem_n13090) );
BUF_X1 MEM_stage_inst_dmem_U9308 ( .A(EX_pipeline_reg_out_13), .Z(MEM_stage_inst_dmem_n13883) );
NAND2_X1 MEM_stage_inst_dmem_U9307 ( .A1(MEM_stage_inst_dmem_ram_312), .A2(MEM_stage_inst_dmem_n13106), .ZN(MEM_stage_inst_dmem_n13091) );
NAND2_X1 MEM_stage_inst_dmem_U9306 ( .A1(MEM_stage_inst_dmem_n13089), .A2(MEM_stage_inst_dmem_n13088), .ZN(MEM_stage_inst_dmem_n12660) );
NAND2_X1 MEM_stage_inst_dmem_U9305 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n13107), .ZN(MEM_stage_inst_dmem_n13088) );
NAND2_X1 MEM_stage_inst_dmem_U9304 ( .A1(MEM_stage_inst_dmem_ram_313), .A2(MEM_stage_inst_dmem_n13106), .ZN(MEM_stage_inst_dmem_n13089) );
NAND2_X1 MEM_stage_inst_dmem_U9303 ( .A1(MEM_stage_inst_dmem_n13087), .A2(MEM_stage_inst_dmem_n13086), .ZN(MEM_stage_inst_dmem_n12661) );
NAND2_X1 MEM_stage_inst_dmem_U9302 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n13107), .ZN(MEM_stage_inst_dmem_n13086) );
NAND2_X1 MEM_stage_inst_dmem_U9301 ( .A1(MEM_stage_inst_dmem_ram_314), .A2(MEM_stage_inst_dmem_n13106), .ZN(MEM_stage_inst_dmem_n13087) );
NAND2_X1 MEM_stage_inst_dmem_U9300 ( .A1(MEM_stage_inst_dmem_n13085), .A2(MEM_stage_inst_dmem_n13084), .ZN(MEM_stage_inst_dmem_n12662) );
NAND2_X1 MEM_stage_inst_dmem_U9299 ( .A1(MEM_stage_inst_dmem_n13874), .A2(MEM_stage_inst_dmem_n13107), .ZN(MEM_stage_inst_dmem_n13084) );
NAND2_X1 MEM_stage_inst_dmem_U9298 ( .A1(MEM_stage_inst_dmem_ram_315), .A2(MEM_stage_inst_dmem_n13106), .ZN(MEM_stage_inst_dmem_n13085) );
NAND2_X1 MEM_stage_inst_dmem_U9297 ( .A1(MEM_stage_inst_dmem_n13083), .A2(MEM_stage_inst_dmem_n13082), .ZN(MEM_stage_inst_dmem_n12663) );
NAND2_X1 MEM_stage_inst_dmem_U9296 ( .A1(MEM_stage_inst_dmem_n13871), .A2(MEM_stage_inst_dmem_n13107), .ZN(MEM_stage_inst_dmem_n13082) );
NAND2_X1 MEM_stage_inst_dmem_U9295 ( .A1(MEM_stage_inst_dmem_ram_316), .A2(MEM_stage_inst_dmem_n13106), .ZN(MEM_stage_inst_dmem_n13083) );
NAND2_X1 MEM_stage_inst_dmem_U9294 ( .A1(MEM_stage_inst_dmem_n13081), .A2(MEM_stage_inst_dmem_n13080), .ZN(MEM_stage_inst_dmem_n12664) );
NAND2_X1 MEM_stage_inst_dmem_U9293 ( .A1(MEM_stage_inst_dmem_n116), .A2(MEM_stage_inst_dmem_n13107), .ZN(MEM_stage_inst_dmem_n13080) );
NAND2_X1 MEM_stage_inst_dmem_U9292 ( .A1(MEM_stage_inst_dmem_ram_317), .A2(MEM_stage_inst_dmem_n13106), .ZN(MEM_stage_inst_dmem_n13081) );
NAND2_X1 MEM_stage_inst_dmem_U9291 ( .A1(MEM_stage_inst_dmem_n13079), .A2(MEM_stage_inst_dmem_n13078), .ZN(MEM_stage_inst_dmem_n12665) );
NAND2_X1 MEM_stage_inst_dmem_U9290 ( .A1(MEM_stage_inst_dmem_n14696), .A2(MEM_stage_inst_dmem_n13107), .ZN(MEM_stage_inst_dmem_n13078) );
NAND2_X1 MEM_stage_inst_dmem_U9289 ( .A1(MEM_stage_inst_dmem_ram_318), .A2(MEM_stage_inst_dmem_n13106), .ZN(MEM_stage_inst_dmem_n13079) );
NAND2_X1 MEM_stage_inst_dmem_U9288 ( .A1(MEM_stage_inst_dmem_n13077), .A2(MEM_stage_inst_dmem_n13076), .ZN(MEM_stage_inst_dmem_n12666) );
NAND2_X1 MEM_stage_inst_dmem_U9287 ( .A1(MEM_stage_inst_dmem_n15110), .A2(MEM_stage_inst_dmem_n13107), .ZN(MEM_stage_inst_dmem_n13076) );
NAND2_X1 MEM_stage_inst_dmem_U9286 ( .A1(MEM_stage_inst_dmem_ram_319), .A2(MEM_stage_inst_dmem_n13106), .ZN(MEM_stage_inst_dmem_n13077) );
NAND2_X1 MEM_stage_inst_dmem_U9285 ( .A1(MEM_stage_inst_dmem_n13182), .A2(MEM_stage_inst_dmem_n21359), .ZN(MEM_stage_inst_dmem_n13106) );
NOR2_X2 MEM_stage_inst_dmem_U9284 ( .A1(MEM_stage_inst_dmem_n13110), .A2(MEM_stage_inst_dmem_n13145), .ZN(MEM_stage_inst_dmem_n21359) );
NAND2_X1 MEM_stage_inst_dmem_U9283 ( .A1(MEM_stage_inst_dmem_n13075), .A2(MEM_stage_inst_dmem_n13074), .ZN(MEM_stage_inst_dmem_n12667) );
NAND2_X1 MEM_stage_inst_dmem_U9282 ( .A1(MEM_stage_inst_dmem_n14732), .A2(MEM_stage_inst_dmem_n13073), .ZN(MEM_stage_inst_dmem_n13074) );
NAND2_X1 MEM_stage_inst_dmem_U9281 ( .A1(MEM_stage_inst_dmem_ram_320), .A2(MEM_stage_inst_dmem_n13072), .ZN(MEM_stage_inst_dmem_n13075) );
NAND2_X1 MEM_stage_inst_dmem_U9280 ( .A1(MEM_stage_inst_dmem_n13071), .A2(MEM_stage_inst_dmem_n13070), .ZN(MEM_stage_inst_dmem_n12668) );
NAND2_X1 MEM_stage_inst_dmem_U9279 ( .A1(EX_pipeline_reg_out_6), .A2(MEM_stage_inst_dmem_n13073), .ZN(MEM_stage_inst_dmem_n13070) );
NAND2_X1 MEM_stage_inst_dmem_U9278 ( .A1(MEM_stage_inst_dmem_ram_321), .A2(MEM_stage_inst_dmem_n13072), .ZN(MEM_stage_inst_dmem_n13071) );
NAND2_X1 MEM_stage_inst_dmem_U9277 ( .A1(MEM_stage_inst_dmem_n13068), .A2(MEM_stage_inst_dmem_n13067), .ZN(MEM_stage_inst_dmem_n12669) );
NAND2_X1 MEM_stage_inst_dmem_U9276 ( .A1(EX_pipeline_reg_out_7), .A2(MEM_stage_inst_dmem_n13073), .ZN(MEM_stage_inst_dmem_n13067) );
NAND2_X1 MEM_stage_inst_dmem_U9275 ( .A1(MEM_stage_inst_dmem_ram_322), .A2(MEM_stage_inst_dmem_n13072), .ZN(MEM_stage_inst_dmem_n13068) );
NAND2_X1 MEM_stage_inst_dmem_U9274 ( .A1(MEM_stage_inst_dmem_n13066), .A2(MEM_stage_inst_dmem_n13065), .ZN(MEM_stage_inst_dmem_n12670) );
NAND2_X1 MEM_stage_inst_dmem_U9273 ( .A1(MEM_stage_inst_dmem_n13064), .A2(MEM_stage_inst_dmem_n13073), .ZN(MEM_stage_inst_dmem_n13065) );
NAND2_X1 MEM_stage_inst_dmem_U9272 ( .A1(MEM_stage_inst_dmem_ram_323), .A2(MEM_stage_inst_dmem_n13072), .ZN(MEM_stage_inst_dmem_n13066) );
NAND2_X1 MEM_stage_inst_dmem_U9271 ( .A1(MEM_stage_inst_dmem_n13063), .A2(MEM_stage_inst_dmem_n13062), .ZN(MEM_stage_inst_dmem_n12671) );
NAND2_X1 MEM_stage_inst_dmem_U9270 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n13073), .ZN(MEM_stage_inst_dmem_n13062) );
NAND2_X1 MEM_stage_inst_dmem_U9269 ( .A1(MEM_stage_inst_dmem_ram_324), .A2(MEM_stage_inst_dmem_n13072), .ZN(MEM_stage_inst_dmem_n13063) );
NAND2_X1 MEM_stage_inst_dmem_U9268 ( .A1(MEM_stage_inst_dmem_n13061), .A2(MEM_stage_inst_dmem_n13060), .ZN(MEM_stage_inst_dmem_n12672) );
NAND2_X1 MEM_stage_inst_dmem_U9267 ( .A1(MEM_stage_inst_dmem_n13059), .A2(MEM_stage_inst_dmem_n13073), .ZN(MEM_stage_inst_dmem_n13060) );
NAND2_X1 MEM_stage_inst_dmem_U9266 ( .A1(MEM_stage_inst_dmem_ram_325), .A2(MEM_stage_inst_dmem_n13072), .ZN(MEM_stage_inst_dmem_n13061) );
NAND2_X1 MEM_stage_inst_dmem_U9265 ( .A1(MEM_stage_inst_dmem_n13058), .A2(MEM_stage_inst_dmem_n13057), .ZN(MEM_stage_inst_dmem_n12673) );
NAND2_X1 MEM_stage_inst_dmem_U9264 ( .A1(MEM_stage_inst_dmem_n13056), .A2(MEM_stage_inst_dmem_n13073), .ZN(MEM_stage_inst_dmem_n13057) );
NAND2_X1 MEM_stage_inst_dmem_U9263 ( .A1(MEM_stage_inst_dmem_ram_326), .A2(MEM_stage_inst_dmem_n13072), .ZN(MEM_stage_inst_dmem_n13058) );
NAND2_X1 MEM_stage_inst_dmem_U9262 ( .A1(MEM_stage_inst_dmem_n13055), .A2(MEM_stage_inst_dmem_n13054), .ZN(MEM_stage_inst_dmem_n12674) );
NAND2_X1 MEM_stage_inst_dmem_U9261 ( .A1(MEM_stage_inst_dmem_n112), .A2(MEM_stage_inst_dmem_n13073), .ZN(MEM_stage_inst_dmem_n13054) );
NAND2_X1 MEM_stage_inst_dmem_U9260 ( .A1(MEM_stage_inst_dmem_ram_327), .A2(MEM_stage_inst_dmem_n13072), .ZN(MEM_stage_inst_dmem_n13055) );
NAND2_X1 MEM_stage_inst_dmem_U9259 ( .A1(MEM_stage_inst_dmem_n13053), .A2(MEM_stage_inst_dmem_n13052), .ZN(MEM_stage_inst_dmem_n12675) );
NAND2_X1 MEM_stage_inst_dmem_U9258 ( .A1(MEM_stage_inst_dmem_n13051), .A2(MEM_stage_inst_dmem_n13073), .ZN(MEM_stage_inst_dmem_n13052) );
NAND2_X1 MEM_stage_inst_dmem_U9257 ( .A1(MEM_stage_inst_dmem_ram_328), .A2(MEM_stage_inst_dmem_n13072), .ZN(MEM_stage_inst_dmem_n13053) );
NAND2_X1 MEM_stage_inst_dmem_U9256 ( .A1(MEM_stage_inst_dmem_n13050), .A2(MEM_stage_inst_dmem_n13049), .ZN(MEM_stage_inst_dmem_n12676) );
NAND2_X1 MEM_stage_inst_dmem_U9255 ( .A1(EX_pipeline_reg_out_14), .A2(MEM_stage_inst_dmem_n13073), .ZN(MEM_stage_inst_dmem_n13049) );
NAND2_X1 MEM_stage_inst_dmem_U9254 ( .A1(MEM_stage_inst_dmem_ram_329), .A2(MEM_stage_inst_dmem_n13072), .ZN(MEM_stage_inst_dmem_n13050) );
NAND2_X1 MEM_stage_inst_dmem_U9253 ( .A1(MEM_stage_inst_dmem_n13048), .A2(MEM_stage_inst_dmem_n13047), .ZN(MEM_stage_inst_dmem_n12677) );
NAND2_X1 MEM_stage_inst_dmem_U9252 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n13073), .ZN(MEM_stage_inst_dmem_n13047) );
NAND2_X1 MEM_stage_inst_dmem_U9251 ( .A1(MEM_stage_inst_dmem_ram_330), .A2(MEM_stage_inst_dmem_n13072), .ZN(MEM_stage_inst_dmem_n13048) );
NAND2_X1 MEM_stage_inst_dmem_U9250 ( .A1(MEM_stage_inst_dmem_n13046), .A2(MEM_stage_inst_dmem_n13045), .ZN(MEM_stage_inst_dmem_n12678) );
NAND2_X1 MEM_stage_inst_dmem_U9249 ( .A1(MEM_stage_inst_dmem_n13044), .A2(MEM_stage_inst_dmem_n13073), .ZN(MEM_stage_inst_dmem_n13045) );
NAND2_X1 MEM_stage_inst_dmem_U9248 ( .A1(MEM_stage_inst_dmem_ram_331), .A2(MEM_stage_inst_dmem_n13072), .ZN(MEM_stage_inst_dmem_n13046) );
NAND2_X1 MEM_stage_inst_dmem_U9247 ( .A1(MEM_stage_inst_dmem_n13043), .A2(MEM_stage_inst_dmem_n13042), .ZN(MEM_stage_inst_dmem_n12679) );
NAND2_X1 MEM_stage_inst_dmem_U9246 ( .A1(MEM_stage_inst_dmem_n13041), .A2(MEM_stage_inst_dmem_n13073), .ZN(MEM_stage_inst_dmem_n13042) );
NAND2_X1 MEM_stage_inst_dmem_U9245 ( .A1(MEM_stage_inst_dmem_ram_332), .A2(MEM_stage_inst_dmem_n13072), .ZN(MEM_stage_inst_dmem_n13043) );
NAND2_X1 MEM_stage_inst_dmem_U9244 ( .A1(MEM_stage_inst_dmem_n13040), .A2(MEM_stage_inst_dmem_n13039), .ZN(MEM_stage_inst_dmem_n12680) );
NAND2_X1 MEM_stage_inst_dmem_U9243 ( .A1(MEM_stage_inst_dmem_n116), .A2(MEM_stage_inst_dmem_n13073), .ZN(MEM_stage_inst_dmem_n13039) );
NAND2_X1 MEM_stage_inst_dmem_U9242 ( .A1(MEM_stage_inst_dmem_ram_333), .A2(MEM_stage_inst_dmem_n13072), .ZN(MEM_stage_inst_dmem_n13040) );
NAND2_X1 MEM_stage_inst_dmem_U9241 ( .A1(MEM_stage_inst_dmem_n13038), .A2(MEM_stage_inst_dmem_n13037), .ZN(MEM_stage_inst_dmem_n12681) );
NAND2_X1 MEM_stage_inst_dmem_U9240 ( .A1(MEM_stage_inst_dmem_n14696), .A2(MEM_stage_inst_dmem_n13073), .ZN(MEM_stage_inst_dmem_n13037) );
NAND2_X1 MEM_stage_inst_dmem_U9239 ( .A1(MEM_stage_inst_dmem_ram_334), .A2(MEM_stage_inst_dmem_n13072), .ZN(MEM_stage_inst_dmem_n13038) );
NAND2_X1 MEM_stage_inst_dmem_U9238 ( .A1(MEM_stage_inst_dmem_n13036), .A2(MEM_stage_inst_dmem_n13035), .ZN(MEM_stage_inst_dmem_n12682) );
NAND2_X1 MEM_stage_inst_dmem_U9237 ( .A1(MEM_stage_inst_dmem_n14693), .A2(MEM_stage_inst_dmem_n13073), .ZN(MEM_stage_inst_dmem_n13035) );
INV_X1 MEM_stage_inst_dmem_U9236 ( .A(MEM_stage_inst_dmem_n13072), .ZN(MEM_stage_inst_dmem_n13073) );
NAND2_X1 MEM_stage_inst_dmem_U9235 ( .A1(MEM_stage_inst_dmem_ram_335), .A2(MEM_stage_inst_dmem_n13072), .ZN(MEM_stage_inst_dmem_n13036) );
NAND2_X1 MEM_stage_inst_dmem_U9234 ( .A1(MEM_stage_inst_dmem_n13182), .A2(MEM_stage_inst_dmem_n21319), .ZN(MEM_stage_inst_dmem_n13072) );
NOR2_X2 MEM_stage_inst_dmem_U9233 ( .A1(MEM_stage_inst_dmem_n13034), .A2(MEM_stage_inst_dmem_n13180), .ZN(MEM_stage_inst_dmem_n21319) );
NAND2_X1 MEM_stage_inst_dmem_U9232 ( .A1(MEM_stage_inst_dmem_n13033), .A2(MEM_stage_inst_dmem_n13032), .ZN(MEM_stage_inst_dmem_n12683) );
NAND2_X1 MEM_stage_inst_dmem_U9231 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n13031), .ZN(MEM_stage_inst_dmem_n13032) );
NAND2_X1 MEM_stage_inst_dmem_U9230 ( .A1(MEM_stage_inst_dmem_ram_336), .A2(MEM_stage_inst_dmem_n13030), .ZN(MEM_stage_inst_dmem_n13033) );
NAND2_X1 MEM_stage_inst_dmem_U9229 ( .A1(MEM_stage_inst_dmem_n13029), .A2(MEM_stage_inst_dmem_n13028), .ZN(MEM_stage_inst_dmem_n12684) );
NAND2_X1 MEM_stage_inst_dmem_U9228 ( .A1(MEM_stage_inst_dmem_n109), .A2(MEM_stage_inst_dmem_n13031), .ZN(MEM_stage_inst_dmem_n13028) );
NAND2_X1 MEM_stage_inst_dmem_U9227 ( .A1(MEM_stage_inst_dmem_ram_337), .A2(MEM_stage_inst_dmem_n13030), .ZN(MEM_stage_inst_dmem_n13029) );
NAND2_X1 MEM_stage_inst_dmem_U9226 ( .A1(MEM_stage_inst_dmem_n13027), .A2(MEM_stage_inst_dmem_n13026), .ZN(MEM_stage_inst_dmem_n12685) );
NAND2_X1 MEM_stage_inst_dmem_U9225 ( .A1(MEM_stage_inst_dmem_n20544), .A2(MEM_stage_inst_dmem_n13031), .ZN(MEM_stage_inst_dmem_n13026) );
NAND2_X1 MEM_stage_inst_dmem_U9224 ( .A1(MEM_stage_inst_dmem_ram_338), .A2(MEM_stage_inst_dmem_n13030), .ZN(MEM_stage_inst_dmem_n13027) );
NAND2_X1 MEM_stage_inst_dmem_U9223 ( .A1(MEM_stage_inst_dmem_n13025), .A2(MEM_stage_inst_dmem_n13024), .ZN(MEM_stage_inst_dmem_n12686) );
NAND2_X1 MEM_stage_inst_dmem_U9222 ( .A1(MEM_stage_inst_dmem_n13064), .A2(MEM_stage_inst_dmem_n13031), .ZN(MEM_stage_inst_dmem_n13024) );
NAND2_X1 MEM_stage_inst_dmem_U9221 ( .A1(MEM_stage_inst_dmem_ram_339), .A2(MEM_stage_inst_dmem_n13030), .ZN(MEM_stage_inst_dmem_n13025) );
NAND2_X1 MEM_stage_inst_dmem_U9220 ( .A1(MEM_stage_inst_dmem_n13023), .A2(MEM_stage_inst_dmem_n13022), .ZN(MEM_stage_inst_dmem_n12687) );
NAND2_X1 MEM_stage_inst_dmem_U9219 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n13031), .ZN(MEM_stage_inst_dmem_n13022) );
NAND2_X1 MEM_stage_inst_dmem_U9218 ( .A1(MEM_stage_inst_dmem_ram_340), .A2(MEM_stage_inst_dmem_n13030), .ZN(MEM_stage_inst_dmem_n13023) );
NAND2_X1 MEM_stage_inst_dmem_U9217 ( .A1(MEM_stage_inst_dmem_n13021), .A2(MEM_stage_inst_dmem_n13020), .ZN(MEM_stage_inst_dmem_n12688) );
NAND2_X1 MEM_stage_inst_dmem_U9216 ( .A1(MEM_stage_inst_dmem_n13059), .A2(MEM_stage_inst_dmem_n13031), .ZN(MEM_stage_inst_dmem_n13020) );
NAND2_X1 MEM_stage_inst_dmem_U9215 ( .A1(MEM_stage_inst_dmem_ram_341), .A2(MEM_stage_inst_dmem_n13030), .ZN(MEM_stage_inst_dmem_n13021) );
NAND2_X1 MEM_stage_inst_dmem_U9214 ( .A1(MEM_stage_inst_dmem_n13019), .A2(MEM_stage_inst_dmem_n13018), .ZN(MEM_stage_inst_dmem_n12689) );
NAND2_X1 MEM_stage_inst_dmem_U9213 ( .A1(MEM_stage_inst_dmem_n13056), .A2(MEM_stage_inst_dmem_n13031), .ZN(MEM_stage_inst_dmem_n13018) );
NAND2_X1 MEM_stage_inst_dmem_U9212 ( .A1(MEM_stage_inst_dmem_ram_342), .A2(MEM_stage_inst_dmem_n13030), .ZN(MEM_stage_inst_dmem_n13019) );
NAND2_X1 MEM_stage_inst_dmem_U9211 ( .A1(MEM_stage_inst_dmem_n13017), .A2(MEM_stage_inst_dmem_n13016), .ZN(MEM_stage_inst_dmem_n12690) );
NAND2_X1 MEM_stage_inst_dmem_U9210 ( .A1(MEM_stage_inst_dmem_n112), .A2(MEM_stage_inst_dmem_n13031), .ZN(MEM_stage_inst_dmem_n13016) );
NAND2_X1 MEM_stage_inst_dmem_U9209 ( .A1(MEM_stage_inst_dmem_ram_343), .A2(MEM_stage_inst_dmem_n13030), .ZN(MEM_stage_inst_dmem_n13017) );
NAND2_X1 MEM_stage_inst_dmem_U9208 ( .A1(MEM_stage_inst_dmem_n13015), .A2(MEM_stage_inst_dmem_n13014), .ZN(MEM_stage_inst_dmem_n12691) );
NAND2_X1 MEM_stage_inst_dmem_U9207 ( .A1(MEM_stage_inst_dmem_n13051), .A2(MEM_stage_inst_dmem_n13031), .ZN(MEM_stage_inst_dmem_n13014) );
NAND2_X1 MEM_stage_inst_dmem_U9206 ( .A1(MEM_stage_inst_dmem_ram_344), .A2(MEM_stage_inst_dmem_n13030), .ZN(MEM_stage_inst_dmem_n13015) );
NAND2_X1 MEM_stage_inst_dmem_U9205 ( .A1(MEM_stage_inst_dmem_n13013), .A2(MEM_stage_inst_dmem_n13012), .ZN(MEM_stage_inst_dmem_n12692) );
NAND2_X1 MEM_stage_inst_dmem_U9204 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n13031), .ZN(MEM_stage_inst_dmem_n13012) );
NAND2_X1 MEM_stage_inst_dmem_U9203 ( .A1(MEM_stage_inst_dmem_ram_345), .A2(MEM_stage_inst_dmem_n13030), .ZN(MEM_stage_inst_dmem_n13013) );
NAND2_X1 MEM_stage_inst_dmem_U9202 ( .A1(MEM_stage_inst_dmem_n13011), .A2(MEM_stage_inst_dmem_n13010), .ZN(MEM_stage_inst_dmem_n12693) );
NAND2_X1 MEM_stage_inst_dmem_U9201 ( .A1(MEM_stage_inst_dmem_n102), .A2(MEM_stage_inst_dmem_n13031), .ZN(MEM_stage_inst_dmem_n13010) );
NAND2_X1 MEM_stage_inst_dmem_U9200 ( .A1(MEM_stage_inst_dmem_ram_346), .A2(MEM_stage_inst_dmem_n13030), .ZN(MEM_stage_inst_dmem_n13011) );
NAND2_X1 MEM_stage_inst_dmem_U9199 ( .A1(MEM_stage_inst_dmem_n13009), .A2(MEM_stage_inst_dmem_n13008), .ZN(MEM_stage_inst_dmem_n12694) );
NAND2_X1 MEM_stage_inst_dmem_U9198 ( .A1(MEM_stage_inst_dmem_n13044), .A2(MEM_stage_inst_dmem_n13031), .ZN(MEM_stage_inst_dmem_n13008) );
NAND2_X1 MEM_stage_inst_dmem_U9197 ( .A1(MEM_stage_inst_dmem_ram_347), .A2(MEM_stage_inst_dmem_n13030), .ZN(MEM_stage_inst_dmem_n13009) );
NAND2_X1 MEM_stage_inst_dmem_U9196 ( .A1(MEM_stage_inst_dmem_n13007), .A2(MEM_stage_inst_dmem_n13006), .ZN(MEM_stage_inst_dmem_n12695) );
NAND2_X1 MEM_stage_inst_dmem_U9195 ( .A1(MEM_stage_inst_dmem_n13041), .A2(MEM_stage_inst_dmem_n13031), .ZN(MEM_stage_inst_dmem_n13006) );
NAND2_X1 MEM_stage_inst_dmem_U9194 ( .A1(MEM_stage_inst_dmem_ram_348), .A2(MEM_stage_inst_dmem_n13030), .ZN(MEM_stage_inst_dmem_n13007) );
NAND2_X1 MEM_stage_inst_dmem_U9193 ( .A1(MEM_stage_inst_dmem_n13005), .A2(MEM_stage_inst_dmem_n13004), .ZN(MEM_stage_inst_dmem_n12696) );
NAND2_X1 MEM_stage_inst_dmem_U9192 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n13031), .ZN(MEM_stage_inst_dmem_n13004) );
NAND2_X1 MEM_stage_inst_dmem_U9191 ( .A1(MEM_stage_inst_dmem_ram_349), .A2(MEM_stage_inst_dmem_n13030), .ZN(MEM_stage_inst_dmem_n13005) );
NAND2_X1 MEM_stage_inst_dmem_U9190 ( .A1(MEM_stage_inst_dmem_n13003), .A2(MEM_stage_inst_dmem_n13002), .ZN(MEM_stage_inst_dmem_n12697) );
NAND2_X1 MEM_stage_inst_dmem_U9189 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n13031), .ZN(MEM_stage_inst_dmem_n13002) );
NAND2_X1 MEM_stage_inst_dmem_U9188 ( .A1(MEM_stage_inst_dmem_ram_350), .A2(MEM_stage_inst_dmem_n13030), .ZN(MEM_stage_inst_dmem_n13003) );
NAND2_X1 MEM_stage_inst_dmem_U9187 ( .A1(MEM_stage_inst_dmem_n13001), .A2(MEM_stage_inst_dmem_n13000), .ZN(MEM_stage_inst_dmem_n12698) );
NAND2_X1 MEM_stage_inst_dmem_U9186 ( .A1(MEM_stage_inst_dmem_n17994), .A2(MEM_stage_inst_dmem_n13031), .ZN(MEM_stage_inst_dmem_n13000) );
INV_X1 MEM_stage_inst_dmem_U9185 ( .A(MEM_stage_inst_dmem_n13030), .ZN(MEM_stage_inst_dmem_n13031) );
NAND2_X1 MEM_stage_inst_dmem_U9184 ( .A1(MEM_stage_inst_dmem_ram_351), .A2(MEM_stage_inst_dmem_n13030), .ZN(MEM_stage_inst_dmem_n13001) );
NAND2_X1 MEM_stage_inst_dmem_U9183 ( .A1(MEM_stage_inst_dmem_n13182), .A2(MEM_stage_inst_dmem_n21284), .ZN(MEM_stage_inst_dmem_n13030) );
NOR2_X2 MEM_stage_inst_dmem_U9182 ( .A1(MEM_stage_inst_dmem_n13034), .A2(MEM_stage_inst_dmem_n13145), .ZN(MEM_stage_inst_dmem_n21284) );
NAND2_X1 MEM_stage_inst_dmem_U9181 ( .A1(MEM_stage_inst_dmem_n12999), .A2(MEM_stage_inst_dmem_n12998), .ZN(MEM_stage_inst_dmem_n12699) );
NAND2_X1 MEM_stage_inst_dmem_U9180 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n12997), .ZN(MEM_stage_inst_dmem_n12998) );
NAND2_X1 MEM_stage_inst_dmem_U9179 ( .A1(MEM_stage_inst_dmem_ram_352), .A2(MEM_stage_inst_dmem_n12996), .ZN(MEM_stage_inst_dmem_n12999) );
NAND2_X1 MEM_stage_inst_dmem_U9178 ( .A1(MEM_stage_inst_dmem_n12995), .A2(MEM_stage_inst_dmem_n12994), .ZN(MEM_stage_inst_dmem_n12700) );
NAND2_X1 MEM_stage_inst_dmem_U9177 ( .A1(MEM_stage_inst_dmem_n109), .A2(MEM_stage_inst_dmem_n12997), .ZN(MEM_stage_inst_dmem_n12994) );
NAND2_X1 MEM_stage_inst_dmem_U9176 ( .A1(MEM_stage_inst_dmem_ram_353), .A2(MEM_stage_inst_dmem_n12996), .ZN(MEM_stage_inst_dmem_n12995) );
NAND2_X1 MEM_stage_inst_dmem_U9175 ( .A1(MEM_stage_inst_dmem_n12993), .A2(MEM_stage_inst_dmem_n12992), .ZN(MEM_stage_inst_dmem_n12701) );
NAND2_X1 MEM_stage_inst_dmem_U9174 ( .A1(MEM_stage_inst_dmem_n18887), .A2(MEM_stage_inst_dmem_n12997), .ZN(MEM_stage_inst_dmem_n12992) );
NAND2_X1 MEM_stage_inst_dmem_U9173 ( .A1(MEM_stage_inst_dmem_ram_354), .A2(MEM_stage_inst_dmem_n12996), .ZN(MEM_stage_inst_dmem_n12993) );
NAND2_X1 MEM_stage_inst_dmem_U9172 ( .A1(MEM_stage_inst_dmem_n12991), .A2(MEM_stage_inst_dmem_n12990), .ZN(MEM_stage_inst_dmem_n12702) );
NAND2_X1 MEM_stage_inst_dmem_U9171 ( .A1(MEM_stage_inst_dmem_n13064), .A2(MEM_stage_inst_dmem_n12997), .ZN(MEM_stage_inst_dmem_n12990) );
NAND2_X1 MEM_stage_inst_dmem_U9170 ( .A1(MEM_stage_inst_dmem_ram_355), .A2(MEM_stage_inst_dmem_n12996), .ZN(MEM_stage_inst_dmem_n12991) );
NAND2_X1 MEM_stage_inst_dmem_U9169 ( .A1(MEM_stage_inst_dmem_n12989), .A2(MEM_stage_inst_dmem_n12988), .ZN(MEM_stage_inst_dmem_n12703) );
NAND2_X1 MEM_stage_inst_dmem_U9168 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n12997), .ZN(MEM_stage_inst_dmem_n12988) );
NAND2_X1 MEM_stage_inst_dmem_U9167 ( .A1(MEM_stage_inst_dmem_ram_356), .A2(MEM_stage_inst_dmem_n12996), .ZN(MEM_stage_inst_dmem_n12989) );
NAND2_X1 MEM_stage_inst_dmem_U9166 ( .A1(MEM_stage_inst_dmem_n12987), .A2(MEM_stage_inst_dmem_n12986), .ZN(MEM_stage_inst_dmem_n12704) );
NAND2_X1 MEM_stage_inst_dmem_U9165 ( .A1(MEM_stage_inst_dmem_n13059), .A2(MEM_stage_inst_dmem_n12997), .ZN(MEM_stage_inst_dmem_n12986) );
NAND2_X1 MEM_stage_inst_dmem_U9164 ( .A1(MEM_stage_inst_dmem_ram_357), .A2(MEM_stage_inst_dmem_n12996), .ZN(MEM_stage_inst_dmem_n12987) );
NAND2_X1 MEM_stage_inst_dmem_U9163 ( .A1(MEM_stage_inst_dmem_n12985), .A2(MEM_stage_inst_dmem_n12984), .ZN(MEM_stage_inst_dmem_n12705) );
NAND2_X1 MEM_stage_inst_dmem_U9162 ( .A1(MEM_stage_inst_dmem_n13056), .A2(MEM_stage_inst_dmem_n12997), .ZN(MEM_stage_inst_dmem_n12984) );
NAND2_X1 MEM_stage_inst_dmem_U9161 ( .A1(MEM_stage_inst_dmem_ram_358), .A2(MEM_stage_inst_dmem_n12996), .ZN(MEM_stage_inst_dmem_n12985) );
NAND2_X1 MEM_stage_inst_dmem_U9160 ( .A1(MEM_stage_inst_dmem_n12983), .A2(MEM_stage_inst_dmem_n12982), .ZN(MEM_stage_inst_dmem_n12706) );
NAND2_X1 MEM_stage_inst_dmem_U9159 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n12997), .ZN(MEM_stage_inst_dmem_n12982) );
NAND2_X1 MEM_stage_inst_dmem_U9158 ( .A1(MEM_stage_inst_dmem_ram_359), .A2(MEM_stage_inst_dmem_n12996), .ZN(MEM_stage_inst_dmem_n12983) );
NAND2_X1 MEM_stage_inst_dmem_U9157 ( .A1(MEM_stage_inst_dmem_n12981), .A2(MEM_stage_inst_dmem_n12980), .ZN(MEM_stage_inst_dmem_n12707) );
NAND2_X1 MEM_stage_inst_dmem_U9156 ( .A1(MEM_stage_inst_dmem_n13051), .A2(MEM_stage_inst_dmem_n12997), .ZN(MEM_stage_inst_dmem_n12980) );
NAND2_X1 MEM_stage_inst_dmem_U9155 ( .A1(MEM_stage_inst_dmem_ram_360), .A2(MEM_stage_inst_dmem_n12996), .ZN(MEM_stage_inst_dmem_n12981) );
NAND2_X1 MEM_stage_inst_dmem_U9154 ( .A1(MEM_stage_inst_dmem_n12979), .A2(MEM_stage_inst_dmem_n12978), .ZN(MEM_stage_inst_dmem_n12708) );
NAND2_X1 MEM_stage_inst_dmem_U9153 ( .A1(MEM_stage_inst_dmem_n19251), .A2(MEM_stage_inst_dmem_n12997), .ZN(MEM_stage_inst_dmem_n12978) );
NAND2_X1 MEM_stage_inst_dmem_U9152 ( .A1(MEM_stage_inst_dmem_ram_361), .A2(MEM_stage_inst_dmem_n12996), .ZN(MEM_stage_inst_dmem_n12979) );
NAND2_X1 MEM_stage_inst_dmem_U9151 ( .A1(MEM_stage_inst_dmem_n12977), .A2(MEM_stage_inst_dmem_n12976), .ZN(MEM_stage_inst_dmem_n12709) );
NAND2_X1 MEM_stage_inst_dmem_U9150 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n12997), .ZN(MEM_stage_inst_dmem_n12976) );
NAND2_X1 MEM_stage_inst_dmem_U9149 ( .A1(MEM_stage_inst_dmem_ram_362), .A2(MEM_stage_inst_dmem_n12996), .ZN(MEM_stage_inst_dmem_n12977) );
NAND2_X1 MEM_stage_inst_dmem_U9148 ( .A1(MEM_stage_inst_dmem_n12975), .A2(MEM_stage_inst_dmem_n12974), .ZN(MEM_stage_inst_dmem_n12710) );
NAND2_X1 MEM_stage_inst_dmem_U9147 ( .A1(MEM_stage_inst_dmem_n13044), .A2(MEM_stage_inst_dmem_n12997), .ZN(MEM_stage_inst_dmem_n12974) );
NAND2_X1 MEM_stage_inst_dmem_U9146 ( .A1(MEM_stage_inst_dmem_ram_363), .A2(MEM_stage_inst_dmem_n12996), .ZN(MEM_stage_inst_dmem_n12975) );
NAND2_X1 MEM_stage_inst_dmem_U9145 ( .A1(MEM_stage_inst_dmem_n12973), .A2(MEM_stage_inst_dmem_n12972), .ZN(MEM_stage_inst_dmem_n12711) );
NAND2_X1 MEM_stage_inst_dmem_U9144 ( .A1(MEM_stage_inst_dmem_n13041), .A2(MEM_stage_inst_dmem_n12997), .ZN(MEM_stage_inst_dmem_n12972) );
NAND2_X1 MEM_stage_inst_dmem_U9143 ( .A1(MEM_stage_inst_dmem_ram_364), .A2(MEM_stage_inst_dmem_n12996), .ZN(MEM_stage_inst_dmem_n12973) );
NAND2_X1 MEM_stage_inst_dmem_U9142 ( .A1(MEM_stage_inst_dmem_n12971), .A2(MEM_stage_inst_dmem_n12970), .ZN(MEM_stage_inst_dmem_n12712) );
NAND2_X1 MEM_stage_inst_dmem_U9141 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n12997), .ZN(MEM_stage_inst_dmem_n12970) );
NAND2_X1 MEM_stage_inst_dmem_U9140 ( .A1(MEM_stage_inst_dmem_ram_365), .A2(MEM_stage_inst_dmem_n12996), .ZN(MEM_stage_inst_dmem_n12971) );
NAND2_X1 MEM_stage_inst_dmem_U9139 ( .A1(MEM_stage_inst_dmem_n12969), .A2(MEM_stage_inst_dmem_n12968), .ZN(MEM_stage_inst_dmem_n12713) );
NAND2_X1 MEM_stage_inst_dmem_U9138 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n12997), .ZN(MEM_stage_inst_dmem_n12968) );
NAND2_X1 MEM_stage_inst_dmem_U9137 ( .A1(MEM_stage_inst_dmem_ram_366), .A2(MEM_stage_inst_dmem_n12996), .ZN(MEM_stage_inst_dmem_n12969) );
NAND2_X1 MEM_stage_inst_dmem_U9136 ( .A1(MEM_stage_inst_dmem_n12967), .A2(MEM_stage_inst_dmem_n12966), .ZN(MEM_stage_inst_dmem_n12714) );
NAND2_X1 MEM_stage_inst_dmem_U9135 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n12997), .ZN(MEM_stage_inst_dmem_n12966) );
NAND2_X1 MEM_stage_inst_dmem_U9134 ( .A1(MEM_stage_inst_dmem_ram_367), .A2(MEM_stage_inst_dmem_n12996), .ZN(MEM_stage_inst_dmem_n12967) );
NAND2_X1 MEM_stage_inst_dmem_U9133 ( .A1(MEM_stage_inst_dmem_n13182), .A2(MEM_stage_inst_dmem_n21249), .ZN(MEM_stage_inst_dmem_n12996) );
NOR2_X2 MEM_stage_inst_dmem_U9132 ( .A1(MEM_stage_inst_dmem_n12965), .A2(MEM_stage_inst_dmem_n13180), .ZN(MEM_stage_inst_dmem_n21249) );
NAND2_X1 MEM_stage_inst_dmem_U9131 ( .A1(MEM_stage_inst_dmem_n12964), .A2(MEM_stage_inst_dmem_n12963), .ZN(MEM_stage_inst_dmem_n13180) );
NAND2_X1 MEM_stage_inst_dmem_U9130 ( .A1(MEM_stage_inst_dmem_n12962), .A2(MEM_stage_inst_dmem_n12961), .ZN(MEM_stage_inst_dmem_n12715) );
NAND2_X1 MEM_stage_inst_dmem_U9129 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n12960), .ZN(MEM_stage_inst_dmem_n12961) );
NAND2_X1 MEM_stage_inst_dmem_U9128 ( .A1(MEM_stage_inst_dmem_ram_368), .A2(MEM_stage_inst_dmem_n12959), .ZN(MEM_stage_inst_dmem_n12962) );
NAND2_X1 MEM_stage_inst_dmem_U9127 ( .A1(MEM_stage_inst_dmem_n12958), .A2(MEM_stage_inst_dmem_n12957), .ZN(MEM_stage_inst_dmem_n12716) );
NAND2_X1 MEM_stage_inst_dmem_U9126 ( .A1(MEM_stage_inst_dmem_n109), .A2(MEM_stage_inst_dmem_n12960), .ZN(MEM_stage_inst_dmem_n12957) );
NAND2_X1 MEM_stage_inst_dmem_U9125 ( .A1(MEM_stage_inst_dmem_ram_369), .A2(MEM_stage_inst_dmem_n12959), .ZN(MEM_stage_inst_dmem_n12958) );
NAND2_X1 MEM_stage_inst_dmem_U9124 ( .A1(MEM_stage_inst_dmem_n12956), .A2(MEM_stage_inst_dmem_n12955), .ZN(MEM_stage_inst_dmem_n12717) );
NAND2_X1 MEM_stage_inst_dmem_U9123 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n12960), .ZN(MEM_stage_inst_dmem_n12955) );
NAND2_X1 MEM_stage_inst_dmem_U9122 ( .A1(MEM_stage_inst_dmem_ram_370), .A2(MEM_stage_inst_dmem_n12959), .ZN(MEM_stage_inst_dmem_n12956) );
NAND2_X1 MEM_stage_inst_dmem_U9121 ( .A1(MEM_stage_inst_dmem_n12954), .A2(MEM_stage_inst_dmem_n12953), .ZN(MEM_stage_inst_dmem_n12718) );
NAND2_X1 MEM_stage_inst_dmem_U9120 ( .A1(MEM_stage_inst_dmem_n13064), .A2(MEM_stage_inst_dmem_n12960), .ZN(MEM_stage_inst_dmem_n12953) );
NAND2_X1 MEM_stage_inst_dmem_U9119 ( .A1(MEM_stage_inst_dmem_ram_371), .A2(MEM_stage_inst_dmem_n12959), .ZN(MEM_stage_inst_dmem_n12954) );
NAND2_X1 MEM_stage_inst_dmem_U9118 ( .A1(MEM_stage_inst_dmem_n12952), .A2(MEM_stage_inst_dmem_n12951), .ZN(MEM_stage_inst_dmem_n12719) );
NAND2_X1 MEM_stage_inst_dmem_U9117 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n12960), .ZN(MEM_stage_inst_dmem_n12951) );
NAND2_X1 MEM_stage_inst_dmem_U9116 ( .A1(MEM_stage_inst_dmem_ram_372), .A2(MEM_stage_inst_dmem_n12959), .ZN(MEM_stage_inst_dmem_n12952) );
NAND2_X1 MEM_stage_inst_dmem_U9115 ( .A1(MEM_stage_inst_dmem_n12950), .A2(MEM_stage_inst_dmem_n12949), .ZN(MEM_stage_inst_dmem_n12720) );
NAND2_X1 MEM_stage_inst_dmem_U9114 ( .A1(MEM_stage_inst_dmem_n13059), .A2(MEM_stage_inst_dmem_n12960), .ZN(MEM_stage_inst_dmem_n12949) );
NAND2_X1 MEM_stage_inst_dmem_U9113 ( .A1(MEM_stage_inst_dmem_ram_373), .A2(MEM_stage_inst_dmem_n12959), .ZN(MEM_stage_inst_dmem_n12950) );
NAND2_X1 MEM_stage_inst_dmem_U9112 ( .A1(MEM_stage_inst_dmem_n12948), .A2(MEM_stage_inst_dmem_n12947), .ZN(MEM_stage_inst_dmem_n12721) );
NAND2_X1 MEM_stage_inst_dmem_U9111 ( .A1(MEM_stage_inst_dmem_n13056), .A2(MEM_stage_inst_dmem_n12960), .ZN(MEM_stage_inst_dmem_n12947) );
NAND2_X1 MEM_stage_inst_dmem_U9110 ( .A1(MEM_stage_inst_dmem_ram_374), .A2(MEM_stage_inst_dmem_n12959), .ZN(MEM_stage_inst_dmem_n12948) );
NAND2_X1 MEM_stage_inst_dmem_U9109 ( .A1(MEM_stage_inst_dmem_n12946), .A2(MEM_stage_inst_dmem_n12945), .ZN(MEM_stage_inst_dmem_n12722) );
NAND2_X1 MEM_stage_inst_dmem_U9108 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n12960), .ZN(MEM_stage_inst_dmem_n12945) );
NAND2_X1 MEM_stage_inst_dmem_U9107 ( .A1(MEM_stage_inst_dmem_ram_375), .A2(MEM_stage_inst_dmem_n12959), .ZN(MEM_stage_inst_dmem_n12946) );
NAND2_X1 MEM_stage_inst_dmem_U9106 ( .A1(MEM_stage_inst_dmem_n12944), .A2(MEM_stage_inst_dmem_n12943), .ZN(MEM_stage_inst_dmem_n12723) );
NAND2_X1 MEM_stage_inst_dmem_U9105 ( .A1(MEM_stage_inst_dmem_n13051), .A2(MEM_stage_inst_dmem_n12960), .ZN(MEM_stage_inst_dmem_n12943) );
NAND2_X1 MEM_stage_inst_dmem_U9104 ( .A1(MEM_stage_inst_dmem_ram_376), .A2(MEM_stage_inst_dmem_n12959), .ZN(MEM_stage_inst_dmem_n12944) );
NAND2_X1 MEM_stage_inst_dmem_U9103 ( .A1(MEM_stage_inst_dmem_n12942), .A2(MEM_stage_inst_dmem_n12941), .ZN(MEM_stage_inst_dmem_n12724) );
NAND2_X1 MEM_stage_inst_dmem_U9102 ( .A1(MEM_stage_inst_dmem_n13880), .A2(MEM_stage_inst_dmem_n12960), .ZN(MEM_stage_inst_dmem_n12941) );
NAND2_X1 MEM_stage_inst_dmem_U9101 ( .A1(MEM_stage_inst_dmem_ram_377), .A2(MEM_stage_inst_dmem_n12959), .ZN(MEM_stage_inst_dmem_n12942) );
NAND2_X1 MEM_stage_inst_dmem_U9100 ( .A1(MEM_stage_inst_dmem_n12940), .A2(MEM_stage_inst_dmem_n12939), .ZN(MEM_stage_inst_dmem_n12725) );
NAND2_X1 MEM_stage_inst_dmem_U9099 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n12960), .ZN(MEM_stage_inst_dmem_n12939) );
NAND2_X1 MEM_stage_inst_dmem_U9098 ( .A1(MEM_stage_inst_dmem_ram_378), .A2(MEM_stage_inst_dmem_n12959), .ZN(MEM_stage_inst_dmem_n12940) );
NAND2_X1 MEM_stage_inst_dmem_U9097 ( .A1(MEM_stage_inst_dmem_n12938), .A2(MEM_stage_inst_dmem_n12937), .ZN(MEM_stage_inst_dmem_n12726) );
NAND2_X1 MEM_stage_inst_dmem_U9096 ( .A1(MEM_stage_inst_dmem_n13044), .A2(MEM_stage_inst_dmem_n12960), .ZN(MEM_stage_inst_dmem_n12937) );
NAND2_X1 MEM_stage_inst_dmem_U9095 ( .A1(MEM_stage_inst_dmem_ram_379), .A2(MEM_stage_inst_dmem_n12959), .ZN(MEM_stage_inst_dmem_n12938) );
NAND2_X1 MEM_stage_inst_dmem_U9094 ( .A1(MEM_stage_inst_dmem_n12936), .A2(MEM_stage_inst_dmem_n12935), .ZN(MEM_stage_inst_dmem_n12727) );
NAND2_X1 MEM_stage_inst_dmem_U9093 ( .A1(MEM_stage_inst_dmem_n13041), .A2(MEM_stage_inst_dmem_n12960), .ZN(MEM_stage_inst_dmem_n12935) );
NAND2_X1 MEM_stage_inst_dmem_U9092 ( .A1(MEM_stage_inst_dmem_ram_380), .A2(MEM_stage_inst_dmem_n12959), .ZN(MEM_stage_inst_dmem_n12936) );
NAND2_X1 MEM_stage_inst_dmem_U9091 ( .A1(MEM_stage_inst_dmem_n12934), .A2(MEM_stage_inst_dmem_n12933), .ZN(MEM_stage_inst_dmem_n12728) );
NAND2_X1 MEM_stage_inst_dmem_U9090 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n12960), .ZN(MEM_stage_inst_dmem_n12933) );
NAND2_X1 MEM_stage_inst_dmem_U9089 ( .A1(MEM_stage_inst_dmem_ram_381), .A2(MEM_stage_inst_dmem_n12959), .ZN(MEM_stage_inst_dmem_n12934) );
NAND2_X1 MEM_stage_inst_dmem_U9088 ( .A1(MEM_stage_inst_dmem_n12932), .A2(MEM_stage_inst_dmem_n12931), .ZN(MEM_stage_inst_dmem_n12729) );
NAND2_X1 MEM_stage_inst_dmem_U9087 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n12960), .ZN(MEM_stage_inst_dmem_n12931) );
NAND2_X1 MEM_stage_inst_dmem_U9086 ( .A1(MEM_stage_inst_dmem_ram_382), .A2(MEM_stage_inst_dmem_n12959), .ZN(MEM_stage_inst_dmem_n12932) );
NAND2_X1 MEM_stage_inst_dmem_U9085 ( .A1(MEM_stage_inst_dmem_n12930), .A2(MEM_stage_inst_dmem_n12929), .ZN(MEM_stage_inst_dmem_n12730) );
NAND2_X1 MEM_stage_inst_dmem_U9084 ( .A1(MEM_stage_inst_dmem_n16343), .A2(MEM_stage_inst_dmem_n12960), .ZN(MEM_stage_inst_dmem_n12929) );
INV_X1 MEM_stage_inst_dmem_U9083 ( .A(MEM_stage_inst_dmem_n12959), .ZN(MEM_stage_inst_dmem_n12960) );
NAND2_X1 MEM_stage_inst_dmem_U9082 ( .A1(MEM_stage_inst_dmem_ram_383), .A2(MEM_stage_inst_dmem_n12959), .ZN(MEM_stage_inst_dmem_n12930) );
NAND2_X1 MEM_stage_inst_dmem_U9081 ( .A1(MEM_stage_inst_dmem_n13182), .A2(MEM_stage_inst_dmem_n21214), .ZN(MEM_stage_inst_dmem_n12959) );
NOR2_X2 MEM_stage_inst_dmem_U9080 ( .A1(MEM_stage_inst_dmem_n12965), .A2(MEM_stage_inst_dmem_n13145), .ZN(MEM_stage_inst_dmem_n21214) );
NAND2_X1 MEM_stage_inst_dmem_U9079 ( .A1(EX_pipeline_reg_out_22), .A2(MEM_stage_inst_dmem_n12964), .ZN(MEM_stage_inst_dmem_n13145) );
NAND2_X1 MEM_stage_inst_dmem_U9078 ( .A1(MEM_stage_inst_dmem_n12928), .A2(MEM_stage_inst_dmem_n12927), .ZN(MEM_stage_inst_dmem_n12731) );
NAND2_X1 MEM_stage_inst_dmem_U9077 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n12926), .ZN(MEM_stage_inst_dmem_n12927) );
NAND2_X1 MEM_stage_inst_dmem_U9076 ( .A1(MEM_stage_inst_dmem_ram_384), .A2(MEM_stage_inst_dmem_n12925), .ZN(MEM_stage_inst_dmem_n12928) );
NAND2_X1 MEM_stage_inst_dmem_U9075 ( .A1(MEM_stage_inst_dmem_n12924), .A2(MEM_stage_inst_dmem_n12923), .ZN(MEM_stage_inst_dmem_n12732) );
NAND2_X1 MEM_stage_inst_dmem_U9074 ( .A1(MEM_stage_inst_dmem_n109), .A2(MEM_stage_inst_dmem_n12926), .ZN(MEM_stage_inst_dmem_n12923) );
NAND2_X1 MEM_stage_inst_dmem_U9073 ( .A1(MEM_stage_inst_dmem_ram_385), .A2(MEM_stage_inst_dmem_n12925), .ZN(MEM_stage_inst_dmem_n12924) );
NAND2_X1 MEM_stage_inst_dmem_U9072 ( .A1(MEM_stage_inst_dmem_n12922), .A2(MEM_stage_inst_dmem_n12921), .ZN(MEM_stage_inst_dmem_n12733) );
NAND2_X1 MEM_stage_inst_dmem_U9071 ( .A1(MEM_stage_inst_dmem_n16789), .A2(MEM_stage_inst_dmem_n12926), .ZN(MEM_stage_inst_dmem_n12921) );
NAND2_X1 MEM_stage_inst_dmem_U9070 ( .A1(MEM_stage_inst_dmem_ram_386), .A2(MEM_stage_inst_dmem_n12925), .ZN(MEM_stage_inst_dmem_n12922) );
NAND2_X1 MEM_stage_inst_dmem_U9069 ( .A1(MEM_stage_inst_dmem_n12920), .A2(MEM_stage_inst_dmem_n12919), .ZN(MEM_stage_inst_dmem_n12734) );
NAND2_X1 MEM_stage_inst_dmem_U9068 ( .A1(MEM_stage_inst_dmem_n13064), .A2(MEM_stage_inst_dmem_n12926), .ZN(MEM_stage_inst_dmem_n12919) );
NAND2_X1 MEM_stage_inst_dmem_U9067 ( .A1(MEM_stage_inst_dmem_ram_387), .A2(MEM_stage_inst_dmem_n12925), .ZN(MEM_stage_inst_dmem_n12920) );
NAND2_X1 MEM_stage_inst_dmem_U9066 ( .A1(MEM_stage_inst_dmem_n12918), .A2(MEM_stage_inst_dmem_n12917), .ZN(MEM_stage_inst_dmem_n12735) );
NAND2_X1 MEM_stage_inst_dmem_U9065 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n12926), .ZN(MEM_stage_inst_dmem_n12917) );
NAND2_X1 MEM_stage_inst_dmem_U9064 ( .A1(MEM_stage_inst_dmem_ram_388), .A2(MEM_stage_inst_dmem_n12925), .ZN(MEM_stage_inst_dmem_n12918) );
NAND2_X1 MEM_stage_inst_dmem_U9063 ( .A1(MEM_stage_inst_dmem_n12916), .A2(MEM_stage_inst_dmem_n12915), .ZN(MEM_stage_inst_dmem_n12736) );
NAND2_X1 MEM_stage_inst_dmem_U9062 ( .A1(MEM_stage_inst_dmem_n13059), .A2(MEM_stage_inst_dmem_n12926), .ZN(MEM_stage_inst_dmem_n12915) );
NAND2_X1 MEM_stage_inst_dmem_U9061 ( .A1(MEM_stage_inst_dmem_ram_389), .A2(MEM_stage_inst_dmem_n12925), .ZN(MEM_stage_inst_dmem_n12916) );
NAND2_X1 MEM_stage_inst_dmem_U9060 ( .A1(MEM_stage_inst_dmem_n12914), .A2(MEM_stage_inst_dmem_n12913), .ZN(MEM_stage_inst_dmem_n12737) );
NAND2_X1 MEM_stage_inst_dmem_U9059 ( .A1(MEM_stage_inst_dmem_n13056), .A2(MEM_stage_inst_dmem_n12926), .ZN(MEM_stage_inst_dmem_n12913) );
NAND2_X1 MEM_stage_inst_dmem_U9058 ( .A1(MEM_stage_inst_dmem_ram_390), .A2(MEM_stage_inst_dmem_n12925), .ZN(MEM_stage_inst_dmem_n12914) );
NAND2_X1 MEM_stage_inst_dmem_U9057 ( .A1(MEM_stage_inst_dmem_n12912), .A2(MEM_stage_inst_dmem_n12911), .ZN(MEM_stage_inst_dmem_n12738) );
NAND2_X1 MEM_stage_inst_dmem_U9056 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n12926), .ZN(MEM_stage_inst_dmem_n12911) );
NAND2_X1 MEM_stage_inst_dmem_U9055 ( .A1(MEM_stage_inst_dmem_ram_391), .A2(MEM_stage_inst_dmem_n12925), .ZN(MEM_stage_inst_dmem_n12912) );
NAND2_X1 MEM_stage_inst_dmem_U9054 ( .A1(MEM_stage_inst_dmem_n12910), .A2(MEM_stage_inst_dmem_n12909), .ZN(MEM_stage_inst_dmem_n12739) );
NAND2_X1 MEM_stage_inst_dmem_U9053 ( .A1(MEM_stage_inst_dmem_n13051), .A2(MEM_stage_inst_dmem_n12926), .ZN(MEM_stage_inst_dmem_n12909) );
NAND2_X1 MEM_stage_inst_dmem_U9052 ( .A1(MEM_stage_inst_dmem_ram_392), .A2(MEM_stage_inst_dmem_n12925), .ZN(MEM_stage_inst_dmem_n12910) );
NAND2_X1 MEM_stage_inst_dmem_U9051 ( .A1(MEM_stage_inst_dmem_n12908), .A2(MEM_stage_inst_dmem_n12907), .ZN(MEM_stage_inst_dmem_n12740) );
NAND2_X1 MEM_stage_inst_dmem_U9050 ( .A1(MEM_stage_inst_dmem_n100), .A2(MEM_stage_inst_dmem_n12926), .ZN(MEM_stage_inst_dmem_n12907) );
NAND2_X1 MEM_stage_inst_dmem_U9049 ( .A1(MEM_stage_inst_dmem_ram_393), .A2(MEM_stage_inst_dmem_n12925), .ZN(MEM_stage_inst_dmem_n12908) );
NAND2_X1 MEM_stage_inst_dmem_U9048 ( .A1(MEM_stage_inst_dmem_n12906), .A2(MEM_stage_inst_dmem_n12905), .ZN(MEM_stage_inst_dmem_n12741) );
NAND2_X1 MEM_stage_inst_dmem_U9047 ( .A1(MEM_stage_inst_dmem_n18007), .A2(MEM_stage_inst_dmem_n12926), .ZN(MEM_stage_inst_dmem_n12905) );
NAND2_X1 MEM_stage_inst_dmem_U9046 ( .A1(MEM_stage_inst_dmem_ram_394), .A2(MEM_stage_inst_dmem_n12925), .ZN(MEM_stage_inst_dmem_n12906) );
NAND2_X1 MEM_stage_inst_dmem_U9045 ( .A1(MEM_stage_inst_dmem_n12904), .A2(MEM_stage_inst_dmem_n12903), .ZN(MEM_stage_inst_dmem_n12742) );
NAND2_X1 MEM_stage_inst_dmem_U9044 ( .A1(MEM_stage_inst_dmem_n13044), .A2(MEM_stage_inst_dmem_n12926), .ZN(MEM_stage_inst_dmem_n12903) );
NAND2_X1 MEM_stage_inst_dmem_U9043 ( .A1(MEM_stage_inst_dmem_ram_395), .A2(MEM_stage_inst_dmem_n12925), .ZN(MEM_stage_inst_dmem_n12904) );
NAND2_X1 MEM_stage_inst_dmem_U9042 ( .A1(MEM_stage_inst_dmem_n12902), .A2(MEM_stage_inst_dmem_n12901), .ZN(MEM_stage_inst_dmem_n12743) );
NAND2_X1 MEM_stage_inst_dmem_U9041 ( .A1(MEM_stage_inst_dmem_n13041), .A2(MEM_stage_inst_dmem_n12926), .ZN(MEM_stage_inst_dmem_n12901) );
NAND2_X1 MEM_stage_inst_dmem_U9040 ( .A1(MEM_stage_inst_dmem_ram_396), .A2(MEM_stage_inst_dmem_n12925), .ZN(MEM_stage_inst_dmem_n12902) );
NAND2_X1 MEM_stage_inst_dmem_U9039 ( .A1(MEM_stage_inst_dmem_n12900), .A2(MEM_stage_inst_dmem_n12899), .ZN(MEM_stage_inst_dmem_n12744) );
NAND2_X1 MEM_stage_inst_dmem_U9038 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n12926), .ZN(MEM_stage_inst_dmem_n12899) );
NAND2_X1 MEM_stage_inst_dmem_U9037 ( .A1(MEM_stage_inst_dmem_ram_397), .A2(MEM_stage_inst_dmem_n12925), .ZN(MEM_stage_inst_dmem_n12900) );
NAND2_X1 MEM_stage_inst_dmem_U9036 ( .A1(MEM_stage_inst_dmem_n12898), .A2(MEM_stage_inst_dmem_n12897), .ZN(MEM_stage_inst_dmem_n12745) );
NAND2_X1 MEM_stage_inst_dmem_U9035 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n12926), .ZN(MEM_stage_inst_dmem_n12897) );
NAND2_X1 MEM_stage_inst_dmem_U9034 ( .A1(MEM_stage_inst_dmem_ram_398), .A2(MEM_stage_inst_dmem_n12925), .ZN(MEM_stage_inst_dmem_n12898) );
NAND2_X1 MEM_stage_inst_dmem_U9033 ( .A1(MEM_stage_inst_dmem_n12896), .A2(MEM_stage_inst_dmem_n12895), .ZN(MEM_stage_inst_dmem_n12746) );
NAND2_X1 MEM_stage_inst_dmem_U9032 ( .A1(MEM_stage_inst_dmem_n14693), .A2(MEM_stage_inst_dmem_n12926), .ZN(MEM_stage_inst_dmem_n12895) );
INV_X1 MEM_stage_inst_dmem_U9031 ( .A(MEM_stage_inst_dmem_n12925), .ZN(MEM_stage_inst_dmem_n12926) );
NAND2_X1 MEM_stage_inst_dmem_U9030 ( .A1(MEM_stage_inst_dmem_ram_399), .A2(MEM_stage_inst_dmem_n12925), .ZN(MEM_stage_inst_dmem_n12896) );
NAND2_X1 MEM_stage_inst_dmem_U9029 ( .A1(MEM_stage_inst_dmem_n13182), .A2(MEM_stage_inst_dmem_n21179), .ZN(MEM_stage_inst_dmem_n12925) );
NOR2_X2 MEM_stage_inst_dmem_U9028 ( .A1(MEM_stage_inst_dmem_n12894), .A2(MEM_stage_inst_dmem_n13181), .ZN(MEM_stage_inst_dmem_n21179) );
NAND2_X1 MEM_stage_inst_dmem_U9027 ( .A1(MEM_stage_inst_dmem_n12893), .A2(MEM_stage_inst_dmem_n12892), .ZN(MEM_stage_inst_dmem_n12747) );
NAND2_X1 MEM_stage_inst_dmem_U9026 ( .A1(MEM_stage_inst_dmem_n15145), .A2(MEM_stage_inst_dmem_n12891), .ZN(MEM_stage_inst_dmem_n12892) );
NAND2_X1 MEM_stage_inst_dmem_U9025 ( .A1(MEM_stage_inst_dmem_ram_400), .A2(MEM_stage_inst_dmem_n12890), .ZN(MEM_stage_inst_dmem_n12893) );
NAND2_X1 MEM_stage_inst_dmem_U9024 ( .A1(MEM_stage_inst_dmem_n12889), .A2(MEM_stage_inst_dmem_n12888), .ZN(MEM_stage_inst_dmem_n12748) );
NAND2_X1 MEM_stage_inst_dmem_U9023 ( .A1(MEM_stage_inst_dmem_n109), .A2(MEM_stage_inst_dmem_n12891), .ZN(MEM_stage_inst_dmem_n12888) );
NAND2_X1 MEM_stage_inst_dmem_U9022 ( .A1(MEM_stage_inst_dmem_ram_401), .A2(MEM_stage_inst_dmem_n12890), .ZN(MEM_stage_inst_dmem_n12889) );
NAND2_X1 MEM_stage_inst_dmem_U9021 ( .A1(MEM_stage_inst_dmem_n12887), .A2(MEM_stage_inst_dmem_n12886), .ZN(MEM_stage_inst_dmem_n12749) );
NAND2_X1 MEM_stage_inst_dmem_U9020 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n12891), .ZN(MEM_stage_inst_dmem_n12886) );
NAND2_X1 MEM_stage_inst_dmem_U9019 ( .A1(MEM_stage_inst_dmem_ram_402), .A2(MEM_stage_inst_dmem_n12890), .ZN(MEM_stage_inst_dmem_n12887) );
NAND2_X1 MEM_stage_inst_dmem_U9018 ( .A1(MEM_stage_inst_dmem_n12885), .A2(MEM_stage_inst_dmem_n12884), .ZN(MEM_stage_inst_dmem_n12750) );
NAND2_X1 MEM_stage_inst_dmem_U9017 ( .A1(MEM_stage_inst_dmem_n13064), .A2(MEM_stage_inst_dmem_n12891), .ZN(MEM_stage_inst_dmem_n12884) );
NAND2_X1 MEM_stage_inst_dmem_U9016 ( .A1(MEM_stage_inst_dmem_ram_403), .A2(MEM_stage_inst_dmem_n12890), .ZN(MEM_stage_inst_dmem_n12885) );
NAND2_X1 MEM_stage_inst_dmem_U9015 ( .A1(MEM_stage_inst_dmem_n12883), .A2(MEM_stage_inst_dmem_n12882), .ZN(MEM_stage_inst_dmem_n12751) );
NAND2_X1 MEM_stage_inst_dmem_U9014 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n12891), .ZN(MEM_stage_inst_dmem_n12882) );
NAND2_X1 MEM_stage_inst_dmem_U9013 ( .A1(MEM_stage_inst_dmem_ram_404), .A2(MEM_stage_inst_dmem_n12890), .ZN(MEM_stage_inst_dmem_n12883) );
NAND2_X1 MEM_stage_inst_dmem_U9012 ( .A1(MEM_stage_inst_dmem_n12881), .A2(MEM_stage_inst_dmem_n12880), .ZN(MEM_stage_inst_dmem_n12752) );
NAND2_X1 MEM_stage_inst_dmem_U9011 ( .A1(MEM_stage_inst_dmem_n13059), .A2(MEM_stage_inst_dmem_n12891), .ZN(MEM_stage_inst_dmem_n12880) );
NAND2_X1 MEM_stage_inst_dmem_U9010 ( .A1(MEM_stage_inst_dmem_ram_405), .A2(MEM_stage_inst_dmem_n12890), .ZN(MEM_stage_inst_dmem_n12881) );
NAND2_X1 MEM_stage_inst_dmem_U9009 ( .A1(MEM_stage_inst_dmem_n12879), .A2(MEM_stage_inst_dmem_n12878), .ZN(MEM_stage_inst_dmem_n12753) );
NAND2_X1 MEM_stage_inst_dmem_U9008 ( .A1(MEM_stage_inst_dmem_n13056), .A2(MEM_stage_inst_dmem_n12891), .ZN(MEM_stage_inst_dmem_n12878) );
NAND2_X1 MEM_stage_inst_dmem_U9007 ( .A1(MEM_stage_inst_dmem_ram_406), .A2(MEM_stage_inst_dmem_n12890), .ZN(MEM_stage_inst_dmem_n12879) );
NAND2_X1 MEM_stage_inst_dmem_U9006 ( .A1(MEM_stage_inst_dmem_n12877), .A2(MEM_stage_inst_dmem_n12876), .ZN(MEM_stage_inst_dmem_n12754) );
NAND2_X1 MEM_stage_inst_dmem_U9005 ( .A1(MEM_stage_inst_dmem_n16361), .A2(MEM_stage_inst_dmem_n12891), .ZN(MEM_stage_inst_dmem_n12876) );
NAND2_X1 MEM_stage_inst_dmem_U9004 ( .A1(MEM_stage_inst_dmem_ram_407), .A2(MEM_stage_inst_dmem_n12890), .ZN(MEM_stage_inst_dmem_n12877) );
NAND2_X1 MEM_stage_inst_dmem_U9003 ( .A1(MEM_stage_inst_dmem_n12875), .A2(MEM_stage_inst_dmem_n12874), .ZN(MEM_stage_inst_dmem_n12755) );
NAND2_X1 MEM_stage_inst_dmem_U9002 ( .A1(MEM_stage_inst_dmem_n13051), .A2(MEM_stage_inst_dmem_n12891), .ZN(MEM_stage_inst_dmem_n12874) );
NAND2_X1 MEM_stage_inst_dmem_U9001 ( .A1(MEM_stage_inst_dmem_ram_408), .A2(MEM_stage_inst_dmem_n12890), .ZN(MEM_stage_inst_dmem_n12875) );
NAND2_X1 MEM_stage_inst_dmem_U9000 ( .A1(MEM_stage_inst_dmem_n12873), .A2(MEM_stage_inst_dmem_n12872), .ZN(MEM_stage_inst_dmem_n12756) );
NAND2_X1 MEM_stage_inst_dmem_U8999 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n12891), .ZN(MEM_stage_inst_dmem_n12872) );
NAND2_X1 MEM_stage_inst_dmem_U8998 ( .A1(MEM_stage_inst_dmem_ram_409), .A2(MEM_stage_inst_dmem_n12890), .ZN(MEM_stage_inst_dmem_n12873) );
NAND2_X1 MEM_stage_inst_dmem_U8997 ( .A1(MEM_stage_inst_dmem_n12871), .A2(MEM_stage_inst_dmem_n12870), .ZN(MEM_stage_inst_dmem_n12757) );
NAND2_X1 MEM_stage_inst_dmem_U8996 ( .A1(MEM_stage_inst_dmem_n13877), .A2(MEM_stage_inst_dmem_n12891), .ZN(MEM_stage_inst_dmem_n12870) );
NAND2_X1 MEM_stage_inst_dmem_U8995 ( .A1(MEM_stage_inst_dmem_ram_410), .A2(MEM_stage_inst_dmem_n12890), .ZN(MEM_stage_inst_dmem_n12871) );
NAND2_X1 MEM_stage_inst_dmem_U8994 ( .A1(MEM_stage_inst_dmem_n12869), .A2(MEM_stage_inst_dmem_n12868), .ZN(MEM_stage_inst_dmem_n12758) );
NAND2_X1 MEM_stage_inst_dmem_U8993 ( .A1(MEM_stage_inst_dmem_n13044), .A2(MEM_stage_inst_dmem_n12891), .ZN(MEM_stage_inst_dmem_n12868) );
NAND2_X1 MEM_stage_inst_dmem_U8992 ( .A1(MEM_stage_inst_dmem_ram_411), .A2(MEM_stage_inst_dmem_n12890), .ZN(MEM_stage_inst_dmem_n12869) );
NAND2_X1 MEM_stage_inst_dmem_U8991 ( .A1(MEM_stage_inst_dmem_n12867), .A2(MEM_stage_inst_dmem_n12866), .ZN(MEM_stage_inst_dmem_n12759) );
NAND2_X1 MEM_stage_inst_dmem_U8990 ( .A1(MEM_stage_inst_dmem_n13041), .A2(MEM_stage_inst_dmem_n12891), .ZN(MEM_stage_inst_dmem_n12866) );
NAND2_X1 MEM_stage_inst_dmem_U8989 ( .A1(MEM_stage_inst_dmem_ram_412), .A2(MEM_stage_inst_dmem_n12890), .ZN(MEM_stage_inst_dmem_n12867) );
NAND2_X1 MEM_stage_inst_dmem_U8988 ( .A1(MEM_stage_inst_dmem_n12865), .A2(MEM_stage_inst_dmem_n12864), .ZN(MEM_stage_inst_dmem_n12760) );
NAND2_X1 MEM_stage_inst_dmem_U8987 ( .A1(MEM_stage_inst_dmem_n15116), .A2(MEM_stage_inst_dmem_n12891), .ZN(MEM_stage_inst_dmem_n12864) );
NAND2_X1 MEM_stage_inst_dmem_U8986 ( .A1(MEM_stage_inst_dmem_ram_413), .A2(MEM_stage_inst_dmem_n12890), .ZN(MEM_stage_inst_dmem_n12865) );
NAND2_X1 MEM_stage_inst_dmem_U8985 ( .A1(MEM_stage_inst_dmem_n12863), .A2(MEM_stage_inst_dmem_n12862), .ZN(MEM_stage_inst_dmem_n12761) );
NAND2_X1 MEM_stage_inst_dmem_U8984 ( .A1(MEM_stage_inst_dmem_n15113), .A2(MEM_stage_inst_dmem_n12891), .ZN(MEM_stage_inst_dmem_n12862) );
NAND2_X1 MEM_stage_inst_dmem_U8983 ( .A1(MEM_stage_inst_dmem_ram_414), .A2(MEM_stage_inst_dmem_n12890), .ZN(MEM_stage_inst_dmem_n12863) );
NAND2_X1 MEM_stage_inst_dmem_U8982 ( .A1(MEM_stage_inst_dmem_n12861), .A2(MEM_stage_inst_dmem_n12860), .ZN(MEM_stage_inst_dmem_n12762) );
NAND2_X1 MEM_stage_inst_dmem_U8981 ( .A1(MEM_stage_inst_dmem_n15110), .A2(MEM_stage_inst_dmem_n12891), .ZN(MEM_stage_inst_dmem_n12860) );
INV_X1 MEM_stage_inst_dmem_U8980 ( .A(MEM_stage_inst_dmem_n12890), .ZN(MEM_stage_inst_dmem_n12891) );
NAND2_X1 MEM_stage_inst_dmem_U8979 ( .A1(MEM_stage_inst_dmem_ram_415), .A2(MEM_stage_inst_dmem_n12890), .ZN(MEM_stage_inst_dmem_n12861) );
NAND2_X1 MEM_stage_inst_dmem_U8978 ( .A1(MEM_stage_inst_dmem_n13182), .A2(MEM_stage_inst_dmem_n21144), .ZN(MEM_stage_inst_dmem_n12890) );
NOR2_X2 MEM_stage_inst_dmem_U8977 ( .A1(MEM_stage_inst_dmem_n12859), .A2(MEM_stage_inst_dmem_n13181), .ZN(MEM_stage_inst_dmem_n21144) );
NAND2_X1 MEM_stage_inst_dmem_U8976 ( .A1(MEM_stage_inst_dmem_n8762), .A2(MEM_stage_inst_dmem_n8761), .ZN(MEM_stage_inst_dmem_n13181) );
NAND2_X1 MEM_stage_inst_dmem_U8975 ( .A1(MEM_stage_inst_dmem_n8760), .A2(MEM_stage_inst_dmem_n8759), .ZN(MEM_stage_inst_dmem_n12763) );
NAND2_X1 MEM_stage_inst_dmem_U8974 ( .A1(EX_pipeline_reg_out_5), .A2(MEM_stage_inst_dmem_n8758), .ZN(MEM_stage_inst_dmem_n8759) );
NAND2_X1 MEM_stage_inst_dmem_U8973 ( .A1(MEM_stage_inst_dmem_ram_416), .A2(MEM_stage_inst_dmem_n8757), .ZN(MEM_stage_inst_dmem_n8760) );
NAND2_X1 MEM_stage_inst_dmem_U8972 ( .A1(MEM_stage_inst_dmem_n8756), .A2(MEM_stage_inst_dmem_n8755), .ZN(MEM_stage_inst_dmem_n12764) );
NAND2_X1 MEM_stage_inst_dmem_U8971 ( .A1(MEM_stage_inst_dmem_n109), .A2(MEM_stage_inst_dmem_n8758), .ZN(MEM_stage_inst_dmem_n8755) );
NAND2_X1 MEM_stage_inst_dmem_U8970 ( .A1(MEM_stage_inst_dmem_ram_417), .A2(MEM_stage_inst_dmem_n8757), .ZN(MEM_stage_inst_dmem_n8756) );
NAND2_X1 MEM_stage_inst_dmem_U8969 ( .A1(MEM_stage_inst_dmem_n8754), .A2(MEM_stage_inst_dmem_n8753), .ZN(MEM_stage_inst_dmem_n12765) );
NAND2_X1 MEM_stage_inst_dmem_U8968 ( .A1(MEM_stage_inst_dmem_n18027), .A2(MEM_stage_inst_dmem_n8758), .ZN(MEM_stage_inst_dmem_n8753) );
NAND2_X1 MEM_stage_inst_dmem_U8967 ( .A1(MEM_stage_inst_dmem_ram_418), .A2(MEM_stage_inst_dmem_n8757), .ZN(MEM_stage_inst_dmem_n8754) );
NAND2_X1 MEM_stage_inst_dmem_U8966 ( .A1(MEM_stage_inst_dmem_n8752), .A2(MEM_stage_inst_dmem_n8751), .ZN(MEM_stage_inst_dmem_n12766) );
NAND2_X1 MEM_stage_inst_dmem_U8965 ( .A1(MEM_stage_inst_dmem_n13064), .A2(MEM_stage_inst_dmem_n8758), .ZN(MEM_stage_inst_dmem_n8751) );
NAND2_X1 MEM_stage_inst_dmem_U8964 ( .A1(MEM_stage_inst_dmem_ram_419), .A2(MEM_stage_inst_dmem_n8757), .ZN(MEM_stage_inst_dmem_n8752) );
NAND2_X1 MEM_stage_inst_dmem_U8963 ( .A1(MEM_stage_inst_dmem_n8750), .A2(MEM_stage_inst_dmem_n8749), .ZN(MEM_stage_inst_dmem_n12767) );
NAND2_X1 MEM_stage_inst_dmem_U8962 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n8758), .ZN(MEM_stage_inst_dmem_n8749) );
NAND2_X1 MEM_stage_inst_dmem_U8961 ( .A1(MEM_stage_inst_dmem_ram_420), .A2(MEM_stage_inst_dmem_n8757), .ZN(MEM_stage_inst_dmem_n8750) );
NAND2_X1 MEM_stage_inst_dmem_U8960 ( .A1(MEM_stage_inst_dmem_n8748), .A2(MEM_stage_inst_dmem_n8747), .ZN(MEM_stage_inst_dmem_n12768) );
NAND2_X1 MEM_stage_inst_dmem_U8959 ( .A1(MEM_stage_inst_dmem_n13059), .A2(MEM_stage_inst_dmem_n8758), .ZN(MEM_stage_inst_dmem_n8747) );
NAND2_X1 MEM_stage_inst_dmem_U8958 ( .A1(MEM_stage_inst_dmem_ram_421), .A2(MEM_stage_inst_dmem_n8757), .ZN(MEM_stage_inst_dmem_n8748) );
NAND2_X1 MEM_stage_inst_dmem_U8957 ( .A1(MEM_stage_inst_dmem_n8746), .A2(MEM_stage_inst_dmem_n8745), .ZN(MEM_stage_inst_dmem_n12769) );
NAND2_X1 MEM_stage_inst_dmem_U8956 ( .A1(MEM_stage_inst_dmem_n13056), .A2(MEM_stage_inst_dmem_n8758), .ZN(MEM_stage_inst_dmem_n8745) );
NAND2_X1 MEM_stage_inst_dmem_U8955 ( .A1(MEM_stage_inst_dmem_ram_422), .A2(MEM_stage_inst_dmem_n8757), .ZN(MEM_stage_inst_dmem_n8746) );
NAND2_X1 MEM_stage_inst_dmem_U8954 ( .A1(MEM_stage_inst_dmem_n8744), .A2(MEM_stage_inst_dmem_n8743), .ZN(MEM_stage_inst_dmem_n12770) );
NAND2_X1 MEM_stage_inst_dmem_U8953 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n8758), .ZN(MEM_stage_inst_dmem_n8743) );
NAND2_X1 MEM_stage_inst_dmem_U8952 ( .A1(MEM_stage_inst_dmem_ram_423), .A2(MEM_stage_inst_dmem_n8757), .ZN(MEM_stage_inst_dmem_n8744) );
NAND2_X1 MEM_stage_inst_dmem_U8951 ( .A1(MEM_stage_inst_dmem_n8742), .A2(MEM_stage_inst_dmem_n8741), .ZN(MEM_stage_inst_dmem_n12771) );
NAND2_X1 MEM_stage_inst_dmem_U8950 ( .A1(MEM_stage_inst_dmem_n13051), .A2(MEM_stage_inst_dmem_n8758), .ZN(MEM_stage_inst_dmem_n8741) );
NAND2_X1 MEM_stage_inst_dmem_U8949 ( .A1(MEM_stage_inst_dmem_ram_424), .A2(MEM_stage_inst_dmem_n8757), .ZN(MEM_stage_inst_dmem_n8742) );
NAND2_X1 MEM_stage_inst_dmem_U8948 ( .A1(MEM_stage_inst_dmem_n8740), .A2(MEM_stage_inst_dmem_n8739), .ZN(MEM_stage_inst_dmem_n12772) );
NAND2_X1 MEM_stage_inst_dmem_U8947 ( .A1(MEM_stage_inst_dmem_n19251), .A2(MEM_stage_inst_dmem_n8758), .ZN(MEM_stage_inst_dmem_n8739) );
NAND2_X1 MEM_stage_inst_dmem_U8946 ( .A1(MEM_stage_inst_dmem_ram_425), .A2(MEM_stage_inst_dmem_n8757), .ZN(MEM_stage_inst_dmem_n8740) );
NAND2_X1 MEM_stage_inst_dmem_U8945 ( .A1(MEM_stage_inst_dmem_n8738), .A2(MEM_stage_inst_dmem_n8737), .ZN(MEM_stage_inst_dmem_n12773) );
NAND2_X1 MEM_stage_inst_dmem_U8944 ( .A1(MEM_stage_inst_dmem_n16769), .A2(MEM_stage_inst_dmem_n8758), .ZN(MEM_stage_inst_dmem_n8737) );
NAND2_X1 MEM_stage_inst_dmem_U8943 ( .A1(MEM_stage_inst_dmem_ram_426), .A2(MEM_stage_inst_dmem_n8757), .ZN(MEM_stage_inst_dmem_n8738) );
NAND2_X1 MEM_stage_inst_dmem_U8942 ( .A1(MEM_stage_inst_dmem_n8736), .A2(MEM_stage_inst_dmem_n8735), .ZN(MEM_stage_inst_dmem_n12774) );
NAND2_X1 MEM_stage_inst_dmem_U8941 ( .A1(MEM_stage_inst_dmem_n13044), .A2(MEM_stage_inst_dmem_n8758), .ZN(MEM_stage_inst_dmem_n8735) );
NAND2_X1 MEM_stage_inst_dmem_U8940 ( .A1(MEM_stage_inst_dmem_ram_427), .A2(MEM_stage_inst_dmem_n8757), .ZN(MEM_stage_inst_dmem_n8736) );
NAND2_X1 MEM_stage_inst_dmem_U8939 ( .A1(MEM_stage_inst_dmem_n8734), .A2(MEM_stage_inst_dmem_n8733), .ZN(MEM_stage_inst_dmem_n12775) );
NAND2_X1 MEM_stage_inst_dmem_U8938 ( .A1(MEM_stage_inst_dmem_n13041), .A2(MEM_stage_inst_dmem_n8758), .ZN(MEM_stage_inst_dmem_n8733) );
NAND2_X1 MEM_stage_inst_dmem_U8937 ( .A1(MEM_stage_inst_dmem_ram_428), .A2(MEM_stage_inst_dmem_n8757), .ZN(MEM_stage_inst_dmem_n8734) );
NAND2_X1 MEM_stage_inst_dmem_U8936 ( .A1(MEM_stage_inst_dmem_n8732), .A2(MEM_stage_inst_dmem_n8731), .ZN(MEM_stage_inst_dmem_n12776) );
NAND2_X1 MEM_stage_inst_dmem_U8935 ( .A1(EX_pipeline_reg_out_18), .A2(MEM_stage_inst_dmem_n8758), .ZN(MEM_stage_inst_dmem_n8731) );
NAND2_X1 MEM_stage_inst_dmem_U8934 ( .A1(MEM_stage_inst_dmem_ram_429), .A2(MEM_stage_inst_dmem_n8757), .ZN(MEM_stage_inst_dmem_n8732) );
NAND2_X1 MEM_stage_inst_dmem_U8933 ( .A1(MEM_stage_inst_dmem_n8730), .A2(MEM_stage_inst_dmem_n8729), .ZN(MEM_stage_inst_dmem_n12777) );
NAND2_X1 MEM_stage_inst_dmem_U8932 ( .A1(EX_pipeline_reg_out_19), .A2(MEM_stage_inst_dmem_n8758), .ZN(MEM_stage_inst_dmem_n8729) );
NAND2_X1 MEM_stage_inst_dmem_U8931 ( .A1(MEM_stage_inst_dmem_ram_430), .A2(MEM_stage_inst_dmem_n8757), .ZN(MEM_stage_inst_dmem_n8730) );
NAND2_X1 MEM_stage_inst_dmem_U8930 ( .A1(MEM_stage_inst_dmem_n8728), .A2(MEM_stage_inst_dmem_n8727), .ZN(MEM_stage_inst_dmem_n12778) );
NAND2_X1 MEM_stage_inst_dmem_U8929 ( .A1(EX_pipeline_reg_out_20), .A2(MEM_stage_inst_dmem_n8758), .ZN(MEM_stage_inst_dmem_n8727) );
INV_X1 MEM_stage_inst_dmem_U8928 ( .A(MEM_stage_inst_dmem_n8757), .ZN(MEM_stage_inst_dmem_n8758) );
NAND2_X1 MEM_stage_inst_dmem_U8927 ( .A1(MEM_stage_inst_dmem_ram_431), .A2(MEM_stage_inst_dmem_n8757), .ZN(MEM_stage_inst_dmem_n8728) );
NAND2_X1 MEM_stage_inst_dmem_U8926 ( .A1(MEM_stage_inst_dmem_n13182), .A2(MEM_stage_inst_dmem_n21109), .ZN(MEM_stage_inst_dmem_n8757) );
NOR2_X2 MEM_stage_inst_dmem_U8925 ( .A1(MEM_stage_inst_dmem_n12894), .A2(MEM_stage_inst_dmem_n13110), .ZN(MEM_stage_inst_dmem_n21109) );
NAND2_X1 MEM_stage_inst_dmem_U8924 ( .A1(MEM_stage_inst_dmem_n8726), .A2(MEM_stage_inst_dmem_n8725), .ZN(MEM_stage_inst_dmem_n12779) );
NAND2_X1 MEM_stage_inst_dmem_U8923 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n8724), .ZN(MEM_stage_inst_dmem_n8725) );
NAND2_X1 MEM_stage_inst_dmem_U8922 ( .A1(MEM_stage_inst_dmem_ram_432), .A2(MEM_stage_inst_dmem_n8723), .ZN(MEM_stage_inst_dmem_n8726) );
NAND2_X1 MEM_stage_inst_dmem_U8921 ( .A1(MEM_stage_inst_dmem_n8722), .A2(MEM_stage_inst_dmem_n8721), .ZN(MEM_stage_inst_dmem_n12780) );
NAND2_X1 MEM_stage_inst_dmem_U8920 ( .A1(MEM_stage_inst_dmem_n109), .A2(MEM_stage_inst_dmem_n8724), .ZN(MEM_stage_inst_dmem_n8721) );
NAND2_X1 MEM_stage_inst_dmem_U8919 ( .A1(MEM_stage_inst_dmem_ram_433), .A2(MEM_stage_inst_dmem_n8723), .ZN(MEM_stage_inst_dmem_n8722) );
NAND2_X1 MEM_stage_inst_dmem_U8918 ( .A1(MEM_stage_inst_dmem_n8720), .A2(MEM_stage_inst_dmem_n8719), .ZN(MEM_stage_inst_dmem_n12781) );
NAND2_X1 MEM_stage_inst_dmem_U8917 ( .A1(MEM_stage_inst_dmem_n13900), .A2(MEM_stage_inst_dmem_n8724), .ZN(MEM_stage_inst_dmem_n8719) );
NAND2_X1 MEM_stage_inst_dmem_U8916 ( .A1(MEM_stage_inst_dmem_ram_434), .A2(MEM_stage_inst_dmem_n8723), .ZN(MEM_stage_inst_dmem_n8720) );
NAND2_X1 MEM_stage_inst_dmem_U8915 ( .A1(MEM_stage_inst_dmem_n8718), .A2(MEM_stage_inst_dmem_n8717), .ZN(MEM_stage_inst_dmem_n12782) );
NAND2_X1 MEM_stage_inst_dmem_U8914 ( .A1(MEM_stage_inst_dmem_n13064), .A2(MEM_stage_inst_dmem_n8724), .ZN(MEM_stage_inst_dmem_n8717) );
NAND2_X1 MEM_stage_inst_dmem_U8913 ( .A1(MEM_stage_inst_dmem_ram_435), .A2(MEM_stage_inst_dmem_n8723), .ZN(MEM_stage_inst_dmem_n8718) );
NAND2_X1 MEM_stage_inst_dmem_U8912 ( .A1(MEM_stage_inst_dmem_n8716), .A2(MEM_stage_inst_dmem_n8715), .ZN(MEM_stage_inst_dmem_n12783) );
NAND2_X1 MEM_stage_inst_dmem_U8911 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n8724), .ZN(MEM_stage_inst_dmem_n8715) );
NAND2_X1 MEM_stage_inst_dmem_U8910 ( .A1(MEM_stage_inst_dmem_ram_436), .A2(MEM_stage_inst_dmem_n8723), .ZN(MEM_stage_inst_dmem_n8716) );
NAND2_X1 MEM_stage_inst_dmem_U8909 ( .A1(MEM_stage_inst_dmem_n8714), .A2(MEM_stage_inst_dmem_n8713), .ZN(MEM_stage_inst_dmem_n12784) );
NAND2_X1 MEM_stage_inst_dmem_U8908 ( .A1(MEM_stage_inst_dmem_n13059), .A2(MEM_stage_inst_dmem_n8724), .ZN(MEM_stage_inst_dmem_n8713) );
NAND2_X1 MEM_stage_inst_dmem_U8907 ( .A1(MEM_stage_inst_dmem_ram_437), .A2(MEM_stage_inst_dmem_n8723), .ZN(MEM_stage_inst_dmem_n8714) );
NAND2_X1 MEM_stage_inst_dmem_U8906 ( .A1(MEM_stage_inst_dmem_n8712), .A2(MEM_stage_inst_dmem_n8711), .ZN(MEM_stage_inst_dmem_n12785) );
NAND2_X1 MEM_stage_inst_dmem_U8905 ( .A1(MEM_stage_inst_dmem_n13056), .A2(MEM_stage_inst_dmem_n8724), .ZN(MEM_stage_inst_dmem_n8711) );
NAND2_X1 MEM_stage_inst_dmem_U8904 ( .A1(MEM_stage_inst_dmem_ram_438), .A2(MEM_stage_inst_dmem_n8723), .ZN(MEM_stage_inst_dmem_n8712) );
NAND2_X1 MEM_stage_inst_dmem_U8903 ( .A1(MEM_stage_inst_dmem_n8710), .A2(MEM_stage_inst_dmem_n8709), .ZN(MEM_stage_inst_dmem_n12786) );
NAND2_X1 MEM_stage_inst_dmem_U8902 ( .A1(MEM_stage_inst_dmem_n17), .A2(MEM_stage_inst_dmem_n8724), .ZN(MEM_stage_inst_dmem_n8709) );
NAND2_X1 MEM_stage_inst_dmem_U8901 ( .A1(MEM_stage_inst_dmem_ram_439), .A2(MEM_stage_inst_dmem_n8723), .ZN(MEM_stage_inst_dmem_n8710) );
NAND2_X1 MEM_stage_inst_dmem_U8900 ( .A1(MEM_stage_inst_dmem_n8708), .A2(MEM_stage_inst_dmem_n8707), .ZN(MEM_stage_inst_dmem_n12787) );
NAND2_X1 MEM_stage_inst_dmem_U8899 ( .A1(MEM_stage_inst_dmem_n13051), .A2(MEM_stage_inst_dmem_n8724), .ZN(MEM_stage_inst_dmem_n8707) );
NAND2_X1 MEM_stage_inst_dmem_U8898 ( .A1(MEM_stage_inst_dmem_ram_440), .A2(MEM_stage_inst_dmem_n8723), .ZN(MEM_stage_inst_dmem_n8708) );
NAND2_X1 MEM_stage_inst_dmem_U8897 ( .A1(MEM_stage_inst_dmem_n8706), .A2(MEM_stage_inst_dmem_n8705), .ZN(MEM_stage_inst_dmem_n12788) );
NAND2_X1 MEM_stage_inst_dmem_U8896 ( .A1(MEM_stage_inst_dmem_n20524), .A2(MEM_stage_inst_dmem_n8724), .ZN(MEM_stage_inst_dmem_n8705) );
NAND2_X1 MEM_stage_inst_dmem_U8895 ( .A1(MEM_stage_inst_dmem_ram_441), .A2(MEM_stage_inst_dmem_n8723), .ZN(MEM_stage_inst_dmem_n8706) );
NAND2_X1 MEM_stage_inst_dmem_U8894 ( .A1(MEM_stage_inst_dmem_n8704), .A2(MEM_stage_inst_dmem_n8703), .ZN(MEM_stage_inst_dmem_n12789) );
NAND2_X1 MEM_stage_inst_dmem_U8893 ( .A1(MEM_stage_inst_dmem_n16354), .A2(MEM_stage_inst_dmem_n8724), .ZN(MEM_stage_inst_dmem_n8703) );
NAND2_X1 MEM_stage_inst_dmem_U8892 ( .A1(MEM_stage_inst_dmem_ram_442), .A2(MEM_stage_inst_dmem_n8723), .ZN(MEM_stage_inst_dmem_n8704) );
NAND2_X1 MEM_stage_inst_dmem_U8891 ( .A1(MEM_stage_inst_dmem_n8702), .A2(MEM_stage_inst_dmem_n8701), .ZN(MEM_stage_inst_dmem_n12790) );
NAND2_X1 MEM_stage_inst_dmem_U8890 ( .A1(MEM_stage_inst_dmem_n13044), .A2(MEM_stage_inst_dmem_n8724), .ZN(MEM_stage_inst_dmem_n8701) );
NAND2_X1 MEM_stage_inst_dmem_U8889 ( .A1(MEM_stage_inst_dmem_ram_443), .A2(MEM_stage_inst_dmem_n8723), .ZN(MEM_stage_inst_dmem_n8702) );
NAND2_X1 MEM_stage_inst_dmem_U8888 ( .A1(MEM_stage_inst_dmem_n8700), .A2(MEM_stage_inst_dmem_n8699), .ZN(MEM_stage_inst_dmem_n12791) );
NAND2_X1 MEM_stage_inst_dmem_U8887 ( .A1(MEM_stage_inst_dmem_n13041), .A2(MEM_stage_inst_dmem_n8724), .ZN(MEM_stage_inst_dmem_n8699) );
NAND2_X1 MEM_stage_inst_dmem_U8886 ( .A1(MEM_stage_inst_dmem_ram_444), .A2(MEM_stage_inst_dmem_n8723), .ZN(MEM_stage_inst_dmem_n8700) );
NAND2_X1 MEM_stage_inst_dmem_U8885 ( .A1(MEM_stage_inst_dmem_n8698), .A2(MEM_stage_inst_dmem_n8697), .ZN(MEM_stage_inst_dmem_n12792) );
NAND2_X1 MEM_stage_inst_dmem_U8884 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n8724), .ZN(MEM_stage_inst_dmem_n8697) );
NAND2_X1 MEM_stage_inst_dmem_U8883 ( .A1(MEM_stage_inst_dmem_ram_445), .A2(MEM_stage_inst_dmem_n8723), .ZN(MEM_stage_inst_dmem_n8698) );
NAND2_X1 MEM_stage_inst_dmem_U8882 ( .A1(MEM_stage_inst_dmem_n8696), .A2(MEM_stage_inst_dmem_n8695), .ZN(MEM_stage_inst_dmem_n12793) );
NAND2_X1 MEM_stage_inst_dmem_U8881 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n8724), .ZN(MEM_stage_inst_dmem_n8695) );
NAND2_X1 MEM_stage_inst_dmem_U8880 ( .A1(MEM_stage_inst_dmem_ram_446), .A2(MEM_stage_inst_dmem_n8723), .ZN(MEM_stage_inst_dmem_n8696) );
NAND2_X1 MEM_stage_inst_dmem_U8879 ( .A1(MEM_stage_inst_dmem_n8694), .A2(MEM_stage_inst_dmem_n8693), .ZN(MEM_stage_inst_dmem_n12794) );
NAND2_X1 MEM_stage_inst_dmem_U8878 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n8724), .ZN(MEM_stage_inst_dmem_n8693) );
INV_X1 MEM_stage_inst_dmem_U8877 ( .A(MEM_stage_inst_dmem_n8723), .ZN(MEM_stage_inst_dmem_n8724) );
NAND2_X1 MEM_stage_inst_dmem_U8876 ( .A1(MEM_stage_inst_dmem_ram_447), .A2(MEM_stage_inst_dmem_n8723), .ZN(MEM_stage_inst_dmem_n8694) );
NAND2_X1 MEM_stage_inst_dmem_U8875 ( .A1(MEM_stage_inst_dmem_n13182), .A2(MEM_stage_inst_dmem_n21074), .ZN(MEM_stage_inst_dmem_n8723) );
NOR2_X2 MEM_stage_inst_dmem_U8874 ( .A1(MEM_stage_inst_dmem_n12859), .A2(MEM_stage_inst_dmem_n13110), .ZN(MEM_stage_inst_dmem_n21074) );
NAND2_X1 MEM_stage_inst_dmem_U8873 ( .A1(EX_pipeline_reg_out_23), .A2(MEM_stage_inst_dmem_n8762), .ZN(MEM_stage_inst_dmem_n13110) );
NAND2_X1 MEM_stage_inst_dmem_U8872 ( .A1(MEM_stage_inst_dmem_n8692), .A2(MEM_stage_inst_dmem_n8691), .ZN(MEM_stage_inst_dmem_n12795) );
NAND2_X1 MEM_stage_inst_dmem_U8871 ( .A1(MEM_stage_inst_dmem_n21501), .A2(MEM_stage_inst_dmem_n8690), .ZN(MEM_stage_inst_dmem_n8691) );
NAND2_X1 MEM_stage_inst_dmem_U8870 ( .A1(MEM_stage_inst_dmem_ram_448), .A2(MEM_stage_inst_dmem_n8689), .ZN(MEM_stage_inst_dmem_n8692) );
NAND2_X1 MEM_stage_inst_dmem_U8869 ( .A1(MEM_stage_inst_dmem_n8688), .A2(MEM_stage_inst_dmem_n8687), .ZN(MEM_stage_inst_dmem_n12796) );
NAND2_X1 MEM_stage_inst_dmem_U8868 ( .A1(MEM_stage_inst_dmem_n109), .A2(MEM_stage_inst_dmem_n8690), .ZN(MEM_stage_inst_dmem_n8687) );
NAND2_X1 MEM_stage_inst_dmem_U8867 ( .A1(MEM_stage_inst_dmem_ram_449), .A2(MEM_stage_inst_dmem_n8689), .ZN(MEM_stage_inst_dmem_n8688) );
NAND2_X1 MEM_stage_inst_dmem_U8866 ( .A1(MEM_stage_inst_dmem_n8686), .A2(MEM_stage_inst_dmem_n8685), .ZN(MEM_stage_inst_dmem_n12797) );
NAND2_X1 MEM_stage_inst_dmem_U8865 ( .A1(MEM_stage_inst_dmem_n16373), .A2(MEM_stage_inst_dmem_n8690), .ZN(MEM_stage_inst_dmem_n8685) );
NAND2_X1 MEM_stage_inst_dmem_U8864 ( .A1(MEM_stage_inst_dmem_ram_450), .A2(MEM_stage_inst_dmem_n8689), .ZN(MEM_stage_inst_dmem_n8686) );
NAND2_X1 MEM_stage_inst_dmem_U8863 ( .A1(MEM_stage_inst_dmem_n8684), .A2(MEM_stage_inst_dmem_n8683), .ZN(MEM_stage_inst_dmem_n12798) );
NAND2_X1 MEM_stage_inst_dmem_U8862 ( .A1(MEM_stage_inst_dmem_n13064), .A2(MEM_stage_inst_dmem_n8690), .ZN(MEM_stage_inst_dmem_n8683) );
NAND2_X1 MEM_stage_inst_dmem_U8861 ( .A1(MEM_stage_inst_dmem_ram_451), .A2(MEM_stage_inst_dmem_n8689), .ZN(MEM_stage_inst_dmem_n8684) );
NAND2_X1 MEM_stage_inst_dmem_U8860 ( .A1(MEM_stage_inst_dmem_n8682), .A2(MEM_stage_inst_dmem_n8681), .ZN(MEM_stage_inst_dmem_n12799) );
NAND2_X1 MEM_stage_inst_dmem_U8859 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n8690), .ZN(MEM_stage_inst_dmem_n8681) );
NAND2_X1 MEM_stage_inst_dmem_U8858 ( .A1(MEM_stage_inst_dmem_ram_452), .A2(MEM_stage_inst_dmem_n8689), .ZN(MEM_stage_inst_dmem_n8682) );
NAND2_X1 MEM_stage_inst_dmem_U8857 ( .A1(MEM_stage_inst_dmem_n8680), .A2(MEM_stage_inst_dmem_n8679), .ZN(MEM_stage_inst_dmem_n12800) );
NAND2_X1 MEM_stage_inst_dmem_U8856 ( .A1(MEM_stage_inst_dmem_n13059), .A2(MEM_stage_inst_dmem_n8690), .ZN(MEM_stage_inst_dmem_n8679) );
NAND2_X1 MEM_stage_inst_dmem_U8855 ( .A1(MEM_stage_inst_dmem_ram_453), .A2(MEM_stage_inst_dmem_n8689), .ZN(MEM_stage_inst_dmem_n8680) );
NAND2_X1 MEM_stage_inst_dmem_U8854 ( .A1(MEM_stage_inst_dmem_n8678), .A2(MEM_stage_inst_dmem_n8677), .ZN(MEM_stage_inst_dmem_n12801) );
NAND2_X1 MEM_stage_inst_dmem_U8853 ( .A1(MEM_stage_inst_dmem_n13056), .A2(MEM_stage_inst_dmem_n8690), .ZN(MEM_stage_inst_dmem_n8677) );
NAND2_X1 MEM_stage_inst_dmem_U8852 ( .A1(MEM_stage_inst_dmem_ram_454), .A2(MEM_stage_inst_dmem_n8689), .ZN(MEM_stage_inst_dmem_n8678) );
NAND2_X1 MEM_stage_inst_dmem_U8851 ( .A1(MEM_stage_inst_dmem_n8676), .A2(MEM_stage_inst_dmem_n8675), .ZN(MEM_stage_inst_dmem_n12802) );
NAND2_X1 MEM_stage_inst_dmem_U8850 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n8690), .ZN(MEM_stage_inst_dmem_n8675) );
NAND2_X1 MEM_stage_inst_dmem_U8849 ( .A1(MEM_stage_inst_dmem_ram_455), .A2(MEM_stage_inst_dmem_n8689), .ZN(MEM_stage_inst_dmem_n8676) );
NAND2_X1 MEM_stage_inst_dmem_U8848 ( .A1(MEM_stage_inst_dmem_n8674), .A2(MEM_stage_inst_dmem_n8673), .ZN(MEM_stage_inst_dmem_n12803) );
NAND2_X1 MEM_stage_inst_dmem_U8847 ( .A1(MEM_stage_inst_dmem_n13051), .A2(MEM_stage_inst_dmem_n8690), .ZN(MEM_stage_inst_dmem_n8673) );
NAND2_X1 MEM_stage_inst_dmem_U8846 ( .A1(MEM_stage_inst_dmem_ram_456), .A2(MEM_stage_inst_dmem_n8689), .ZN(MEM_stage_inst_dmem_n8674) );
NAND2_X1 MEM_stage_inst_dmem_U8845 ( .A1(MEM_stage_inst_dmem_n8672), .A2(MEM_stage_inst_dmem_n8671), .ZN(MEM_stage_inst_dmem_n12804) );
NAND2_X1 MEM_stage_inst_dmem_U8844 ( .A1(EX_pipeline_reg_out_14), .A2(MEM_stage_inst_dmem_n8690), .ZN(MEM_stage_inst_dmem_n8671) );
NAND2_X1 MEM_stage_inst_dmem_U8843 ( .A1(MEM_stage_inst_dmem_ram_457), .A2(MEM_stage_inst_dmem_n8689), .ZN(MEM_stage_inst_dmem_n8672) );
NAND2_X1 MEM_stage_inst_dmem_U8842 ( .A1(MEM_stage_inst_dmem_n8670), .A2(MEM_stage_inst_dmem_n8669), .ZN(MEM_stage_inst_dmem_n12805) );
NAND2_X1 MEM_stage_inst_dmem_U8841 ( .A1(MEM_stage_inst_dmem_n18867), .A2(MEM_stage_inst_dmem_n8690), .ZN(MEM_stage_inst_dmem_n8669) );
NAND2_X1 MEM_stage_inst_dmem_U8840 ( .A1(MEM_stage_inst_dmem_ram_458), .A2(MEM_stage_inst_dmem_n8689), .ZN(MEM_stage_inst_dmem_n8670) );
NAND2_X1 MEM_stage_inst_dmem_U8839 ( .A1(MEM_stage_inst_dmem_n8668), .A2(MEM_stage_inst_dmem_n8667), .ZN(MEM_stage_inst_dmem_n12806) );
NAND2_X1 MEM_stage_inst_dmem_U8838 ( .A1(MEM_stage_inst_dmem_n13044), .A2(MEM_stage_inst_dmem_n8690), .ZN(MEM_stage_inst_dmem_n8667) );
NAND2_X1 MEM_stage_inst_dmem_U8837 ( .A1(MEM_stage_inst_dmem_ram_459), .A2(MEM_stage_inst_dmem_n8689), .ZN(MEM_stage_inst_dmem_n8668) );
NAND2_X1 MEM_stage_inst_dmem_U8836 ( .A1(MEM_stage_inst_dmem_n8666), .A2(MEM_stage_inst_dmem_n8665), .ZN(MEM_stage_inst_dmem_n12807) );
NAND2_X1 MEM_stage_inst_dmem_U8835 ( .A1(MEM_stage_inst_dmem_n13041), .A2(MEM_stage_inst_dmem_n8690), .ZN(MEM_stage_inst_dmem_n8665) );
NAND2_X1 MEM_stage_inst_dmem_U8834 ( .A1(MEM_stage_inst_dmem_ram_460), .A2(MEM_stage_inst_dmem_n8689), .ZN(MEM_stage_inst_dmem_n8666) );
NAND2_X1 MEM_stage_inst_dmem_U8833 ( .A1(MEM_stage_inst_dmem_n8664), .A2(MEM_stage_inst_dmem_n8663), .ZN(MEM_stage_inst_dmem_n12808) );
NAND2_X1 MEM_stage_inst_dmem_U8832 ( .A1(MEM_stage_inst_dmem_n21471), .A2(MEM_stage_inst_dmem_n8690), .ZN(MEM_stage_inst_dmem_n8663) );
NAND2_X1 MEM_stage_inst_dmem_U8831 ( .A1(MEM_stage_inst_dmem_ram_461), .A2(MEM_stage_inst_dmem_n8689), .ZN(MEM_stage_inst_dmem_n8664) );
NAND2_X1 MEM_stage_inst_dmem_U8830 ( .A1(MEM_stage_inst_dmem_n8662), .A2(MEM_stage_inst_dmem_n8661), .ZN(MEM_stage_inst_dmem_n12809) );
NAND2_X1 MEM_stage_inst_dmem_U8829 ( .A1(MEM_stage_inst_dmem_n21468), .A2(MEM_stage_inst_dmem_n8690), .ZN(MEM_stage_inst_dmem_n8661) );
NAND2_X1 MEM_stage_inst_dmem_U8828 ( .A1(MEM_stage_inst_dmem_ram_462), .A2(MEM_stage_inst_dmem_n8689), .ZN(MEM_stage_inst_dmem_n8662) );
NAND2_X1 MEM_stage_inst_dmem_U8827 ( .A1(MEM_stage_inst_dmem_n8660), .A2(MEM_stage_inst_dmem_n8659), .ZN(MEM_stage_inst_dmem_n12810) );
NAND2_X1 MEM_stage_inst_dmem_U8826 ( .A1(MEM_stage_inst_dmem_n14693), .A2(MEM_stage_inst_dmem_n8690), .ZN(MEM_stage_inst_dmem_n8659) );
INV_X1 MEM_stage_inst_dmem_U8825 ( .A(MEM_stage_inst_dmem_n8689), .ZN(MEM_stage_inst_dmem_n8690) );
NAND2_X1 MEM_stage_inst_dmem_U8824 ( .A1(MEM_stage_inst_dmem_ram_463), .A2(MEM_stage_inst_dmem_n8689), .ZN(MEM_stage_inst_dmem_n8660) );
NAND2_X1 MEM_stage_inst_dmem_U8823 ( .A1(MEM_stage_inst_dmem_n13182), .A2(MEM_stage_inst_dmem_n21039), .ZN(MEM_stage_inst_dmem_n8689) );
NOR2_X2 MEM_stage_inst_dmem_U8822 ( .A1(MEM_stage_inst_dmem_n12894), .A2(MEM_stage_inst_dmem_n13034), .ZN(MEM_stage_inst_dmem_n21039) );
NAND2_X1 MEM_stage_inst_dmem_U8821 ( .A1(MEM_stage_inst_dmem_n8658), .A2(MEM_stage_inst_dmem_n8657), .ZN(MEM_stage_inst_dmem_n12811) );
NAND2_X1 MEM_stage_inst_dmem_U8820 ( .A1(MEM_stage_inst_dmem_n8), .A2(MEM_stage_inst_dmem_n8656), .ZN(MEM_stage_inst_dmem_n8657) );
NAND2_X1 MEM_stage_inst_dmem_U8819 ( .A1(MEM_stage_inst_dmem_ram_464), .A2(MEM_stage_inst_dmem_n8655), .ZN(MEM_stage_inst_dmem_n8658) );
NAND2_X1 MEM_stage_inst_dmem_U8818 ( .A1(MEM_stage_inst_dmem_n8654), .A2(MEM_stage_inst_dmem_n8653), .ZN(MEM_stage_inst_dmem_n12812) );
NAND2_X1 MEM_stage_inst_dmem_U8817 ( .A1(MEM_stage_inst_dmem_n109), .A2(MEM_stage_inst_dmem_n8656), .ZN(MEM_stage_inst_dmem_n8653) );
NAND2_X1 MEM_stage_inst_dmem_U8816 ( .A1(MEM_stage_inst_dmem_ram_465), .A2(MEM_stage_inst_dmem_n8655), .ZN(MEM_stage_inst_dmem_n8654) );
NAND2_X1 MEM_stage_inst_dmem_U8815 ( .A1(MEM_stage_inst_dmem_n8652), .A2(MEM_stage_inst_dmem_n8651), .ZN(MEM_stage_inst_dmem_n12813) );
NAND2_X1 MEM_stage_inst_dmem_U8814 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n8656), .ZN(MEM_stage_inst_dmem_n8651) );
NAND2_X1 MEM_stage_inst_dmem_U8813 ( .A1(MEM_stage_inst_dmem_ram_466), .A2(MEM_stage_inst_dmem_n8655), .ZN(MEM_stage_inst_dmem_n8652) );
NAND2_X1 MEM_stage_inst_dmem_U8812 ( .A1(MEM_stage_inst_dmem_n8650), .A2(MEM_stage_inst_dmem_n8649), .ZN(MEM_stage_inst_dmem_n12814) );
NAND2_X1 MEM_stage_inst_dmem_U8811 ( .A1(MEM_stage_inst_dmem_n13064), .A2(MEM_stage_inst_dmem_n8656), .ZN(MEM_stage_inst_dmem_n8649) );
NAND2_X1 MEM_stage_inst_dmem_U8810 ( .A1(MEM_stage_inst_dmem_ram_467), .A2(MEM_stage_inst_dmem_n8655), .ZN(MEM_stage_inst_dmem_n8650) );
NAND2_X1 MEM_stage_inst_dmem_U8809 ( .A1(MEM_stage_inst_dmem_n8648), .A2(MEM_stage_inst_dmem_n8647), .ZN(MEM_stage_inst_dmem_n12815) );
NAND2_X1 MEM_stage_inst_dmem_U8808 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n8656), .ZN(MEM_stage_inst_dmem_n8647) );
NAND2_X1 MEM_stage_inst_dmem_U8807 ( .A1(MEM_stage_inst_dmem_ram_468), .A2(MEM_stage_inst_dmem_n8655), .ZN(MEM_stage_inst_dmem_n8648) );
NAND2_X1 MEM_stage_inst_dmem_U8806 ( .A1(MEM_stage_inst_dmem_n8646), .A2(MEM_stage_inst_dmem_n8645), .ZN(MEM_stage_inst_dmem_n12816) );
NAND2_X1 MEM_stage_inst_dmem_U8805 ( .A1(MEM_stage_inst_dmem_n13059), .A2(MEM_stage_inst_dmem_n8656), .ZN(MEM_stage_inst_dmem_n8645) );
NAND2_X1 MEM_stage_inst_dmem_U8804 ( .A1(MEM_stage_inst_dmem_ram_469), .A2(MEM_stage_inst_dmem_n8655), .ZN(MEM_stage_inst_dmem_n8646) );
NAND2_X1 MEM_stage_inst_dmem_U8803 ( .A1(MEM_stage_inst_dmem_n8644), .A2(MEM_stage_inst_dmem_n8643), .ZN(MEM_stage_inst_dmem_n12817) );
NAND2_X1 MEM_stage_inst_dmem_U8802 ( .A1(MEM_stage_inst_dmem_n13056), .A2(MEM_stage_inst_dmem_n8656), .ZN(MEM_stage_inst_dmem_n8643) );
NAND2_X1 MEM_stage_inst_dmem_U8801 ( .A1(MEM_stage_inst_dmem_ram_470), .A2(MEM_stage_inst_dmem_n8655), .ZN(MEM_stage_inst_dmem_n8644) );
NAND2_X1 MEM_stage_inst_dmem_U8800 ( .A1(MEM_stage_inst_dmem_n8642), .A2(MEM_stage_inst_dmem_n8641), .ZN(MEM_stage_inst_dmem_n12818) );
NAND2_X1 MEM_stage_inst_dmem_U8799 ( .A1(MEM_stage_inst_dmem_n101), .A2(MEM_stage_inst_dmem_n8656), .ZN(MEM_stage_inst_dmem_n8641) );
NAND2_X1 MEM_stage_inst_dmem_U8798 ( .A1(MEM_stage_inst_dmem_ram_471), .A2(MEM_stage_inst_dmem_n8655), .ZN(MEM_stage_inst_dmem_n8642) );
NAND2_X1 MEM_stage_inst_dmem_U8797 ( .A1(MEM_stage_inst_dmem_n8640), .A2(MEM_stage_inst_dmem_n8639), .ZN(MEM_stage_inst_dmem_n12819) );
NAND2_X1 MEM_stage_inst_dmem_U8796 ( .A1(MEM_stage_inst_dmem_n13051), .A2(MEM_stage_inst_dmem_n8656), .ZN(MEM_stage_inst_dmem_n8639) );
NAND2_X1 MEM_stage_inst_dmem_U8795 ( .A1(MEM_stage_inst_dmem_ram_472), .A2(MEM_stage_inst_dmem_n8655), .ZN(MEM_stage_inst_dmem_n8640) );
NAND2_X1 MEM_stage_inst_dmem_U8794 ( .A1(MEM_stage_inst_dmem_n8638), .A2(MEM_stage_inst_dmem_n8637), .ZN(MEM_stage_inst_dmem_n12820) );
NAND2_X1 MEM_stage_inst_dmem_U8793 ( .A1(MEM_stage_inst_dmem_n2), .A2(MEM_stage_inst_dmem_n8656), .ZN(MEM_stage_inst_dmem_n8637) );
NAND2_X1 MEM_stage_inst_dmem_U8792 ( .A1(MEM_stage_inst_dmem_ram_473), .A2(MEM_stage_inst_dmem_n8655), .ZN(MEM_stage_inst_dmem_n8638) );
NAND2_X1 MEM_stage_inst_dmem_U8791 ( .A1(MEM_stage_inst_dmem_n8636), .A2(MEM_stage_inst_dmem_n8635), .ZN(MEM_stage_inst_dmem_n12821) );
NAND2_X1 MEM_stage_inst_dmem_U8790 ( .A1(MEM_stage_inst_dmem_n20521), .A2(MEM_stage_inst_dmem_n8656), .ZN(MEM_stage_inst_dmem_n8635) );
NAND2_X1 MEM_stage_inst_dmem_U8789 ( .A1(MEM_stage_inst_dmem_ram_474), .A2(MEM_stage_inst_dmem_n8655), .ZN(MEM_stage_inst_dmem_n8636) );
NAND2_X1 MEM_stage_inst_dmem_U8788 ( .A1(MEM_stage_inst_dmem_n8634), .A2(MEM_stage_inst_dmem_n8633), .ZN(MEM_stage_inst_dmem_n12822) );
NAND2_X1 MEM_stage_inst_dmem_U8787 ( .A1(MEM_stage_inst_dmem_n13044), .A2(MEM_stage_inst_dmem_n8656), .ZN(MEM_stage_inst_dmem_n8633) );
NAND2_X1 MEM_stage_inst_dmem_U8786 ( .A1(MEM_stage_inst_dmem_ram_475), .A2(MEM_stage_inst_dmem_n8655), .ZN(MEM_stage_inst_dmem_n8634) );
NAND2_X1 MEM_stage_inst_dmem_U8785 ( .A1(MEM_stage_inst_dmem_n8632), .A2(MEM_stage_inst_dmem_n8631), .ZN(MEM_stage_inst_dmem_n12823) );
NAND2_X1 MEM_stage_inst_dmem_U8784 ( .A1(MEM_stage_inst_dmem_n13041), .A2(MEM_stage_inst_dmem_n8656), .ZN(MEM_stage_inst_dmem_n8631) );
NAND2_X1 MEM_stage_inst_dmem_U8783 ( .A1(MEM_stage_inst_dmem_ram_476), .A2(MEM_stage_inst_dmem_n8655), .ZN(MEM_stage_inst_dmem_n8632) );
NAND2_X1 MEM_stage_inst_dmem_U8782 ( .A1(MEM_stage_inst_dmem_n8630), .A2(MEM_stage_inst_dmem_n8629), .ZN(MEM_stage_inst_dmem_n12824) );
NAND2_X1 MEM_stage_inst_dmem_U8781 ( .A1(MEM_stage_inst_dmem_n12), .A2(MEM_stage_inst_dmem_n8656), .ZN(MEM_stage_inst_dmem_n8629) );
NAND2_X1 MEM_stage_inst_dmem_U8780 ( .A1(MEM_stage_inst_dmem_ram_477), .A2(MEM_stage_inst_dmem_n8655), .ZN(MEM_stage_inst_dmem_n8630) );
NAND2_X1 MEM_stage_inst_dmem_U8779 ( .A1(MEM_stage_inst_dmem_n8628), .A2(MEM_stage_inst_dmem_n8627), .ZN(MEM_stage_inst_dmem_n12825) );
NAND2_X1 MEM_stage_inst_dmem_U8778 ( .A1(MEM_stage_inst_dmem_n10), .A2(MEM_stage_inst_dmem_n8656), .ZN(MEM_stage_inst_dmem_n8627) );
NAND2_X1 MEM_stage_inst_dmem_U8777 ( .A1(MEM_stage_inst_dmem_ram_478), .A2(MEM_stage_inst_dmem_n8655), .ZN(MEM_stage_inst_dmem_n8628) );
NAND2_X1 MEM_stage_inst_dmem_U8776 ( .A1(MEM_stage_inst_dmem_n8626), .A2(MEM_stage_inst_dmem_n8625), .ZN(MEM_stage_inst_dmem_n12826) );
NAND2_X1 MEM_stage_inst_dmem_U8775 ( .A1(MEM_stage_inst_dmem_n15110), .A2(MEM_stage_inst_dmem_n8656), .ZN(MEM_stage_inst_dmem_n8625) );
NAND2_X1 MEM_stage_inst_dmem_U8774 ( .A1(MEM_stage_inst_dmem_ram_479), .A2(MEM_stage_inst_dmem_n8655), .ZN(MEM_stage_inst_dmem_n8626) );
NAND2_X1 MEM_stage_inst_dmem_U8773 ( .A1(MEM_stage_inst_dmem_n13182), .A2(MEM_stage_inst_dmem_n21004), .ZN(MEM_stage_inst_dmem_n8655) );
NOR2_X2 MEM_stage_inst_dmem_U8772 ( .A1(MEM_stage_inst_dmem_n12859), .A2(MEM_stage_inst_dmem_n13034), .ZN(MEM_stage_inst_dmem_n21004) );
NAND2_X1 MEM_stage_inst_dmem_U8771 ( .A1(EX_pipeline_reg_out_24), .A2(MEM_stage_inst_dmem_n8761), .ZN(MEM_stage_inst_dmem_n13034) );
NAND2_X1 MEM_stage_inst_dmem_U8770 ( .A1(MEM_stage_inst_dmem_n8624), .A2(MEM_stage_inst_dmem_n8623), .ZN(MEM_stage_inst_dmem_n12827) );
NAND2_X1 MEM_stage_inst_dmem_U8769 ( .A1(MEM_stage_inst_dmem_n15145), .A2(MEM_stage_inst_dmem_n8622), .ZN(MEM_stage_inst_dmem_n8623) );
NAND2_X1 MEM_stage_inst_dmem_U8768 ( .A1(MEM_stage_inst_dmem_ram_480), .A2(MEM_stage_inst_dmem_n8621), .ZN(MEM_stage_inst_dmem_n8624) );
NAND2_X1 MEM_stage_inst_dmem_U8767 ( .A1(MEM_stage_inst_dmem_n8620), .A2(MEM_stage_inst_dmem_n8619), .ZN(MEM_stage_inst_dmem_n12828) );
NAND2_X1 MEM_stage_inst_dmem_U8766 ( .A1(MEM_stage_inst_dmem_n109), .A2(MEM_stage_inst_dmem_n8622), .ZN(MEM_stage_inst_dmem_n8619) );
NAND2_X1 MEM_stage_inst_dmem_U8765 ( .A1(MEM_stage_inst_dmem_ram_481), .A2(MEM_stage_inst_dmem_n8621), .ZN(MEM_stage_inst_dmem_n8620) );
NAND2_X1 MEM_stage_inst_dmem_U8764 ( .A1(MEM_stage_inst_dmem_n8618), .A2(MEM_stage_inst_dmem_n8617), .ZN(MEM_stage_inst_dmem_n12829) );
NAND2_X1 MEM_stage_inst_dmem_U8763 ( .A1(MEM_stage_inst_dmem_n113), .A2(MEM_stage_inst_dmem_n8622), .ZN(MEM_stage_inst_dmem_n8617) );
NAND2_X1 MEM_stage_inst_dmem_U8762 ( .A1(MEM_stage_inst_dmem_ram_482), .A2(MEM_stage_inst_dmem_n8621), .ZN(MEM_stage_inst_dmem_n8618) );
NAND2_X1 MEM_stage_inst_dmem_U8761 ( .A1(MEM_stage_inst_dmem_n8616), .A2(MEM_stage_inst_dmem_n8615), .ZN(MEM_stage_inst_dmem_n12830) );
NAND2_X1 MEM_stage_inst_dmem_U8760 ( .A1(MEM_stage_inst_dmem_n13064), .A2(MEM_stage_inst_dmem_n8622), .ZN(MEM_stage_inst_dmem_n8615) );
NAND2_X1 MEM_stage_inst_dmem_U8759 ( .A1(MEM_stage_inst_dmem_ram_483), .A2(MEM_stage_inst_dmem_n8621), .ZN(MEM_stage_inst_dmem_n8616) );
NAND2_X1 MEM_stage_inst_dmem_U8758 ( .A1(MEM_stage_inst_dmem_n8614), .A2(MEM_stage_inst_dmem_n8613), .ZN(MEM_stage_inst_dmem_n12831) );
NAND2_X1 MEM_stage_inst_dmem_U8757 ( .A1(MEM_stage_inst_dmem_n6), .A2(MEM_stage_inst_dmem_n8622), .ZN(MEM_stage_inst_dmem_n8613) );
NAND2_X1 MEM_stage_inst_dmem_U8756 ( .A1(MEM_stage_inst_dmem_ram_484), .A2(MEM_stage_inst_dmem_n8621), .ZN(MEM_stage_inst_dmem_n8614) );
NAND2_X1 MEM_stage_inst_dmem_U8755 ( .A1(MEM_stage_inst_dmem_n8612), .A2(MEM_stage_inst_dmem_n8611), .ZN(MEM_stage_inst_dmem_n12832) );
NAND2_X1 MEM_stage_inst_dmem_U8754 ( .A1(MEM_stage_inst_dmem_n13059), .A2(MEM_stage_inst_dmem_n8622), .ZN(MEM_stage_inst_dmem_n8611) );
NAND2_X1 MEM_stage_inst_dmem_U8753 ( .A1(MEM_stage_inst_dmem_ram_485), .A2(MEM_stage_inst_dmem_n8621), .ZN(MEM_stage_inst_dmem_n8612) );
NAND2_X1 MEM_stage_inst_dmem_U8752 ( .A1(MEM_stage_inst_dmem_n8610), .A2(MEM_stage_inst_dmem_n8609), .ZN(MEM_stage_inst_dmem_n12833) );
NAND2_X1 MEM_stage_inst_dmem_U8751 ( .A1(MEM_stage_inst_dmem_n13056), .A2(MEM_stage_inst_dmem_n8622), .ZN(MEM_stage_inst_dmem_n8609) );
NAND2_X1 MEM_stage_inst_dmem_U8750 ( .A1(MEM_stage_inst_dmem_ram_486), .A2(MEM_stage_inst_dmem_n8621), .ZN(MEM_stage_inst_dmem_n8610) );
NAND2_X1 MEM_stage_inst_dmem_U8749 ( .A1(MEM_stage_inst_dmem_n8608), .A2(MEM_stage_inst_dmem_n8607), .ZN(MEM_stage_inst_dmem_n12834) );
NAND2_X1 MEM_stage_inst_dmem_U8748 ( .A1(MEM_stage_inst_dmem_n16361), .A2(MEM_stage_inst_dmem_n8622), .ZN(MEM_stage_inst_dmem_n8607) );
NAND2_X1 MEM_stage_inst_dmem_U8747 ( .A1(MEM_stage_inst_dmem_ram_487), .A2(MEM_stage_inst_dmem_n8621), .ZN(MEM_stage_inst_dmem_n8608) );
NAND2_X1 MEM_stage_inst_dmem_U8746 ( .A1(MEM_stage_inst_dmem_n8606), .A2(MEM_stage_inst_dmem_n8605), .ZN(MEM_stage_inst_dmem_n12835) );
NAND2_X1 MEM_stage_inst_dmem_U8745 ( .A1(MEM_stage_inst_dmem_n13051), .A2(MEM_stage_inst_dmem_n8622), .ZN(MEM_stage_inst_dmem_n8605) );
NAND2_X1 MEM_stage_inst_dmem_U8744 ( .A1(MEM_stage_inst_dmem_ram_488), .A2(MEM_stage_inst_dmem_n8621), .ZN(MEM_stage_inst_dmem_n8606) );
NAND2_X1 MEM_stage_inst_dmem_U8743 ( .A1(MEM_stage_inst_dmem_n8604), .A2(MEM_stage_inst_dmem_n8603), .ZN(MEM_stage_inst_dmem_n12836) );
NAND2_X1 MEM_stage_inst_dmem_U8742 ( .A1(MEM_stage_inst_dmem_n19251), .A2(MEM_stage_inst_dmem_n8622), .ZN(MEM_stage_inst_dmem_n8603) );
NAND2_X1 MEM_stage_inst_dmem_U8741 ( .A1(MEM_stage_inst_dmem_ram_489), .A2(MEM_stage_inst_dmem_n8621), .ZN(MEM_stage_inst_dmem_n8604) );
NAND2_X1 MEM_stage_inst_dmem_U8740 ( .A1(MEM_stage_inst_dmem_n8602), .A2(MEM_stage_inst_dmem_n8601), .ZN(MEM_stage_inst_dmem_n12837) );
NAND2_X1 MEM_stage_inst_dmem_U8739 ( .A1(EX_pipeline_reg_out_15), .A2(MEM_stage_inst_dmem_n8622), .ZN(MEM_stage_inst_dmem_n8601) );
NAND2_X1 MEM_stage_inst_dmem_U8738 ( .A1(MEM_stage_inst_dmem_ram_490), .A2(MEM_stage_inst_dmem_n8621), .ZN(MEM_stage_inst_dmem_n8602) );
NAND2_X1 MEM_stage_inst_dmem_U8737 ( .A1(MEM_stage_inst_dmem_n8600), .A2(MEM_stage_inst_dmem_n8599), .ZN(MEM_stage_inst_dmem_n12838) );
NAND2_X1 MEM_stage_inst_dmem_U8736 ( .A1(MEM_stage_inst_dmem_n13044), .A2(MEM_stage_inst_dmem_n8622), .ZN(MEM_stage_inst_dmem_n8599) );
NAND2_X1 MEM_stage_inst_dmem_U8735 ( .A1(MEM_stage_inst_dmem_ram_491), .A2(MEM_stage_inst_dmem_n8621), .ZN(MEM_stage_inst_dmem_n8600) );
NAND2_X1 MEM_stage_inst_dmem_U8734 ( .A1(MEM_stage_inst_dmem_n8598), .A2(MEM_stage_inst_dmem_n8597), .ZN(MEM_stage_inst_dmem_n12839) );
NAND2_X1 MEM_stage_inst_dmem_U8733 ( .A1(MEM_stage_inst_dmem_n13041), .A2(MEM_stage_inst_dmem_n8622), .ZN(MEM_stage_inst_dmem_n8597) );
NAND2_X1 MEM_stage_inst_dmem_U8732 ( .A1(MEM_stage_inst_dmem_ram_492), .A2(MEM_stage_inst_dmem_n8621), .ZN(MEM_stage_inst_dmem_n8598) );
NAND2_X1 MEM_stage_inst_dmem_U8731 ( .A1(MEM_stage_inst_dmem_n8596), .A2(MEM_stage_inst_dmem_n8595), .ZN(MEM_stage_inst_dmem_n12840) );
NAND2_X1 MEM_stage_inst_dmem_U8730 ( .A1(MEM_stage_inst_dmem_n15116), .A2(MEM_stage_inst_dmem_n8622), .ZN(MEM_stage_inst_dmem_n8595) );
NAND2_X1 MEM_stage_inst_dmem_U8729 ( .A1(MEM_stage_inst_dmem_ram_493), .A2(MEM_stage_inst_dmem_n8621), .ZN(MEM_stage_inst_dmem_n8596) );
NAND2_X1 MEM_stage_inst_dmem_U8728 ( .A1(MEM_stage_inst_dmem_n8594), .A2(MEM_stage_inst_dmem_n8593), .ZN(MEM_stage_inst_dmem_n12841) );
NAND2_X1 MEM_stage_inst_dmem_U8727 ( .A1(MEM_stage_inst_dmem_n15113), .A2(MEM_stage_inst_dmem_n8622), .ZN(MEM_stage_inst_dmem_n8593) );
NAND2_X1 MEM_stage_inst_dmem_U8726 ( .A1(MEM_stage_inst_dmem_ram_494), .A2(MEM_stage_inst_dmem_n8621), .ZN(MEM_stage_inst_dmem_n8594) );
NAND2_X1 MEM_stage_inst_dmem_U8725 ( .A1(MEM_stage_inst_dmem_n8592), .A2(MEM_stage_inst_dmem_n8591), .ZN(MEM_stage_inst_dmem_n12842) );
NAND2_X1 MEM_stage_inst_dmem_U8724 ( .A1(MEM_stage_inst_dmem_n114), .A2(MEM_stage_inst_dmem_n8622), .ZN(MEM_stage_inst_dmem_n8591) );
INV_X1 MEM_stage_inst_dmem_U8723 ( .A(MEM_stage_inst_dmem_n8621), .ZN(MEM_stage_inst_dmem_n8622) );
NAND2_X1 MEM_stage_inst_dmem_U8722 ( .A1(MEM_stage_inst_dmem_ram_495), .A2(MEM_stage_inst_dmem_n8621), .ZN(MEM_stage_inst_dmem_n8592) );
NAND2_X1 MEM_stage_inst_dmem_U8721 ( .A1(MEM_stage_inst_dmem_n13182), .A2(MEM_stage_inst_dmem_n20969), .ZN(MEM_stage_inst_dmem_n8621) );
NOR2_X2 MEM_stage_inst_dmem_U8720 ( .A1(MEM_stage_inst_dmem_n12965), .A2(MEM_stage_inst_dmem_n12894), .ZN(MEM_stage_inst_dmem_n20969) );
NAND2_X1 MEM_stage_inst_dmem_U8719 ( .A1(EX_pipeline_reg_out_25), .A2(MEM_stage_inst_dmem_n12963), .ZN(MEM_stage_inst_dmem_n12894) );
NAND2_X1 MEM_stage_inst_dmem_U8718 ( .A1(MEM_stage_inst_dmem_n8590), .A2(MEM_stage_inst_dmem_n8589), .ZN(MEM_stage_inst_dmem_n12843) );
NAND2_X1 MEM_stage_inst_dmem_U8717 ( .A1(MEM_stage_inst_dmem_n8588), .A2(MEM_stage_inst_dmem_n14732), .ZN(MEM_stage_inst_dmem_n8589) );
NAND2_X1 MEM_stage_inst_dmem_U8716 ( .A1(MEM_stage_inst_dmem_ram_496), .A2(MEM_stage_inst_dmem_n8587), .ZN(MEM_stage_inst_dmem_n8590) );
NAND2_X1 MEM_stage_inst_dmem_U8715 ( .A1(MEM_stage_inst_dmem_n8586), .A2(MEM_stage_inst_dmem_n8585), .ZN(MEM_stage_inst_dmem_n12844) );
NAND2_X1 MEM_stage_inst_dmem_U8714 ( .A1(MEM_stage_inst_dmem_n8588), .A2(MEM_stage_inst_dmem_n109), .ZN(MEM_stage_inst_dmem_n8585) );
NAND2_X1 MEM_stage_inst_dmem_U8712 ( .A1(MEM_stage_inst_dmem_ram_497), .A2(MEM_stage_inst_dmem_n8587), .ZN(MEM_stage_inst_dmem_n8586) );
NAND2_X1 MEM_stage_inst_dmem_U8711 ( .A1(MEM_stage_inst_dmem_n8584), .A2(MEM_stage_inst_dmem_n8583), .ZN(MEM_stage_inst_dmem_n12845) );
NAND2_X1 MEM_stage_inst_dmem_U8710 ( .A1(MEM_stage_inst_dmem_n8588), .A2(MEM_stage_inst_dmem_n18887), .ZN(MEM_stage_inst_dmem_n8583) );
NAND2_X1 MEM_stage_inst_dmem_U8709 ( .A1(MEM_stage_inst_dmem_ram_498), .A2(MEM_stage_inst_dmem_n8587), .ZN(MEM_stage_inst_dmem_n8584) );
NAND2_X1 MEM_stage_inst_dmem_U8708 ( .A1(MEM_stage_inst_dmem_n8582), .A2(MEM_stage_inst_dmem_n8581), .ZN(MEM_stage_inst_dmem_n12846) );
NAND2_X1 MEM_stage_inst_dmem_U8707 ( .A1(MEM_stage_inst_dmem_n8588), .A2(MEM_stage_inst_dmem_n13064), .ZN(MEM_stage_inst_dmem_n8581) );
BUF_X1 MEM_stage_inst_dmem_U8706 ( .A(MEM_stage_inst_dmem_n21506), .Z(MEM_stage_inst_dmem_n13064) );
NAND2_X1 MEM_stage_inst_dmem_U8705 ( .A1(MEM_stage_inst_dmem_ram_499), .A2(MEM_stage_inst_dmem_n8587), .ZN(MEM_stage_inst_dmem_n8582) );
NAND2_X1 MEM_stage_inst_dmem_U8704 ( .A1(MEM_stage_inst_dmem_n8580), .A2(MEM_stage_inst_dmem_n8579), .ZN(MEM_stage_inst_dmem_n12847) );
NAND2_X1 MEM_stage_inst_dmem_U8703 ( .A1(MEM_stage_inst_dmem_n8588), .A2(EX_pipeline_reg_out_9), .ZN(MEM_stage_inst_dmem_n8579) );
NAND2_X1 MEM_stage_inst_dmem_U8702 ( .A1(MEM_stage_inst_dmem_ram_500), .A2(MEM_stage_inst_dmem_n8587), .ZN(MEM_stage_inst_dmem_n8580) );
NAND2_X1 MEM_stage_inst_dmem_U8701 ( .A1(MEM_stage_inst_dmem_n8578), .A2(MEM_stage_inst_dmem_n8577), .ZN(MEM_stage_inst_dmem_n12848) );
NAND2_X1 MEM_stage_inst_dmem_U8700 ( .A1(MEM_stage_inst_dmem_n8588), .A2(MEM_stage_inst_dmem_n13059), .ZN(MEM_stage_inst_dmem_n8577) );
BUF_X1 MEM_stage_inst_dmem_U8699 ( .A(MEM_stage_inst_dmem_n21508), .Z(MEM_stage_inst_dmem_n13059) );
NAND2_X1 MEM_stage_inst_dmem_U8698 ( .A1(MEM_stage_inst_dmem_ram_501), .A2(MEM_stage_inst_dmem_n8587), .ZN(MEM_stage_inst_dmem_n8578) );
NAND2_X1 MEM_stage_inst_dmem_U8697 ( .A1(MEM_stage_inst_dmem_n8576), .A2(MEM_stage_inst_dmem_n8575), .ZN(MEM_stage_inst_dmem_n12849) );
NAND2_X1 MEM_stage_inst_dmem_U8696 ( .A1(MEM_stage_inst_dmem_n8588), .A2(MEM_stage_inst_dmem_n13056), .ZN(MEM_stage_inst_dmem_n8575) );
BUF_X1 MEM_stage_inst_dmem_U8695 ( .A(MEM_stage_inst_dmem_n21340), .Z(MEM_stage_inst_dmem_n13056) );
NAND2_X1 MEM_stage_inst_dmem_U8694 ( .A1(MEM_stage_inst_dmem_ram_502), .A2(MEM_stage_inst_dmem_n8587), .ZN(MEM_stage_inst_dmem_n8576) );
NAND2_X1 MEM_stage_inst_dmem_U8693 ( .A1(MEM_stage_inst_dmem_n8574), .A2(MEM_stage_inst_dmem_n8573), .ZN(MEM_stage_inst_dmem_n12850) );
NAND2_X1 MEM_stage_inst_dmem_U8692 ( .A1(MEM_stage_inst_dmem_n8588), .A2(MEM_stage_inst_dmem_n101), .ZN(MEM_stage_inst_dmem_n8573) );
NAND2_X1 MEM_stage_inst_dmem_U8691 ( .A1(MEM_stage_inst_dmem_ram_503), .A2(MEM_stage_inst_dmem_n8587), .ZN(MEM_stage_inst_dmem_n8574) );
NAND2_X1 MEM_stage_inst_dmem_U8690 ( .A1(MEM_stage_inst_dmem_n8572), .A2(MEM_stage_inst_dmem_n8571), .ZN(MEM_stage_inst_dmem_n12851) );
NAND2_X1 MEM_stage_inst_dmem_U8689 ( .A1(MEM_stage_inst_dmem_n8588), .A2(MEM_stage_inst_dmem_n13051), .ZN(MEM_stage_inst_dmem_n8571) );
BUF_X1 MEM_stage_inst_dmem_U8688 ( .A(EX_pipeline_reg_out_13), .Z(MEM_stage_inst_dmem_n13051) );
NAND2_X1 MEM_stage_inst_dmem_U8687 ( .A1(MEM_stage_inst_dmem_ram_504), .A2(MEM_stage_inst_dmem_n8587), .ZN(MEM_stage_inst_dmem_n8572) );
NAND2_X1 MEM_stage_inst_dmem_U8686 ( .A1(MEM_stage_inst_dmem_n8570), .A2(MEM_stage_inst_dmem_n8569), .ZN(MEM_stage_inst_dmem_n12852) );
NAND2_X1 MEM_stage_inst_dmem_U8685 ( .A1(MEM_stage_inst_dmem_n8588), .A2(MEM_stage_inst_dmem_n20524), .ZN(MEM_stage_inst_dmem_n8569) );
NAND2_X1 MEM_stage_inst_dmem_U8684 ( .A1(MEM_stage_inst_dmem_ram_505), .A2(MEM_stage_inst_dmem_n8587), .ZN(MEM_stage_inst_dmem_n8570) );
NAND2_X1 MEM_stage_inst_dmem_U8683 ( .A1(MEM_stage_inst_dmem_n8568), .A2(MEM_stage_inst_dmem_n8567), .ZN(MEM_stage_inst_dmem_n12853) );
NAND2_X1 MEM_stage_inst_dmem_U8682 ( .A1(MEM_stage_inst_dmem_n8588), .A2(MEM_stage_inst_dmem_n18867), .ZN(MEM_stage_inst_dmem_n8567) );
NAND2_X1 MEM_stage_inst_dmem_U8681 ( .A1(MEM_stage_inst_dmem_ram_506), .A2(MEM_stage_inst_dmem_n8587), .ZN(MEM_stage_inst_dmem_n8568) );
NAND2_X1 MEM_stage_inst_dmem_U8680 ( .A1(MEM_stage_inst_dmem_n8566), .A2(MEM_stage_inst_dmem_n8565), .ZN(MEM_stage_inst_dmem_n12854) );
NAND2_X1 MEM_stage_inst_dmem_U8679 ( .A1(MEM_stage_inst_dmem_n8588), .A2(MEM_stage_inst_dmem_n13044), .ZN(MEM_stage_inst_dmem_n8565) );
BUF_X1 MEM_stage_inst_dmem_U8678 ( .A(EX_pipeline_reg_out_16), .Z(MEM_stage_inst_dmem_n13044) );
NAND2_X1 MEM_stage_inst_dmem_U8677 ( .A1(MEM_stage_inst_dmem_ram_507), .A2(MEM_stage_inst_dmem_n8587), .ZN(MEM_stage_inst_dmem_n8566) );
NAND2_X1 MEM_stage_inst_dmem_U8676 ( .A1(MEM_stage_inst_dmem_n8564), .A2(MEM_stage_inst_dmem_n8563), .ZN(MEM_stage_inst_dmem_n12855) );
NAND2_X1 MEM_stage_inst_dmem_U8675 ( .A1(MEM_stage_inst_dmem_n8588), .A2(MEM_stage_inst_dmem_n13041), .ZN(MEM_stage_inst_dmem_n8563) );
BUF_X1 MEM_stage_inst_dmem_U8674 ( .A(EX_pipeline_reg_out_17), .Z(MEM_stage_inst_dmem_n13041) );
NAND2_X1 MEM_stage_inst_dmem_U8673 ( .A1(MEM_stage_inst_dmem_ram_508), .A2(MEM_stage_inst_dmem_n8587), .ZN(MEM_stage_inst_dmem_n8564) );
NAND2_X1 MEM_stage_inst_dmem_U8672 ( .A1(MEM_stage_inst_dmem_n8562), .A2(MEM_stage_inst_dmem_n8561), .ZN(MEM_stage_inst_dmem_n12856) );
NAND2_X1 MEM_stage_inst_dmem_U8671 ( .A1(MEM_stage_inst_dmem_n8588), .A2(MEM_stage_inst_dmem_n116), .ZN(MEM_stage_inst_dmem_n8561) );
NAND2_X1 MEM_stage_inst_dmem_U8670 ( .A1(MEM_stage_inst_dmem_ram_509), .A2(MEM_stage_inst_dmem_n8587), .ZN(MEM_stage_inst_dmem_n8562) );
NAND2_X1 MEM_stage_inst_dmem_U8669 ( .A1(MEM_stage_inst_dmem_n8560), .A2(MEM_stage_inst_dmem_n8559), .ZN(MEM_stage_inst_dmem_n12857) );
NAND2_X1 MEM_stage_inst_dmem_U8668 ( .A1(MEM_stage_inst_dmem_n8588), .A2(MEM_stage_inst_dmem_n14696), .ZN(MEM_stage_inst_dmem_n8559) );
NAND2_X1 MEM_stage_inst_dmem_U8667 ( .A1(MEM_stage_inst_dmem_ram_510), .A2(MEM_stage_inst_dmem_n8587), .ZN(MEM_stage_inst_dmem_n8560) );
NAND2_X1 MEM_stage_inst_dmem_U8666 ( .A1(MEM_stage_inst_dmem_n8558), .A2(MEM_stage_inst_dmem_n8557), .ZN(MEM_stage_inst_dmem_n12858) );
NAND2_X1 MEM_stage_inst_dmem_U8665 ( .A1(MEM_stage_inst_dmem_n8588), .A2(MEM_stage_inst_dmem_n114), .ZN(MEM_stage_inst_dmem_n8557) );
INV_X1 MEM_stage_inst_dmem_U8664 ( .A(MEM_stage_inst_dmem_n8587), .ZN(MEM_stage_inst_dmem_n8588) );
NAND2_X1 MEM_stage_inst_dmem_U8663 ( .A1(MEM_stage_inst_dmem_ram_511), .A2(MEM_stage_inst_dmem_n8587), .ZN(MEM_stage_inst_dmem_n8558) );
NAND2_X1 MEM_stage_inst_dmem_U8662 ( .A1(MEM_stage_inst_dmem_n20934), .A2(MEM_stage_inst_dmem_n13182), .ZN(MEM_stage_inst_dmem_n8587) );
NOR2_X2 MEM_stage_inst_dmem_U8661 ( .A1(MEM_stage_inst_dmem_n17619), .A2(MEM_stage_inst_dmem_n15968), .ZN(MEM_stage_inst_dmem_n13182) );
NAND2_X1 MEM_stage_inst_dmem_U8660 ( .A1(EX_pipeline_reg_out_26), .A2(MEM_stage_inst_dmem_n13217), .ZN(MEM_stage_inst_dmem_n15968) );
NOR2_X1 MEM_stage_inst_dmem_U8659 ( .A1(n3522), .A2(MEM_stage_inst_dmem_n8556), .ZN(MEM_stage_inst_dmem_n13217) );
INV_X1 MEM_stage_inst_dmem_U8658 ( .A(EX_pipeline_reg_out_29), .ZN(MEM_stage_inst_dmem_n8556) );
NAND2_X1 MEM_stage_inst_dmem_U8657 ( .A1(EX_pipeline_reg_out_28), .A2(EX_pipeline_reg_out_27), .ZN(MEM_stage_inst_dmem_n17619) );
NOR2_X2 MEM_stage_inst_dmem_U8656 ( .A1(MEM_stage_inst_dmem_n12965), .A2(MEM_stage_inst_dmem_n12859), .ZN(MEM_stage_inst_dmem_n20934) );
NAND2_X1 MEM_stage_inst_dmem_U8655 ( .A1(EX_pipeline_reg_out_25), .A2(EX_pipeline_reg_out_22), .ZN(MEM_stage_inst_dmem_n12859) );
NAND2_X1 MEM_stage_inst_dmem_U8654 ( .A1(EX_pipeline_reg_out_24), .A2(EX_pipeline_reg_out_23), .ZN(MEM_stage_inst_dmem_n12965) );
NAND2_X1 MEM_stage_inst_dmem_U8653 ( .A1(MEM_stage_inst_dmem_n8555), .A2(MEM_stage_inst_dmem_n8554), .ZN(MEM_stage_inst_mem_read_data_15) );
NOR2_X1 MEM_stage_inst_dmem_U8652 ( .A1(MEM_stage_inst_dmem_n8553), .A2(MEM_stage_inst_dmem_n8552), .ZN(MEM_stage_inst_dmem_n8554) );
NOR2_X1 MEM_stage_inst_dmem_U8651 ( .A1(MEM_stage_inst_dmem_n8551), .A2(MEM_stage_inst_dmem_n8550), .ZN(MEM_stage_inst_dmem_n8552) );
NOR2_X1 MEM_stage_inst_dmem_U8650 ( .A1(MEM_stage_inst_dmem_n8549), .A2(MEM_stage_inst_dmem_n8548), .ZN(MEM_stage_inst_dmem_n8550) );
NAND2_X1 MEM_stage_inst_dmem_U8649 ( .A1(MEM_stage_inst_dmem_n8547), .A2(MEM_stage_inst_dmem_n8546), .ZN(MEM_stage_inst_dmem_n8548) );
NOR2_X1 MEM_stage_inst_dmem_U8648 ( .A1(MEM_stage_inst_dmem_n8545), .A2(MEM_stage_inst_dmem_n8544), .ZN(MEM_stage_inst_dmem_n8546) );
NAND2_X1 MEM_stage_inst_dmem_U8647 ( .A1(MEM_stage_inst_dmem_n8543), .A2(MEM_stage_inst_dmem_n8542), .ZN(MEM_stage_inst_dmem_n8544) );
NOR2_X1 MEM_stage_inst_dmem_U8646 ( .A1(MEM_stage_inst_dmem_n8541), .A2(MEM_stage_inst_dmem_n8540), .ZN(MEM_stage_inst_dmem_n8542) );
NAND2_X1 MEM_stage_inst_dmem_U8645 ( .A1(MEM_stage_inst_dmem_n8539), .A2(MEM_stage_inst_dmem_n8538), .ZN(MEM_stage_inst_dmem_n8540) );
NAND2_X1 MEM_stage_inst_dmem_U8644 ( .A1(MEM_stage_inst_dmem_n43), .A2(MEM_stage_inst_dmem_ram_447), .ZN(MEM_stage_inst_dmem_n8538) );
NAND2_X1 MEM_stage_inst_dmem_U8643 ( .A1(MEM_stage_inst_dmem_n40), .A2(MEM_stage_inst_dmem_ram_95), .ZN(MEM_stage_inst_dmem_n8539) );
NAND2_X1 MEM_stage_inst_dmem_U8642 ( .A1(MEM_stage_inst_dmem_n8537), .A2(MEM_stage_inst_dmem_n8536), .ZN(MEM_stage_inst_dmem_n8541) );
NAND2_X1 MEM_stage_inst_dmem_U8641 ( .A1(MEM_stage_inst_dmem_ram_511), .A2(MEM_stage_inst_dmem_n8535), .ZN(MEM_stage_inst_dmem_n8536) );
NAND2_X1 MEM_stage_inst_dmem_U8640 ( .A1(MEM_stage_inst_dmem_ram_239), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n8537) );
NOR2_X1 MEM_stage_inst_dmem_U8639 ( .A1(MEM_stage_inst_dmem_n8534), .A2(MEM_stage_inst_dmem_n8533), .ZN(MEM_stage_inst_dmem_n8543) );
NAND2_X1 MEM_stage_inst_dmem_U8638 ( .A1(MEM_stage_inst_dmem_n8532), .A2(MEM_stage_inst_dmem_n8531), .ZN(MEM_stage_inst_dmem_n8533) );
NAND2_X1 MEM_stage_inst_dmem_U8637 ( .A1(MEM_stage_inst_dmem_ram_495), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n8531) );
NAND2_X1 MEM_stage_inst_dmem_U8636 ( .A1(MEM_stage_inst_dmem_ram_463), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n8532) );
NAND2_X1 MEM_stage_inst_dmem_U8635 ( .A1(MEM_stage_inst_dmem_n8530), .A2(MEM_stage_inst_dmem_n8529), .ZN(MEM_stage_inst_dmem_n8534) );
NAND2_X1 MEM_stage_inst_dmem_U8634 ( .A1(MEM_stage_inst_dmem_ram_911), .A2(MEM_stage_inst_dmem_n72), .ZN(MEM_stage_inst_dmem_n8529) );
NAND2_X1 MEM_stage_inst_dmem_U8633 ( .A1(MEM_stage_inst_dmem_ram_159), .A2(MEM_stage_inst_dmem_n44), .ZN(MEM_stage_inst_dmem_n8530) );
NAND2_X1 MEM_stage_inst_dmem_U8632 ( .A1(MEM_stage_inst_dmem_n8528), .A2(MEM_stage_inst_dmem_n8527), .ZN(MEM_stage_inst_dmem_n8545) );
NOR2_X1 MEM_stage_inst_dmem_U8631 ( .A1(MEM_stage_inst_dmem_n8526), .A2(MEM_stage_inst_dmem_n8525), .ZN(MEM_stage_inst_dmem_n8527) );
NAND2_X1 MEM_stage_inst_dmem_U8630 ( .A1(MEM_stage_inst_dmem_n8524), .A2(MEM_stage_inst_dmem_n8523), .ZN(MEM_stage_inst_dmem_n8525) );
NAND2_X1 MEM_stage_inst_dmem_U8629 ( .A1(MEM_stage_inst_dmem_ram_479), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n8523) );
NAND2_X1 MEM_stage_inst_dmem_U8628 ( .A1(MEM_stage_inst_dmem_ram_111), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n8524) );
NAND2_X1 MEM_stage_inst_dmem_U8627 ( .A1(MEM_stage_inst_dmem_n8522), .A2(MEM_stage_inst_dmem_n8521), .ZN(MEM_stage_inst_dmem_n8526) );
NAND2_X1 MEM_stage_inst_dmem_U8626 ( .A1(MEM_stage_inst_dmem_ram_255), .A2(MEM_stage_inst_dmem_n39), .ZN(MEM_stage_inst_dmem_n8521) );
NAND2_X1 MEM_stage_inst_dmem_U8625 ( .A1(MEM_stage_inst_dmem_ram_671), .A2(MEM_stage_inst_dmem_n3076), .ZN(MEM_stage_inst_dmem_n8522) );
NOR2_X1 MEM_stage_inst_dmem_U8624 ( .A1(MEM_stage_inst_dmem_n8520), .A2(MEM_stage_inst_dmem_n8519), .ZN(MEM_stage_inst_dmem_n8528) );
NAND2_X1 MEM_stage_inst_dmem_U8623 ( .A1(MEM_stage_inst_dmem_n8518), .A2(MEM_stage_inst_dmem_n8517), .ZN(MEM_stage_inst_dmem_n8519) );
NAND2_X1 MEM_stage_inst_dmem_U8622 ( .A1(MEM_stage_inst_dmem_ram_223), .A2(MEM_stage_inst_dmem_n51), .ZN(MEM_stage_inst_dmem_n8517) );
NAND2_X1 MEM_stage_inst_dmem_U8621 ( .A1(MEM_stage_inst_dmem_ram_271), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n8518) );
NAND2_X1 MEM_stage_inst_dmem_U8620 ( .A1(MEM_stage_inst_dmem_n8516), .A2(MEM_stage_inst_dmem_n8515), .ZN(MEM_stage_inst_dmem_n8520) );
NAND2_X1 MEM_stage_inst_dmem_U8619 ( .A1(MEM_stage_inst_dmem_ram_655), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n8515) );
NAND2_X1 MEM_stage_inst_dmem_U8618 ( .A1(MEM_stage_inst_dmem_ram_927), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n8516) );
NOR2_X1 MEM_stage_inst_dmem_U8617 ( .A1(MEM_stage_inst_dmem_n8514), .A2(MEM_stage_inst_dmem_n8513), .ZN(MEM_stage_inst_dmem_n8547) );
NAND2_X1 MEM_stage_inst_dmem_U8616 ( .A1(MEM_stage_inst_dmem_n8512), .A2(MEM_stage_inst_dmem_n8511), .ZN(MEM_stage_inst_dmem_n8513) );
NOR2_X1 MEM_stage_inst_dmem_U8615 ( .A1(MEM_stage_inst_dmem_n8510), .A2(MEM_stage_inst_dmem_n8509), .ZN(MEM_stage_inst_dmem_n8511) );
NAND2_X1 MEM_stage_inst_dmem_U8614 ( .A1(MEM_stage_inst_dmem_n8508), .A2(MEM_stage_inst_dmem_n8507), .ZN(MEM_stage_inst_dmem_n8509) );
NAND2_X1 MEM_stage_inst_dmem_U8613 ( .A1(MEM_stage_inst_dmem_ram_63), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n8507) );
NAND2_X1 MEM_stage_inst_dmem_U8612 ( .A1(MEM_stage_inst_dmem_ram_559), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n8508) );
NAND2_X1 MEM_stage_inst_dmem_U8611 ( .A1(MEM_stage_inst_dmem_n8506), .A2(MEM_stage_inst_dmem_n8505), .ZN(MEM_stage_inst_dmem_n8510) );
NAND2_X1 MEM_stage_inst_dmem_U8610 ( .A1(MEM_stage_inst_dmem_ram_335), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n8505) );
NAND2_X1 MEM_stage_inst_dmem_U8609 ( .A1(MEM_stage_inst_dmem_ram_607), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n8506) );
NOR2_X1 MEM_stage_inst_dmem_U8608 ( .A1(MEM_stage_inst_dmem_n8504), .A2(MEM_stage_inst_dmem_n8503), .ZN(MEM_stage_inst_dmem_n8512) );
NAND2_X1 MEM_stage_inst_dmem_U8607 ( .A1(MEM_stage_inst_dmem_n8502), .A2(MEM_stage_inst_dmem_n8501), .ZN(MEM_stage_inst_dmem_n8503) );
NAND2_X1 MEM_stage_inst_dmem_U8606 ( .A1(MEM_stage_inst_dmem_ram_319), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n8501) );
NAND2_X1 MEM_stage_inst_dmem_U8605 ( .A1(MEM_stage_inst_dmem_ram_31), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n8502) );
NAND2_X1 MEM_stage_inst_dmem_U8604 ( .A1(MEM_stage_inst_dmem_n8500), .A2(MEM_stage_inst_dmem_n8499), .ZN(MEM_stage_inst_dmem_n8504) );
NAND2_X1 MEM_stage_inst_dmem_U8603 ( .A1(MEM_stage_inst_dmem_ram_127), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n8499) );
NAND2_X1 MEM_stage_inst_dmem_U8602 ( .A1(MEM_stage_inst_dmem_ram_527), .A2(MEM_stage_inst_dmem_n71), .ZN(MEM_stage_inst_dmem_n8500) );
NAND2_X1 MEM_stage_inst_dmem_U8601 ( .A1(MEM_stage_inst_dmem_n8498), .A2(MEM_stage_inst_dmem_n8497), .ZN(MEM_stage_inst_dmem_n8514) );
NOR2_X1 MEM_stage_inst_dmem_U8600 ( .A1(MEM_stage_inst_dmem_n8496), .A2(MEM_stage_inst_dmem_n8495), .ZN(MEM_stage_inst_dmem_n8497) );
NAND2_X1 MEM_stage_inst_dmem_U8599 ( .A1(MEM_stage_inst_dmem_n8494), .A2(MEM_stage_inst_dmem_n8493), .ZN(MEM_stage_inst_dmem_n8495) );
NAND2_X1 MEM_stage_inst_dmem_U8598 ( .A1(MEM_stage_inst_dmem_ram_895), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n8493) );
NAND2_X1 MEM_stage_inst_dmem_U8597 ( .A1(MEM_stage_inst_dmem_ram_399), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n8494) );
NAND2_X1 MEM_stage_inst_dmem_U8596 ( .A1(MEM_stage_inst_dmem_n8492), .A2(MEM_stage_inst_dmem_n8491), .ZN(MEM_stage_inst_dmem_n8496) );
NAND2_X1 MEM_stage_inst_dmem_U8595 ( .A1(MEM_stage_inst_dmem_ram_575), .A2(MEM_stage_inst_dmem_n41), .ZN(MEM_stage_inst_dmem_n8491) );
NAND2_X1 MEM_stage_inst_dmem_U8594 ( .A1(MEM_stage_inst_dmem_ram_623), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n8492) );
NOR2_X1 MEM_stage_inst_dmem_U8593 ( .A1(MEM_stage_inst_dmem_n8490), .A2(MEM_stage_inst_dmem_n8489), .ZN(MEM_stage_inst_dmem_n8498) );
NAND2_X1 MEM_stage_inst_dmem_U8592 ( .A1(MEM_stage_inst_dmem_n8488), .A2(MEM_stage_inst_dmem_n8487), .ZN(MEM_stage_inst_dmem_n8489) );
NAND2_X1 MEM_stage_inst_dmem_U8591 ( .A1(MEM_stage_inst_dmem_ram_815), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n8487) );
NAND2_X1 MEM_stage_inst_dmem_U8590 ( .A1(MEM_stage_inst_dmem_ram_735), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n8488) );
NAND2_X1 MEM_stage_inst_dmem_U8589 ( .A1(MEM_stage_inst_dmem_n8486), .A2(MEM_stage_inst_dmem_n8485), .ZN(MEM_stage_inst_dmem_n8490) );
NAND2_X1 MEM_stage_inst_dmem_U8588 ( .A1(MEM_stage_inst_dmem_n46), .A2(MEM_stage_inst_dmem_ram_831), .ZN(MEM_stage_inst_dmem_n8485) );
NAND2_X1 MEM_stage_inst_dmem_U8587 ( .A1(MEM_stage_inst_dmem_n22), .A2(MEM_stage_inst_dmem_ram_751), .ZN(MEM_stage_inst_dmem_n8486) );
NAND2_X1 MEM_stage_inst_dmem_U8586 ( .A1(MEM_stage_inst_dmem_n8484), .A2(MEM_stage_inst_dmem_n8483), .ZN(MEM_stage_inst_dmem_n8549) );
NOR2_X1 MEM_stage_inst_dmem_U8585 ( .A1(MEM_stage_inst_dmem_n8482), .A2(MEM_stage_inst_dmem_n8481), .ZN(MEM_stage_inst_dmem_n8483) );
NAND2_X1 MEM_stage_inst_dmem_U8584 ( .A1(MEM_stage_inst_dmem_n8480), .A2(MEM_stage_inst_dmem_n8479), .ZN(MEM_stage_inst_dmem_n8481) );
NOR2_X1 MEM_stage_inst_dmem_U8583 ( .A1(MEM_stage_inst_dmem_n8478), .A2(MEM_stage_inst_dmem_n8477), .ZN(MEM_stage_inst_dmem_n8479) );
NAND2_X1 MEM_stage_inst_dmem_U8582 ( .A1(MEM_stage_inst_dmem_n8476), .A2(MEM_stage_inst_dmem_n8475), .ZN(MEM_stage_inst_dmem_n8477) );
NAND2_X1 MEM_stage_inst_dmem_U8581 ( .A1(MEM_stage_inst_dmem_ram_959), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n8475) );
NAND2_X1 MEM_stage_inst_dmem_U8580 ( .A1(MEM_stage_inst_dmem_ram_543), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n8476) );
NAND2_X1 MEM_stage_inst_dmem_U8579 ( .A1(MEM_stage_inst_dmem_n8474), .A2(MEM_stage_inst_dmem_n8473), .ZN(MEM_stage_inst_dmem_n8478) );
NAND2_X1 MEM_stage_inst_dmem_U8578 ( .A1(MEM_stage_inst_dmem_ram_783), .A2(MEM_stage_inst_dmem_n8472), .ZN(MEM_stage_inst_dmem_n8473) );
NAND2_X1 MEM_stage_inst_dmem_U8577 ( .A1(MEM_stage_inst_dmem_ram_767), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n8474) );
NOR2_X1 MEM_stage_inst_dmem_U8576 ( .A1(MEM_stage_inst_dmem_n8471), .A2(MEM_stage_inst_dmem_n8470), .ZN(MEM_stage_inst_dmem_n8480) );
NAND2_X1 MEM_stage_inst_dmem_U8575 ( .A1(MEM_stage_inst_dmem_n8469), .A2(MEM_stage_inst_dmem_n8468), .ZN(MEM_stage_inst_dmem_n8470) );
NAND2_X1 MEM_stage_inst_dmem_U8574 ( .A1(MEM_stage_inst_dmem_ram_47), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n8468) );
NAND2_X1 MEM_stage_inst_dmem_U8573 ( .A1(MEM_stage_inst_dmem_ram_943), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n8469) );
NAND2_X1 MEM_stage_inst_dmem_U8572 ( .A1(MEM_stage_inst_dmem_n8467), .A2(MEM_stage_inst_dmem_n8466), .ZN(MEM_stage_inst_dmem_n8471) );
NAND2_X1 MEM_stage_inst_dmem_U8571 ( .A1(MEM_stage_inst_dmem_ram_975), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n8466) );
NAND2_X1 MEM_stage_inst_dmem_U8570 ( .A1(MEM_stage_inst_dmem_ram_143), .A2(MEM_stage_inst_dmem_n61), .ZN(MEM_stage_inst_dmem_n8467) );
NAND2_X1 MEM_stage_inst_dmem_U8569 ( .A1(MEM_stage_inst_dmem_n8465), .A2(MEM_stage_inst_dmem_n8464), .ZN(MEM_stage_inst_dmem_n8482) );
NOR2_X1 MEM_stage_inst_dmem_U8568 ( .A1(MEM_stage_inst_dmem_n8463), .A2(MEM_stage_inst_dmem_n8462), .ZN(MEM_stage_inst_dmem_n8464) );
NAND2_X1 MEM_stage_inst_dmem_U8567 ( .A1(MEM_stage_inst_dmem_n8461), .A2(MEM_stage_inst_dmem_n8460), .ZN(MEM_stage_inst_dmem_n8462) );
NAND2_X1 MEM_stage_inst_dmem_U8566 ( .A1(MEM_stage_inst_dmem_ram_847), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n8460) );
NAND2_X1 MEM_stage_inst_dmem_U8565 ( .A1(MEM_stage_inst_dmem_ram_287), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n8461) );
NAND2_X1 MEM_stage_inst_dmem_U8564 ( .A1(MEM_stage_inst_dmem_n8459), .A2(MEM_stage_inst_dmem_n8458), .ZN(MEM_stage_inst_dmem_n8463) );
NAND2_X1 MEM_stage_inst_dmem_U8563 ( .A1(MEM_stage_inst_dmem_ram_303), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n8458) );
NAND2_X1 MEM_stage_inst_dmem_U8562 ( .A1(MEM_stage_inst_dmem_ram_799), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n8459) );
NOR2_X1 MEM_stage_inst_dmem_U8561 ( .A1(MEM_stage_inst_dmem_n8457), .A2(MEM_stage_inst_dmem_n8456), .ZN(MEM_stage_inst_dmem_n8465) );
NAND2_X1 MEM_stage_inst_dmem_U8560 ( .A1(MEM_stage_inst_dmem_n8455), .A2(MEM_stage_inst_dmem_n8454), .ZN(MEM_stage_inst_dmem_n8456) );
NAND2_X1 MEM_stage_inst_dmem_U8559 ( .A1(MEM_stage_inst_dmem_ram_367), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n8454) );
NAND2_X1 MEM_stage_inst_dmem_U8558 ( .A1(MEM_stage_inst_dmem_ram_687), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n8455) );
NAND2_X1 MEM_stage_inst_dmem_U8557 ( .A1(MEM_stage_inst_dmem_n8453), .A2(MEM_stage_inst_dmem_n8452), .ZN(MEM_stage_inst_dmem_n8457) );
NAND2_X1 MEM_stage_inst_dmem_U8556 ( .A1(MEM_stage_inst_dmem_ram_207), .A2(MEM_stage_inst_dmem_n36), .ZN(MEM_stage_inst_dmem_n8452) );
NAND2_X1 MEM_stage_inst_dmem_U8555 ( .A1(MEM_stage_inst_dmem_ram_351), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n8453) );
NOR2_X1 MEM_stage_inst_dmem_U8554 ( .A1(MEM_stage_inst_dmem_n8450), .A2(MEM_stage_inst_dmem_n8449), .ZN(MEM_stage_inst_dmem_n8484) );
NAND2_X1 MEM_stage_inst_dmem_U8553 ( .A1(MEM_stage_inst_dmem_n8448), .A2(MEM_stage_inst_dmem_n8447), .ZN(MEM_stage_inst_dmem_n8449) );
NOR2_X1 MEM_stage_inst_dmem_U8552 ( .A1(MEM_stage_inst_dmem_n8446), .A2(MEM_stage_inst_dmem_n8445), .ZN(MEM_stage_inst_dmem_n8447) );
NAND2_X1 MEM_stage_inst_dmem_U8551 ( .A1(MEM_stage_inst_dmem_n8444), .A2(MEM_stage_inst_dmem_n8443), .ZN(MEM_stage_inst_dmem_n8445) );
NAND2_X1 MEM_stage_inst_dmem_U8550 ( .A1(MEM_stage_inst_dmem_ram_879), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n8443) );
NAND2_X1 MEM_stage_inst_dmem_U8549 ( .A1(MEM_stage_inst_dmem_ram_991), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n8444) );
NAND2_X1 MEM_stage_inst_dmem_U8548 ( .A1(MEM_stage_inst_dmem_n8442), .A2(MEM_stage_inst_dmem_n8441), .ZN(MEM_stage_inst_dmem_n8446) );
NAND2_X1 MEM_stage_inst_dmem_U8547 ( .A1(MEM_stage_inst_dmem_ram_415), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n8441) );
NAND2_X1 MEM_stage_inst_dmem_U8546 ( .A1(MEM_stage_inst_dmem_ram_79), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n8442) );
NOR2_X1 MEM_stage_inst_dmem_U8545 ( .A1(MEM_stage_inst_dmem_n8440), .A2(MEM_stage_inst_dmem_n8439), .ZN(MEM_stage_inst_dmem_n8448) );
NAND2_X1 MEM_stage_inst_dmem_U8544 ( .A1(MEM_stage_inst_dmem_n8438), .A2(MEM_stage_inst_dmem_n8437), .ZN(MEM_stage_inst_dmem_n8439) );
NAND2_X1 MEM_stage_inst_dmem_U8543 ( .A1(MEM_stage_inst_dmem_ram_703), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n8437) );
NAND2_X1 MEM_stage_inst_dmem_U8542 ( .A1(MEM_stage_inst_dmem_ram_175), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n8438) );
NAND2_X1 MEM_stage_inst_dmem_U8541 ( .A1(MEM_stage_inst_dmem_n8436), .A2(MEM_stage_inst_dmem_n8435), .ZN(MEM_stage_inst_dmem_n8440) );
NAND2_X1 MEM_stage_inst_dmem_U8540 ( .A1(MEM_stage_inst_dmem_n27), .A2(MEM_stage_inst_dmem_ram_591), .ZN(MEM_stage_inst_dmem_n8435) );
NAND2_X1 MEM_stage_inst_dmem_U8539 ( .A1(MEM_stage_inst_dmem_n8434), .A2(MEM_stage_inst_dmem_ram_191), .ZN(MEM_stage_inst_dmem_n8436) );
NAND2_X1 MEM_stage_inst_dmem_U8538 ( .A1(MEM_stage_inst_dmem_n8433), .A2(MEM_stage_inst_dmem_n8432), .ZN(MEM_stage_inst_dmem_n8450) );
NOR2_X1 MEM_stage_inst_dmem_U8537 ( .A1(MEM_stage_inst_dmem_n8431), .A2(MEM_stage_inst_dmem_n8430), .ZN(MEM_stage_inst_dmem_n8432) );
NAND2_X1 MEM_stage_inst_dmem_U8536 ( .A1(MEM_stage_inst_dmem_n8429), .A2(MEM_stage_inst_dmem_n8428), .ZN(MEM_stage_inst_dmem_n8430) );
NAND2_X1 MEM_stage_inst_dmem_U8535 ( .A1(MEM_stage_inst_dmem_ram_719), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n8428) );
NAND2_X1 MEM_stage_inst_dmem_U8534 ( .A1(MEM_stage_inst_dmem_ram_1023), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n8429) );
NAND2_X1 MEM_stage_inst_dmem_U8533 ( .A1(MEM_stage_inst_dmem_n8427), .A2(MEM_stage_inst_dmem_n8426), .ZN(MEM_stage_inst_dmem_n8431) );
NAND2_X1 MEM_stage_inst_dmem_U8532 ( .A1(MEM_stage_inst_dmem_ram_863), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n8426) );
NAND2_X1 MEM_stage_inst_dmem_U8531 ( .A1(MEM_stage_inst_dmem_ram_1007), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n8427) );
NOR2_X1 MEM_stage_inst_dmem_U8530 ( .A1(MEM_stage_inst_dmem_n8425), .A2(MEM_stage_inst_dmem_n8424), .ZN(MEM_stage_inst_dmem_n8433) );
NAND2_X1 MEM_stage_inst_dmem_U8529 ( .A1(MEM_stage_inst_dmem_n8423), .A2(MEM_stage_inst_dmem_n8422), .ZN(MEM_stage_inst_dmem_n8424) );
NAND2_X1 MEM_stage_inst_dmem_U8528 ( .A1(MEM_stage_inst_dmem_n8421), .A2(MEM_stage_inst_dmem_ram_431), .ZN(MEM_stage_inst_dmem_n8422) );
NAND2_X1 MEM_stage_inst_dmem_U8527 ( .A1(MEM_stage_inst_dmem_n77), .A2(MEM_stage_inst_dmem_ram_15), .ZN(MEM_stage_inst_dmem_n8423) );
NAND2_X1 MEM_stage_inst_dmem_U8526 ( .A1(MEM_stage_inst_dmem_n8420), .A2(MEM_stage_inst_dmem_n8419), .ZN(MEM_stage_inst_dmem_n8425) );
NAND2_X1 MEM_stage_inst_dmem_U8525 ( .A1(MEM_stage_inst_dmem_n32), .A2(MEM_stage_inst_dmem_ram_639), .ZN(MEM_stage_inst_dmem_n8419) );
NAND2_X1 MEM_stage_inst_dmem_U8524 ( .A1(MEM_stage_inst_dmem_n33), .A2(MEM_stage_inst_dmem_ram_383), .ZN(MEM_stage_inst_dmem_n8420) );
NOR2_X1 MEM_stage_inst_dmem_U8523 ( .A1(MEM_stage_inst_dmem_n8418), .A2(MEM_stage_inst_dmem_n8417), .ZN(MEM_stage_inst_dmem_n8553) );
NOR2_X1 MEM_stage_inst_dmem_U8522 ( .A1(MEM_stage_inst_dmem_n8416), .A2(MEM_stage_inst_dmem_n8415), .ZN(MEM_stage_inst_dmem_n8418) );
NAND2_X1 MEM_stage_inst_dmem_U8521 ( .A1(MEM_stage_inst_dmem_n8414), .A2(MEM_stage_inst_dmem_n8413), .ZN(MEM_stage_inst_dmem_n8415) );
NOR2_X1 MEM_stage_inst_dmem_U8520 ( .A1(MEM_stage_inst_dmem_n8412), .A2(MEM_stage_inst_dmem_n8411), .ZN(MEM_stage_inst_dmem_n8413) );
NAND2_X1 MEM_stage_inst_dmem_U8519 ( .A1(MEM_stage_inst_dmem_n8410), .A2(MEM_stage_inst_dmem_n8409), .ZN(MEM_stage_inst_dmem_n8411) );
NOR2_X1 MEM_stage_inst_dmem_U8518 ( .A1(MEM_stage_inst_dmem_n8408), .A2(MEM_stage_inst_dmem_n8407), .ZN(MEM_stage_inst_dmem_n8409) );
NAND2_X1 MEM_stage_inst_dmem_U8517 ( .A1(MEM_stage_inst_dmem_n8406), .A2(MEM_stage_inst_dmem_n8405), .ZN(MEM_stage_inst_dmem_n8407) );
NAND2_X1 MEM_stage_inst_dmem_U8516 ( .A1(MEM_stage_inst_dmem_ram_3727), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n8405) );
NAND2_X1 MEM_stage_inst_dmem_U8515 ( .A1(MEM_stage_inst_dmem_ram_3999), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n8406) );
NAND2_X1 MEM_stage_inst_dmem_U8514 ( .A1(MEM_stage_inst_dmem_n8404), .A2(MEM_stage_inst_dmem_n8403), .ZN(MEM_stage_inst_dmem_n8408) );
NAND2_X1 MEM_stage_inst_dmem_U8513 ( .A1(MEM_stage_inst_dmem_ram_4047), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n8403) );
NAND2_X1 MEM_stage_inst_dmem_U8512 ( .A1(MEM_stage_inst_dmem_ram_3839), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n8404) );
NOR2_X1 MEM_stage_inst_dmem_U8511 ( .A1(MEM_stage_inst_dmem_n8402), .A2(MEM_stage_inst_dmem_n8401), .ZN(MEM_stage_inst_dmem_n8410) );
NAND2_X1 MEM_stage_inst_dmem_U8510 ( .A1(MEM_stage_inst_dmem_n8400), .A2(MEM_stage_inst_dmem_n8399), .ZN(MEM_stage_inst_dmem_n8401) );
NAND2_X1 MEM_stage_inst_dmem_U8509 ( .A1(MEM_stage_inst_dmem_ram_3791), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n8399) );
NAND2_X1 MEM_stage_inst_dmem_U8508 ( .A1(MEM_stage_inst_dmem_ram_4031), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n8400) );
NAND2_X1 MEM_stage_inst_dmem_U8507 ( .A1(MEM_stage_inst_dmem_n8398), .A2(MEM_stage_inst_dmem_n8397), .ZN(MEM_stage_inst_dmem_n8402) );
NAND2_X1 MEM_stage_inst_dmem_U8506 ( .A1(MEM_stage_inst_dmem_ram_3151), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n8397) );
NAND2_X1 MEM_stage_inst_dmem_U8505 ( .A1(MEM_stage_inst_dmem_ram_4079), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n8398) );
NAND2_X1 MEM_stage_inst_dmem_U8504 ( .A1(MEM_stage_inst_dmem_n8396), .A2(MEM_stage_inst_dmem_n8395), .ZN(MEM_stage_inst_dmem_n8412) );
NOR2_X1 MEM_stage_inst_dmem_U8503 ( .A1(MEM_stage_inst_dmem_n8394), .A2(MEM_stage_inst_dmem_n8393), .ZN(MEM_stage_inst_dmem_n8395) );
NAND2_X1 MEM_stage_inst_dmem_U8502 ( .A1(MEM_stage_inst_dmem_n8392), .A2(MEM_stage_inst_dmem_n8391), .ZN(MEM_stage_inst_dmem_n8393) );
NAND2_X1 MEM_stage_inst_dmem_U8501 ( .A1(MEM_stage_inst_dmem_ram_3631), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n8391) );
NAND2_X1 MEM_stage_inst_dmem_U8500 ( .A1(MEM_stage_inst_dmem_ram_4063), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n8392) );
NAND2_X1 MEM_stage_inst_dmem_U8499 ( .A1(MEM_stage_inst_dmem_n8390), .A2(MEM_stage_inst_dmem_n8389), .ZN(MEM_stage_inst_dmem_n8394) );
NAND2_X1 MEM_stage_inst_dmem_U8498 ( .A1(MEM_stage_inst_dmem_ram_3119), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n8389) );
NAND2_X1 MEM_stage_inst_dmem_U8497 ( .A1(MEM_stage_inst_dmem_ram_3359), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n8390) );
NOR2_X1 MEM_stage_inst_dmem_U8496 ( .A1(MEM_stage_inst_dmem_n8388), .A2(MEM_stage_inst_dmem_n8387), .ZN(MEM_stage_inst_dmem_n8396) );
NAND2_X1 MEM_stage_inst_dmem_U8495 ( .A1(MEM_stage_inst_dmem_n8386), .A2(MEM_stage_inst_dmem_n8385), .ZN(MEM_stage_inst_dmem_n8387) );
NAND2_X1 MEM_stage_inst_dmem_U8494 ( .A1(MEM_stage_inst_dmem_ram_3503), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n8385) );
NAND2_X1 MEM_stage_inst_dmem_U8493 ( .A1(MEM_stage_inst_dmem_ram_3215), .A2(MEM_stage_inst_dmem_n61), .ZN(MEM_stage_inst_dmem_n8386) );
NAND2_X1 MEM_stage_inst_dmem_U8492 ( .A1(MEM_stage_inst_dmem_n8384), .A2(MEM_stage_inst_dmem_n8383), .ZN(MEM_stage_inst_dmem_n8388) );
NAND2_X1 MEM_stage_inst_dmem_U8491 ( .A1(MEM_stage_inst_dmem_ram_3983), .A2(MEM_stage_inst_dmem_n72), .ZN(MEM_stage_inst_dmem_n8383) );
NAND2_X1 MEM_stage_inst_dmem_U8490 ( .A1(MEM_stage_inst_dmem_ram_3327), .A2(MEM_stage_inst_dmem_n39), .ZN(MEM_stage_inst_dmem_n8384) );
NOR2_X1 MEM_stage_inst_dmem_U8489 ( .A1(MEM_stage_inst_dmem_n8382), .A2(MEM_stage_inst_dmem_n8381), .ZN(MEM_stage_inst_dmem_n8414) );
NAND2_X1 MEM_stage_inst_dmem_U8488 ( .A1(MEM_stage_inst_dmem_n8380), .A2(MEM_stage_inst_dmem_n8379), .ZN(MEM_stage_inst_dmem_n8381) );
NOR2_X1 MEM_stage_inst_dmem_U8487 ( .A1(MEM_stage_inst_dmem_n8378), .A2(MEM_stage_inst_dmem_n8377), .ZN(MEM_stage_inst_dmem_n8379) );
NAND2_X1 MEM_stage_inst_dmem_U8486 ( .A1(MEM_stage_inst_dmem_n8376), .A2(MEM_stage_inst_dmem_n8375), .ZN(MEM_stage_inst_dmem_n8377) );
NAND2_X1 MEM_stage_inst_dmem_U8485 ( .A1(MEM_stage_inst_dmem_ram_3583), .A2(MEM_stage_inst_dmem_n64), .ZN(MEM_stage_inst_dmem_n8375) );
NAND2_X1 MEM_stage_inst_dmem_U8484 ( .A1(MEM_stage_inst_dmem_ram_3519), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n8376) );
NAND2_X1 MEM_stage_inst_dmem_U8483 ( .A1(MEM_stage_inst_dmem_n8374), .A2(MEM_stage_inst_dmem_n8373), .ZN(MEM_stage_inst_dmem_n8378) );
NAND2_X1 MEM_stage_inst_dmem_U8482 ( .A1(MEM_stage_inst_dmem_ram_3407), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n8373) );
NAND2_X1 MEM_stage_inst_dmem_U8481 ( .A1(MEM_stage_inst_dmem_ram_3935), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n8374) );
NOR2_X1 MEM_stage_inst_dmem_U8480 ( .A1(MEM_stage_inst_dmem_n8371), .A2(MEM_stage_inst_dmem_n8370), .ZN(MEM_stage_inst_dmem_n8380) );
NAND2_X1 MEM_stage_inst_dmem_U8479 ( .A1(MEM_stage_inst_dmem_n8369), .A2(MEM_stage_inst_dmem_n8368), .ZN(MEM_stage_inst_dmem_n8370) );
NAND2_X1 MEM_stage_inst_dmem_U8478 ( .A1(MEM_stage_inst_dmem_ram_3967), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n8368) );
NAND2_X1 MEM_stage_inst_dmem_U8477 ( .A1(MEM_stage_inst_dmem_ram_3279), .A2(MEM_stage_inst_dmem_n36), .ZN(MEM_stage_inst_dmem_n8369) );
NAND2_X1 MEM_stage_inst_dmem_U8476 ( .A1(MEM_stage_inst_dmem_n8367), .A2(MEM_stage_inst_dmem_n8366), .ZN(MEM_stage_inst_dmem_n8371) );
NAND2_X1 MEM_stage_inst_dmem_U8475 ( .A1(MEM_stage_inst_dmem_n8472), .A2(MEM_stage_inst_dmem_ram_3855), .ZN(MEM_stage_inst_dmem_n8366) );
NAND2_X1 MEM_stage_inst_dmem_U8474 ( .A1(MEM_stage_inst_dmem_n63), .A2(MEM_stage_inst_dmem_ram_3951), .ZN(MEM_stage_inst_dmem_n8367) );
NAND2_X1 MEM_stage_inst_dmem_U8473 ( .A1(MEM_stage_inst_dmem_n8365), .A2(MEM_stage_inst_dmem_n8364), .ZN(MEM_stage_inst_dmem_n8382) );
NOR2_X1 MEM_stage_inst_dmem_U8472 ( .A1(MEM_stage_inst_dmem_n8363), .A2(MEM_stage_inst_dmem_n8362), .ZN(MEM_stage_inst_dmem_n8364) );
NAND2_X1 MEM_stage_inst_dmem_U8471 ( .A1(MEM_stage_inst_dmem_n8361), .A2(MEM_stage_inst_dmem_n8360), .ZN(MEM_stage_inst_dmem_n8362) );
NAND2_X1 MEM_stage_inst_dmem_U8470 ( .A1(MEM_stage_inst_dmem_ram_3391), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n8360) );
NAND2_X1 MEM_stage_inst_dmem_U8469 ( .A1(MEM_stage_inst_dmem_ram_3135), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n8361) );
NAND2_X1 MEM_stage_inst_dmem_U8468 ( .A1(MEM_stage_inst_dmem_n8359), .A2(MEM_stage_inst_dmem_n8358), .ZN(MEM_stage_inst_dmem_n8363) );
NAND2_X1 MEM_stage_inst_dmem_U8467 ( .A1(MEM_stage_inst_dmem_ram_3567), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n8358) );
NAND2_X1 MEM_stage_inst_dmem_U8466 ( .A1(MEM_stage_inst_dmem_ram_3487), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n8359) );
NOR2_X1 MEM_stage_inst_dmem_U8465 ( .A1(MEM_stage_inst_dmem_n8357), .A2(MEM_stage_inst_dmem_n8356), .ZN(MEM_stage_inst_dmem_n8365) );
NAND2_X1 MEM_stage_inst_dmem_U8464 ( .A1(MEM_stage_inst_dmem_n8355), .A2(MEM_stage_inst_dmem_n8354), .ZN(MEM_stage_inst_dmem_n8356) );
NAND2_X1 MEM_stage_inst_dmem_U8463 ( .A1(MEM_stage_inst_dmem_ram_3439), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n8354) );
NAND2_X1 MEM_stage_inst_dmem_U8462 ( .A1(MEM_stage_inst_dmem_ram_3647), .A2(MEM_stage_inst_dmem_n41), .ZN(MEM_stage_inst_dmem_n8355) );
NAND2_X1 MEM_stage_inst_dmem_U8461 ( .A1(MEM_stage_inst_dmem_n8353), .A2(MEM_stage_inst_dmem_n8352), .ZN(MEM_stage_inst_dmem_n8357) );
NAND2_X1 MEM_stage_inst_dmem_U8460 ( .A1(MEM_stage_inst_dmem_ram_3919), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n8352) );
NAND2_X1 MEM_stage_inst_dmem_U8459 ( .A1(MEM_stage_inst_dmem_ram_3311), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n8353) );
NAND2_X1 MEM_stage_inst_dmem_U8458 ( .A1(MEM_stage_inst_dmem_n8351), .A2(MEM_stage_inst_dmem_n8350), .ZN(MEM_stage_inst_dmem_n8416) );
NOR2_X1 MEM_stage_inst_dmem_U8457 ( .A1(MEM_stage_inst_dmem_n8349), .A2(MEM_stage_inst_dmem_n8348), .ZN(MEM_stage_inst_dmem_n8350) );
NAND2_X1 MEM_stage_inst_dmem_U8456 ( .A1(MEM_stage_inst_dmem_n8347), .A2(MEM_stage_inst_dmem_n8346), .ZN(MEM_stage_inst_dmem_n8348) );
NOR2_X1 MEM_stage_inst_dmem_U8455 ( .A1(MEM_stage_inst_dmem_n8345), .A2(MEM_stage_inst_dmem_n8344), .ZN(MEM_stage_inst_dmem_n8346) );
NAND2_X1 MEM_stage_inst_dmem_U8454 ( .A1(MEM_stage_inst_dmem_n8343), .A2(MEM_stage_inst_dmem_n8342), .ZN(MEM_stage_inst_dmem_n8344) );
NAND2_X1 MEM_stage_inst_dmem_U8453 ( .A1(MEM_stage_inst_dmem_ram_3615), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n8342) );
NAND2_X1 MEM_stage_inst_dmem_U8452 ( .A1(MEM_stage_inst_dmem_ram_3423), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n8343) );
NAND2_X1 MEM_stage_inst_dmem_U8451 ( .A1(MEM_stage_inst_dmem_n8341), .A2(MEM_stage_inst_dmem_n8340), .ZN(MEM_stage_inst_dmem_n8345) );
NAND2_X1 MEM_stage_inst_dmem_U8450 ( .A1(MEM_stage_inst_dmem_ram_3599), .A2(MEM_stage_inst_dmem_n71), .ZN(MEM_stage_inst_dmem_n8340) );
NAND2_X1 MEM_stage_inst_dmem_U8449 ( .A1(MEM_stage_inst_dmem_ram_3679), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n8341) );
NOR2_X1 MEM_stage_inst_dmem_U8448 ( .A1(MEM_stage_inst_dmem_n8339), .A2(MEM_stage_inst_dmem_n8338), .ZN(MEM_stage_inst_dmem_n8347) );
NAND2_X1 MEM_stage_inst_dmem_U8447 ( .A1(MEM_stage_inst_dmem_n8337), .A2(MEM_stage_inst_dmem_n8336), .ZN(MEM_stage_inst_dmem_n8338) );
NAND2_X1 MEM_stage_inst_dmem_U8446 ( .A1(MEM_stage_inst_dmem_ram_3375), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n8336) );
NAND2_X1 MEM_stage_inst_dmem_U8445 ( .A1(MEM_stage_inst_dmem_ram_3247), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n8337) );
NAND2_X1 MEM_stage_inst_dmem_U8444 ( .A1(MEM_stage_inst_dmem_n8335), .A2(MEM_stage_inst_dmem_n8334), .ZN(MEM_stage_inst_dmem_n8339) );
NAND2_X1 MEM_stage_inst_dmem_U8443 ( .A1(MEM_stage_inst_dmem_ram_3711), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n8334) );
NAND2_X1 MEM_stage_inst_dmem_U8442 ( .A1(MEM_stage_inst_dmem_ram_3871), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n8335) );
NAND2_X1 MEM_stage_inst_dmem_U8441 ( .A1(MEM_stage_inst_dmem_n8333), .A2(MEM_stage_inst_dmem_n8332), .ZN(MEM_stage_inst_dmem_n8349) );
NOR2_X1 MEM_stage_inst_dmem_U8440 ( .A1(MEM_stage_inst_dmem_n8331), .A2(MEM_stage_inst_dmem_n8330), .ZN(MEM_stage_inst_dmem_n8332) );
NAND2_X1 MEM_stage_inst_dmem_U8439 ( .A1(MEM_stage_inst_dmem_n8329), .A2(MEM_stage_inst_dmem_n8328), .ZN(MEM_stage_inst_dmem_n8330) );
NAND2_X1 MEM_stage_inst_dmem_U8438 ( .A1(MEM_stage_inst_dmem_n27), .A2(MEM_stage_inst_dmem_ram_3663), .ZN(MEM_stage_inst_dmem_n8328) );
NAND2_X1 MEM_stage_inst_dmem_U8437 ( .A1(MEM_stage_inst_dmem_n7898), .A2(MEM_stage_inst_dmem_ram_3343), .ZN(MEM_stage_inst_dmem_n8329) );
NAND2_X1 MEM_stage_inst_dmem_U8436 ( .A1(MEM_stage_inst_dmem_n8327), .A2(MEM_stage_inst_dmem_n8326), .ZN(MEM_stage_inst_dmem_n8331) );
NAND2_X1 MEM_stage_inst_dmem_U8435 ( .A1(MEM_stage_inst_dmem_ram_3743), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n8326) );
NAND2_X1 MEM_stage_inst_dmem_U8434 ( .A1(MEM_stage_inst_dmem_ram_3823), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n8327) );
NOR2_X1 MEM_stage_inst_dmem_U8433 ( .A1(MEM_stage_inst_dmem_n8324), .A2(MEM_stage_inst_dmem_n8323), .ZN(MEM_stage_inst_dmem_n8333) );
NAND2_X1 MEM_stage_inst_dmem_U8432 ( .A1(MEM_stage_inst_dmem_n8322), .A2(MEM_stage_inst_dmem_n8321), .ZN(MEM_stage_inst_dmem_n8323) );
NAND2_X1 MEM_stage_inst_dmem_U8431 ( .A1(MEM_stage_inst_dmem_ram_3087), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n8321) );
NAND2_X1 MEM_stage_inst_dmem_U8430 ( .A1(MEM_stage_inst_dmem_ram_3807), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n8322) );
NAND2_X1 MEM_stage_inst_dmem_U8429 ( .A1(MEM_stage_inst_dmem_n8320), .A2(MEM_stage_inst_dmem_n8319), .ZN(MEM_stage_inst_dmem_n8324) );
NAND2_X1 MEM_stage_inst_dmem_U8428 ( .A1(MEM_stage_inst_dmem_ram_3455), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n8319) );
NAND2_X1 MEM_stage_inst_dmem_U8427 ( .A1(MEM_stage_inst_dmem_ram_3183), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n8320) );
NOR2_X1 MEM_stage_inst_dmem_U8426 ( .A1(MEM_stage_inst_dmem_n8318), .A2(MEM_stage_inst_dmem_n8317), .ZN(MEM_stage_inst_dmem_n8351) );
NAND2_X1 MEM_stage_inst_dmem_U8425 ( .A1(MEM_stage_inst_dmem_n8316), .A2(MEM_stage_inst_dmem_n8315), .ZN(MEM_stage_inst_dmem_n8317) );
NOR2_X1 MEM_stage_inst_dmem_U8424 ( .A1(MEM_stage_inst_dmem_n8314), .A2(MEM_stage_inst_dmem_n8313), .ZN(MEM_stage_inst_dmem_n8315) );
NAND2_X1 MEM_stage_inst_dmem_U8423 ( .A1(MEM_stage_inst_dmem_n8312), .A2(MEM_stage_inst_dmem_n8311), .ZN(MEM_stage_inst_dmem_n8313) );
NAND2_X1 MEM_stage_inst_dmem_U8422 ( .A1(MEM_stage_inst_dmem_n70), .A2(MEM_stage_inst_dmem_ram_3103), .ZN(MEM_stage_inst_dmem_n8311) );
NAND2_X1 MEM_stage_inst_dmem_U8421 ( .A1(MEM_stage_inst_dmem_n50), .A2(MEM_stage_inst_dmem_ram_3775), .ZN(MEM_stage_inst_dmem_n8312) );
NAND2_X1 MEM_stage_inst_dmem_U8420 ( .A1(MEM_stage_inst_dmem_n8310), .A2(MEM_stage_inst_dmem_n8309), .ZN(MEM_stage_inst_dmem_n8314) );
NAND2_X1 MEM_stage_inst_dmem_U8419 ( .A1(MEM_stage_inst_dmem_ram_3167), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n8309) );
NAND2_X1 MEM_stage_inst_dmem_U8418 ( .A1(MEM_stage_inst_dmem_ram_3551), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n8310) );
NOR2_X1 MEM_stage_inst_dmem_U8417 ( .A1(MEM_stage_inst_dmem_n8308), .A2(MEM_stage_inst_dmem_n8307), .ZN(MEM_stage_inst_dmem_n8316) );
NAND2_X1 MEM_stage_inst_dmem_U8416 ( .A1(MEM_stage_inst_dmem_n8306), .A2(MEM_stage_inst_dmem_n8305), .ZN(MEM_stage_inst_dmem_n8307) );
NAND2_X1 MEM_stage_inst_dmem_U8415 ( .A1(MEM_stage_inst_dmem_ram_3887), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n8305) );
NAND2_X1 MEM_stage_inst_dmem_U8414 ( .A1(MEM_stage_inst_dmem_ram_3759), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n8306) );
NAND2_X1 MEM_stage_inst_dmem_U8413 ( .A1(MEM_stage_inst_dmem_n8304), .A2(MEM_stage_inst_dmem_n8303), .ZN(MEM_stage_inst_dmem_n8308) );
NAND2_X1 MEM_stage_inst_dmem_U8412 ( .A1(MEM_stage_inst_dmem_n52), .A2(MEM_stage_inst_dmem_ram_3199), .ZN(MEM_stage_inst_dmem_n8303) );
NAND2_X1 MEM_stage_inst_dmem_U8411 ( .A1(MEM_stage_inst_dmem_n46), .A2(MEM_stage_inst_dmem_ram_3903), .ZN(MEM_stage_inst_dmem_n8304) );
NAND2_X1 MEM_stage_inst_dmem_U8410 ( .A1(MEM_stage_inst_dmem_n8302), .A2(MEM_stage_inst_dmem_n8301), .ZN(MEM_stage_inst_dmem_n8318) );
NOR2_X1 MEM_stage_inst_dmem_U8409 ( .A1(MEM_stage_inst_dmem_n8300), .A2(MEM_stage_inst_dmem_n8299), .ZN(MEM_stage_inst_dmem_n8301) );
NAND2_X1 MEM_stage_inst_dmem_U8408 ( .A1(MEM_stage_inst_dmem_n8298), .A2(MEM_stage_inst_dmem_n8297), .ZN(MEM_stage_inst_dmem_n8299) );
NAND2_X1 MEM_stage_inst_dmem_U8407 ( .A1(MEM_stage_inst_dmem_n76), .A2(MEM_stage_inst_dmem_ram_4015), .ZN(MEM_stage_inst_dmem_n8297) );
NAND2_X1 MEM_stage_inst_dmem_U8406 ( .A1(MEM_stage_inst_dmem_n44), .A2(MEM_stage_inst_dmem_ram_3231), .ZN(MEM_stage_inst_dmem_n8298) );
NAND2_X1 MEM_stage_inst_dmem_U8405 ( .A1(MEM_stage_inst_dmem_n8296), .A2(MEM_stage_inst_dmem_n8295), .ZN(MEM_stage_inst_dmem_n8300) );
NAND2_X1 MEM_stage_inst_dmem_U8404 ( .A1(MEM_stage_inst_dmem_ram_3695), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n8295) );
NAND2_X1 MEM_stage_inst_dmem_U8403 ( .A1(MEM_stage_inst_dmem_ram_3263), .A2(MEM_stage_inst_dmem_n8434), .ZN(MEM_stage_inst_dmem_n8296) );
NOR2_X1 MEM_stage_inst_dmem_U8402 ( .A1(MEM_stage_inst_dmem_n8294), .A2(MEM_stage_inst_dmem_n8293), .ZN(MEM_stage_inst_dmem_n8302) );
NAND2_X1 MEM_stage_inst_dmem_U8401 ( .A1(MEM_stage_inst_dmem_n8292), .A2(MEM_stage_inst_dmem_n8291), .ZN(MEM_stage_inst_dmem_n8293) );
NAND2_X1 MEM_stage_inst_dmem_U8400 ( .A1(MEM_stage_inst_dmem_ram_3471), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n8291) );
NAND2_X1 MEM_stage_inst_dmem_U8399 ( .A1(MEM_stage_inst_dmem_ram_3295), .A2(MEM_stage_inst_dmem_n51), .ZN(MEM_stage_inst_dmem_n8292) );
NAND2_X1 MEM_stage_inst_dmem_U8398 ( .A1(MEM_stage_inst_dmem_n8290), .A2(MEM_stage_inst_dmem_n8289), .ZN(MEM_stage_inst_dmem_n8294) );
NAND2_X1 MEM_stage_inst_dmem_U8397 ( .A1(MEM_stage_inst_dmem_ram_4095), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n8289) );
NAND2_X1 MEM_stage_inst_dmem_U8396 ( .A1(MEM_stage_inst_dmem_ram_3535), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n8290) );
NOR2_X1 MEM_stage_inst_dmem_U8395 ( .A1(MEM_stage_inst_dmem_n8288), .A2(MEM_stage_inst_dmem_n8287), .ZN(MEM_stage_inst_dmem_n8555) );
NOR2_X1 MEM_stage_inst_dmem_U8394 ( .A1(MEM_stage_inst_dmem_n8286), .A2(MEM_stage_inst_dmem_n8285), .ZN(MEM_stage_inst_dmem_n8287) );
NOR2_X1 MEM_stage_inst_dmem_U8393 ( .A1(MEM_stage_inst_dmem_n8284), .A2(MEM_stage_inst_dmem_n8283), .ZN(MEM_stage_inst_dmem_n8285) );
NAND2_X1 MEM_stage_inst_dmem_U8392 ( .A1(MEM_stage_inst_dmem_n8282), .A2(MEM_stage_inst_dmem_n8281), .ZN(MEM_stage_inst_dmem_n8283) );
NOR2_X1 MEM_stage_inst_dmem_U8391 ( .A1(MEM_stage_inst_dmem_n8280), .A2(MEM_stage_inst_dmem_n8279), .ZN(MEM_stage_inst_dmem_n8281) );
NAND2_X1 MEM_stage_inst_dmem_U8390 ( .A1(MEM_stage_inst_dmem_n8278), .A2(MEM_stage_inst_dmem_n8277), .ZN(MEM_stage_inst_dmem_n8279) );
NOR2_X1 MEM_stage_inst_dmem_U8389 ( .A1(MEM_stage_inst_dmem_n8276), .A2(MEM_stage_inst_dmem_n8275), .ZN(MEM_stage_inst_dmem_n8277) );
NAND2_X1 MEM_stage_inst_dmem_U8388 ( .A1(MEM_stage_inst_dmem_n8274), .A2(MEM_stage_inst_dmem_n8273), .ZN(MEM_stage_inst_dmem_n8275) );
NAND2_X1 MEM_stage_inst_dmem_U8387 ( .A1(MEM_stage_inst_dmem_ram_2911), .A2(MEM_stage_inst_dmem_n3141), .ZN(MEM_stage_inst_dmem_n8273) );
NAND2_X1 MEM_stage_inst_dmem_U8386 ( .A1(MEM_stage_inst_dmem_ram_3055), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n8274) );
NAND2_X1 MEM_stage_inst_dmem_U8385 ( .A1(MEM_stage_inst_dmem_n8272), .A2(MEM_stage_inst_dmem_n8271), .ZN(MEM_stage_inst_dmem_n8276) );
NAND2_X1 MEM_stage_inst_dmem_U8384 ( .A1(MEM_stage_inst_dmem_ram_2559), .A2(MEM_stage_inst_dmem_n64), .ZN(MEM_stage_inst_dmem_n8271) );
NAND2_X1 MEM_stage_inst_dmem_U8383 ( .A1(MEM_stage_inst_dmem_ram_2511), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n8272) );
NOR2_X1 MEM_stage_inst_dmem_U8382 ( .A1(MEM_stage_inst_dmem_n8270), .A2(MEM_stage_inst_dmem_n8269), .ZN(MEM_stage_inst_dmem_n8278) );
NAND2_X1 MEM_stage_inst_dmem_U8381 ( .A1(MEM_stage_inst_dmem_n8268), .A2(MEM_stage_inst_dmem_n8267), .ZN(MEM_stage_inst_dmem_n8269) );
NAND2_X1 MEM_stage_inst_dmem_U8380 ( .A1(MEM_stage_inst_dmem_ram_2079), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n8267) );
NAND2_X1 MEM_stage_inst_dmem_U8379 ( .A1(MEM_stage_inst_dmem_ram_2399), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n8268) );
NAND2_X1 MEM_stage_inst_dmem_U8378 ( .A1(MEM_stage_inst_dmem_n8266), .A2(MEM_stage_inst_dmem_n8265), .ZN(MEM_stage_inst_dmem_n8270) );
NAND2_X1 MEM_stage_inst_dmem_U8377 ( .A1(MEM_stage_inst_dmem_ram_2831), .A2(MEM_stage_inst_dmem_n8472), .ZN(MEM_stage_inst_dmem_n8265) );
NAND2_X1 MEM_stage_inst_dmem_U8376 ( .A1(MEM_stage_inst_dmem_ram_2975), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n8266) );
NAND2_X1 MEM_stage_inst_dmem_U8375 ( .A1(MEM_stage_inst_dmem_n8264), .A2(MEM_stage_inst_dmem_n8263), .ZN(MEM_stage_inst_dmem_n8280) );
NOR2_X1 MEM_stage_inst_dmem_U8374 ( .A1(MEM_stage_inst_dmem_n8262), .A2(MEM_stage_inst_dmem_n8261), .ZN(MEM_stage_inst_dmem_n8263) );
NAND2_X1 MEM_stage_inst_dmem_U8373 ( .A1(MEM_stage_inst_dmem_n8260), .A2(MEM_stage_inst_dmem_n8259), .ZN(MEM_stage_inst_dmem_n8261) );
NAND2_X1 MEM_stage_inst_dmem_U8372 ( .A1(MEM_stage_inst_dmem_ram_2127), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n8259) );
NAND2_X1 MEM_stage_inst_dmem_U8371 ( .A1(MEM_stage_inst_dmem_ram_2175), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n8260) );
NAND2_X1 MEM_stage_inst_dmem_U8370 ( .A1(MEM_stage_inst_dmem_n8258), .A2(MEM_stage_inst_dmem_n8257), .ZN(MEM_stage_inst_dmem_n8262) );
NAND2_X1 MEM_stage_inst_dmem_U8369 ( .A1(MEM_stage_inst_dmem_ram_2943), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n8257) );
NAND2_X1 MEM_stage_inst_dmem_U8368 ( .A1(MEM_stage_inst_dmem_ram_2255), .A2(MEM_stage_inst_dmem_n8256), .ZN(MEM_stage_inst_dmem_n8258) );
NOR2_X1 MEM_stage_inst_dmem_U8367 ( .A1(MEM_stage_inst_dmem_n8255), .A2(MEM_stage_inst_dmem_n8254), .ZN(MEM_stage_inst_dmem_n8264) );
NAND2_X1 MEM_stage_inst_dmem_U8366 ( .A1(MEM_stage_inst_dmem_n8253), .A2(MEM_stage_inst_dmem_n8252), .ZN(MEM_stage_inst_dmem_n8254) );
NAND2_X1 MEM_stage_inst_dmem_U8365 ( .A1(MEM_stage_inst_dmem_ram_2415), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n8252) );
NAND2_X1 MEM_stage_inst_dmem_U8364 ( .A1(MEM_stage_inst_dmem_ram_2287), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n8253) );
NAND2_X1 MEM_stage_inst_dmem_U8363 ( .A1(MEM_stage_inst_dmem_n8251), .A2(MEM_stage_inst_dmem_n8250), .ZN(MEM_stage_inst_dmem_n8255) );
NAND2_X1 MEM_stage_inst_dmem_U8362 ( .A1(MEM_stage_inst_dmem_n8421), .A2(MEM_stage_inst_dmem_ram_2479), .ZN(MEM_stage_inst_dmem_n8250) );
NAND2_X1 MEM_stage_inst_dmem_U8361 ( .A1(MEM_stage_inst_dmem_n75), .A2(MEM_stage_inst_dmem_ram_2447), .ZN(MEM_stage_inst_dmem_n8251) );
NOR2_X1 MEM_stage_inst_dmem_U8360 ( .A1(MEM_stage_inst_dmem_n8249), .A2(MEM_stage_inst_dmem_n8248), .ZN(MEM_stage_inst_dmem_n8282) );
NAND2_X1 MEM_stage_inst_dmem_U8359 ( .A1(MEM_stage_inst_dmem_n8247), .A2(MEM_stage_inst_dmem_n8246), .ZN(MEM_stage_inst_dmem_n8248) );
NOR2_X1 MEM_stage_inst_dmem_U8358 ( .A1(MEM_stage_inst_dmem_n8245), .A2(MEM_stage_inst_dmem_n8244), .ZN(MEM_stage_inst_dmem_n8246) );
NAND2_X1 MEM_stage_inst_dmem_U8357 ( .A1(MEM_stage_inst_dmem_n8243), .A2(MEM_stage_inst_dmem_n8242), .ZN(MEM_stage_inst_dmem_n8244) );
NAND2_X1 MEM_stage_inst_dmem_U8356 ( .A1(MEM_stage_inst_dmem_ram_2335), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n8242) );
NAND2_X1 MEM_stage_inst_dmem_U8355 ( .A1(MEM_stage_inst_dmem_ram_2719), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n8243) );
NAND2_X1 MEM_stage_inst_dmem_U8354 ( .A1(MEM_stage_inst_dmem_n8241), .A2(MEM_stage_inst_dmem_n8240), .ZN(MEM_stage_inst_dmem_n8245) );
NAND2_X1 MEM_stage_inst_dmem_U8353 ( .A1(MEM_stage_inst_dmem_ram_2223), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n8240) );
NAND2_X1 MEM_stage_inst_dmem_U8352 ( .A1(MEM_stage_inst_dmem_ram_2655), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n8241) );
NOR2_X1 MEM_stage_inst_dmem_U8351 ( .A1(MEM_stage_inst_dmem_n8239), .A2(MEM_stage_inst_dmem_n8238), .ZN(MEM_stage_inst_dmem_n8247) );
NAND2_X1 MEM_stage_inst_dmem_U8350 ( .A1(MEM_stage_inst_dmem_n8237), .A2(MEM_stage_inst_dmem_n8236), .ZN(MEM_stage_inst_dmem_n8238) );
NAND2_X1 MEM_stage_inst_dmem_U8349 ( .A1(MEM_stage_inst_dmem_ram_2111), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n8236) );
NAND2_X1 MEM_stage_inst_dmem_U8348 ( .A1(MEM_stage_inst_dmem_ram_2143), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n8237) );
NAND2_X1 MEM_stage_inst_dmem_U8347 ( .A1(MEM_stage_inst_dmem_n8235), .A2(MEM_stage_inst_dmem_n8234), .ZN(MEM_stage_inst_dmem_n8239) );
NAND2_X1 MEM_stage_inst_dmem_U8346 ( .A1(MEM_stage_inst_dmem_ram_2863), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n8234) );
NAND2_X1 MEM_stage_inst_dmem_U8345 ( .A1(MEM_stage_inst_dmem_ram_2239), .A2(MEM_stage_inst_dmem_n8434), .ZN(MEM_stage_inst_dmem_n8235) );
NAND2_X1 MEM_stage_inst_dmem_U8344 ( .A1(MEM_stage_inst_dmem_n8233), .A2(MEM_stage_inst_dmem_n8232), .ZN(MEM_stage_inst_dmem_n8249) );
NOR2_X1 MEM_stage_inst_dmem_U8343 ( .A1(MEM_stage_inst_dmem_n8231), .A2(MEM_stage_inst_dmem_n8230), .ZN(MEM_stage_inst_dmem_n8232) );
NAND2_X1 MEM_stage_inst_dmem_U8342 ( .A1(MEM_stage_inst_dmem_n8229), .A2(MEM_stage_inst_dmem_n8228), .ZN(MEM_stage_inst_dmem_n8230) );
NAND2_X1 MEM_stage_inst_dmem_U8341 ( .A1(MEM_stage_inst_dmem_ram_2383), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n8228) );
NAND2_X1 MEM_stage_inst_dmem_U8340 ( .A1(MEM_stage_inst_dmem_ram_2095), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n8229) );
NAND2_X1 MEM_stage_inst_dmem_U8339 ( .A1(MEM_stage_inst_dmem_n8227), .A2(MEM_stage_inst_dmem_n8226), .ZN(MEM_stage_inst_dmem_n8231) );
NAND2_X1 MEM_stage_inst_dmem_U8338 ( .A1(MEM_stage_inst_dmem_ram_2575), .A2(MEM_stage_inst_dmem_n8225), .ZN(MEM_stage_inst_dmem_n8226) );
NAND2_X1 MEM_stage_inst_dmem_U8337 ( .A1(MEM_stage_inst_dmem_ram_2783), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n8227) );
NOR2_X1 MEM_stage_inst_dmem_U8336 ( .A1(MEM_stage_inst_dmem_n8224), .A2(MEM_stage_inst_dmem_n8223), .ZN(MEM_stage_inst_dmem_n8233) );
NAND2_X1 MEM_stage_inst_dmem_U8335 ( .A1(MEM_stage_inst_dmem_n8222), .A2(MEM_stage_inst_dmem_n8221), .ZN(MEM_stage_inst_dmem_n8223) );
NAND2_X1 MEM_stage_inst_dmem_U8334 ( .A1(MEM_stage_inst_dmem_ram_2895), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n8221) );
NAND2_X1 MEM_stage_inst_dmem_U8333 ( .A1(MEM_stage_inst_dmem_ram_2159), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n8222) );
NAND2_X1 MEM_stage_inst_dmem_U8332 ( .A1(MEM_stage_inst_dmem_n8220), .A2(MEM_stage_inst_dmem_n8219), .ZN(MEM_stage_inst_dmem_n8224) );
NAND2_X1 MEM_stage_inst_dmem_U8331 ( .A1(MEM_stage_inst_dmem_ram_2767), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n8219) );
NAND2_X1 MEM_stage_inst_dmem_U8330 ( .A1(MEM_stage_inst_dmem_ram_2319), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n8220) );
NAND2_X1 MEM_stage_inst_dmem_U8329 ( .A1(MEM_stage_inst_dmem_n8218), .A2(MEM_stage_inst_dmem_n8217), .ZN(MEM_stage_inst_dmem_n8284) );
NOR2_X1 MEM_stage_inst_dmem_U8328 ( .A1(MEM_stage_inst_dmem_n8216), .A2(MEM_stage_inst_dmem_n8215), .ZN(MEM_stage_inst_dmem_n8217) );
NAND2_X1 MEM_stage_inst_dmem_U8327 ( .A1(MEM_stage_inst_dmem_n8214), .A2(MEM_stage_inst_dmem_n8213), .ZN(MEM_stage_inst_dmem_n8215) );
NOR2_X1 MEM_stage_inst_dmem_U8326 ( .A1(MEM_stage_inst_dmem_n8212), .A2(MEM_stage_inst_dmem_n8211), .ZN(MEM_stage_inst_dmem_n8213) );
NAND2_X1 MEM_stage_inst_dmem_U8325 ( .A1(MEM_stage_inst_dmem_n8210), .A2(MEM_stage_inst_dmem_n8209), .ZN(MEM_stage_inst_dmem_n8211) );
NAND2_X1 MEM_stage_inst_dmem_U8324 ( .A1(MEM_stage_inst_dmem_n27), .A2(MEM_stage_inst_dmem_ram_2639), .ZN(MEM_stage_inst_dmem_n8209) );
NAND2_X1 MEM_stage_inst_dmem_U8323 ( .A1(MEM_stage_inst_dmem_n32), .A2(MEM_stage_inst_dmem_ram_2687), .ZN(MEM_stage_inst_dmem_n8210) );
NAND2_X1 MEM_stage_inst_dmem_U8322 ( .A1(MEM_stage_inst_dmem_n8208), .A2(MEM_stage_inst_dmem_n8207), .ZN(MEM_stage_inst_dmem_n8212) );
NAND2_X1 MEM_stage_inst_dmem_U8321 ( .A1(MEM_stage_inst_dmem_ram_2271), .A2(MEM_stage_inst_dmem_n8206), .ZN(MEM_stage_inst_dmem_n8207) );
NAND2_X1 MEM_stage_inst_dmem_U8320 ( .A1(MEM_stage_inst_dmem_ram_2799), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n8208) );
NOR2_X1 MEM_stage_inst_dmem_U8319 ( .A1(MEM_stage_inst_dmem_n8205), .A2(MEM_stage_inst_dmem_n8204), .ZN(MEM_stage_inst_dmem_n8214) );
NAND2_X1 MEM_stage_inst_dmem_U8318 ( .A1(MEM_stage_inst_dmem_n8203), .A2(MEM_stage_inst_dmem_n8202), .ZN(MEM_stage_inst_dmem_n8204) );
NAND2_X1 MEM_stage_inst_dmem_U8317 ( .A1(MEM_stage_inst_dmem_ram_2351), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n8202) );
NAND2_X1 MEM_stage_inst_dmem_U8316 ( .A1(MEM_stage_inst_dmem_ram_2063), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n8203) );
NAND2_X1 MEM_stage_inst_dmem_U8315 ( .A1(MEM_stage_inst_dmem_n8201), .A2(MEM_stage_inst_dmem_n8200), .ZN(MEM_stage_inst_dmem_n8205) );
NAND2_X1 MEM_stage_inst_dmem_U8314 ( .A1(MEM_stage_inst_dmem_n19), .A2(MEM_stage_inst_dmem_ram_2543), .ZN(MEM_stage_inst_dmem_n8200) );
NAND2_X1 MEM_stage_inst_dmem_U8313 ( .A1(MEM_stage_inst_dmem_n35), .A2(MEM_stage_inst_dmem_ram_3039), .ZN(MEM_stage_inst_dmem_n8201) );
NAND2_X1 MEM_stage_inst_dmem_U8312 ( .A1(MEM_stage_inst_dmem_n8199), .A2(MEM_stage_inst_dmem_n8198), .ZN(MEM_stage_inst_dmem_n8216) );
NOR2_X1 MEM_stage_inst_dmem_U8311 ( .A1(MEM_stage_inst_dmem_n8197), .A2(MEM_stage_inst_dmem_n8196), .ZN(MEM_stage_inst_dmem_n8198) );
NAND2_X1 MEM_stage_inst_dmem_U8310 ( .A1(MEM_stage_inst_dmem_n8195), .A2(MEM_stage_inst_dmem_n8194), .ZN(MEM_stage_inst_dmem_n8196) );
NAND2_X1 MEM_stage_inst_dmem_U8309 ( .A1(MEM_stage_inst_dmem_ram_2495), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n8194) );
NAND2_X1 MEM_stage_inst_dmem_U8308 ( .A1(MEM_stage_inst_dmem_ram_2959), .A2(MEM_stage_inst_dmem_n8193), .ZN(MEM_stage_inst_dmem_n8195) );
NAND2_X1 MEM_stage_inst_dmem_U8307 ( .A1(MEM_stage_inst_dmem_n8192), .A2(MEM_stage_inst_dmem_n8191), .ZN(MEM_stage_inst_dmem_n8197) );
NAND2_X1 MEM_stage_inst_dmem_U8306 ( .A1(MEM_stage_inst_dmem_ram_3023), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n8191) );
NAND2_X1 MEM_stage_inst_dmem_U8305 ( .A1(MEM_stage_inst_dmem_ram_2607), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n8192) );
NOR2_X1 MEM_stage_inst_dmem_U8304 ( .A1(MEM_stage_inst_dmem_n8190), .A2(MEM_stage_inst_dmem_n8189), .ZN(MEM_stage_inst_dmem_n8199) );
NAND2_X1 MEM_stage_inst_dmem_U8303 ( .A1(MEM_stage_inst_dmem_n8188), .A2(MEM_stage_inst_dmem_n8187), .ZN(MEM_stage_inst_dmem_n8189) );
NAND2_X1 MEM_stage_inst_dmem_U8302 ( .A1(MEM_stage_inst_dmem_ram_3007), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n8187) );
NAND2_X1 MEM_stage_inst_dmem_U8301 ( .A1(MEM_stage_inst_dmem_ram_2815), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n8188) );
NAND2_X1 MEM_stage_inst_dmem_U8300 ( .A1(MEM_stage_inst_dmem_n8186), .A2(MEM_stage_inst_dmem_n8185), .ZN(MEM_stage_inst_dmem_n8190) );
NAND2_X1 MEM_stage_inst_dmem_U8299 ( .A1(MEM_stage_inst_dmem_ram_2735), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n8185) );
NAND2_X1 MEM_stage_inst_dmem_U8298 ( .A1(MEM_stage_inst_dmem_ram_2847), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n8186) );
NOR2_X1 MEM_stage_inst_dmem_U8297 ( .A1(MEM_stage_inst_dmem_n8184), .A2(MEM_stage_inst_dmem_n8183), .ZN(MEM_stage_inst_dmem_n8218) );
NAND2_X1 MEM_stage_inst_dmem_U8296 ( .A1(MEM_stage_inst_dmem_n8182), .A2(MEM_stage_inst_dmem_n8181), .ZN(MEM_stage_inst_dmem_n8183) );
NOR2_X1 MEM_stage_inst_dmem_U8295 ( .A1(MEM_stage_inst_dmem_n8180), .A2(MEM_stage_inst_dmem_n8179), .ZN(MEM_stage_inst_dmem_n8181) );
NAND2_X1 MEM_stage_inst_dmem_U8294 ( .A1(MEM_stage_inst_dmem_n8178), .A2(MEM_stage_inst_dmem_n8177), .ZN(MEM_stage_inst_dmem_n8179) );
NAND2_X1 MEM_stage_inst_dmem_U8293 ( .A1(MEM_stage_inst_dmem_ram_3071), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n8177) );
NAND2_X1 MEM_stage_inst_dmem_U8292 ( .A1(MEM_stage_inst_dmem_ram_2207), .A2(MEM_stage_inst_dmem_n44), .ZN(MEM_stage_inst_dmem_n8178) );
NAND2_X1 MEM_stage_inst_dmem_U8291 ( .A1(MEM_stage_inst_dmem_n8176), .A2(MEM_stage_inst_dmem_n8175), .ZN(MEM_stage_inst_dmem_n8180) );
NAND2_X1 MEM_stage_inst_dmem_U8290 ( .A1(MEM_stage_inst_dmem_ram_2191), .A2(MEM_stage_inst_dmem_n8174), .ZN(MEM_stage_inst_dmem_n8175) );
NAND2_X1 MEM_stage_inst_dmem_U8289 ( .A1(MEM_stage_inst_dmem_ram_2527), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n8176) );
NOR2_X1 MEM_stage_inst_dmem_U8288 ( .A1(MEM_stage_inst_dmem_n8173), .A2(MEM_stage_inst_dmem_n8172), .ZN(MEM_stage_inst_dmem_n8182) );
NAND2_X1 MEM_stage_inst_dmem_U8287 ( .A1(MEM_stage_inst_dmem_n8171), .A2(MEM_stage_inst_dmem_n8170), .ZN(MEM_stage_inst_dmem_n8172) );
NAND2_X1 MEM_stage_inst_dmem_U8286 ( .A1(MEM_stage_inst_dmem_ram_2623), .A2(MEM_stage_inst_dmem_n8169), .ZN(MEM_stage_inst_dmem_n8170) );
NAND2_X1 MEM_stage_inst_dmem_U8285 ( .A1(MEM_stage_inst_dmem_ram_2463), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n8171) );
NAND2_X1 MEM_stage_inst_dmem_U8284 ( .A1(MEM_stage_inst_dmem_n8168), .A2(MEM_stage_inst_dmem_n8167), .ZN(MEM_stage_inst_dmem_n8173) );
NAND2_X1 MEM_stage_inst_dmem_U8283 ( .A1(MEM_stage_inst_dmem_n33), .A2(MEM_stage_inst_dmem_ram_2431), .ZN(MEM_stage_inst_dmem_n8167) );
NAND2_X1 MEM_stage_inst_dmem_U8282 ( .A1(MEM_stage_inst_dmem_n49), .A2(MEM_stage_inst_dmem_ram_2703), .ZN(MEM_stage_inst_dmem_n8168) );
NAND2_X1 MEM_stage_inst_dmem_U8281 ( .A1(MEM_stage_inst_dmem_n8166), .A2(MEM_stage_inst_dmem_n8165), .ZN(MEM_stage_inst_dmem_n8184) );
NOR2_X1 MEM_stage_inst_dmem_U8280 ( .A1(MEM_stage_inst_dmem_n8164), .A2(MEM_stage_inst_dmem_n8163), .ZN(MEM_stage_inst_dmem_n8165) );
NAND2_X1 MEM_stage_inst_dmem_U8279 ( .A1(MEM_stage_inst_dmem_n8162), .A2(MEM_stage_inst_dmem_n8161), .ZN(MEM_stage_inst_dmem_n8163) );
NAND2_X1 MEM_stage_inst_dmem_U8278 ( .A1(MEM_stage_inst_dmem_n76), .A2(MEM_stage_inst_dmem_ram_2991), .ZN(MEM_stage_inst_dmem_n8161) );
NAND2_X1 MEM_stage_inst_dmem_U8277 ( .A1(MEM_stage_inst_dmem_n45), .A2(MEM_stage_inst_dmem_ram_2591), .ZN(MEM_stage_inst_dmem_n8162) );
NAND2_X1 MEM_stage_inst_dmem_U8276 ( .A1(MEM_stage_inst_dmem_n8160), .A2(MEM_stage_inst_dmem_n8159), .ZN(MEM_stage_inst_dmem_n8164) );
NAND2_X1 MEM_stage_inst_dmem_U8275 ( .A1(MEM_stage_inst_dmem_ram_2367), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n8159) );
NAND2_X1 MEM_stage_inst_dmem_U8274 ( .A1(MEM_stage_inst_dmem_ram_2671), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n8160) );
NOR2_X1 MEM_stage_inst_dmem_U8273 ( .A1(MEM_stage_inst_dmem_n8158), .A2(MEM_stage_inst_dmem_n8157), .ZN(MEM_stage_inst_dmem_n8166) );
NAND2_X1 MEM_stage_inst_dmem_U8272 ( .A1(MEM_stage_inst_dmem_n8156), .A2(MEM_stage_inst_dmem_n8155), .ZN(MEM_stage_inst_dmem_n8157) );
NAND2_X1 MEM_stage_inst_dmem_U8271 ( .A1(MEM_stage_inst_dmem_n46), .A2(MEM_stage_inst_dmem_ram_2879), .ZN(MEM_stage_inst_dmem_n8155) );
NAND2_X1 MEM_stage_inst_dmem_U8270 ( .A1(MEM_stage_inst_dmem_n50), .A2(MEM_stage_inst_dmem_ram_2751), .ZN(MEM_stage_inst_dmem_n8156) );
NAND2_X1 MEM_stage_inst_dmem_U8269 ( .A1(MEM_stage_inst_dmem_n8154), .A2(MEM_stage_inst_dmem_n8153), .ZN(MEM_stage_inst_dmem_n8158) );
NAND2_X1 MEM_stage_inst_dmem_U8268 ( .A1(MEM_stage_inst_dmem_n63), .A2(MEM_stage_inst_dmem_ram_2927), .ZN(MEM_stage_inst_dmem_n8153) );
NAND2_X1 MEM_stage_inst_dmem_U8267 ( .A1(MEM_stage_inst_dmem_n39), .A2(MEM_stage_inst_dmem_ram_2303), .ZN(MEM_stage_inst_dmem_n8154) );
NOR2_X1 MEM_stage_inst_dmem_U8266 ( .A1(MEM_stage_inst_dmem_n8152), .A2(MEM_stage_inst_dmem_n8151), .ZN(MEM_stage_inst_dmem_n8288) );
NOR2_X1 MEM_stage_inst_dmem_U8265 ( .A1(MEM_stage_inst_dmem_n8150), .A2(MEM_stage_inst_dmem_n8149), .ZN(MEM_stage_inst_dmem_n8151) );
NAND2_X1 MEM_stage_inst_dmem_U8264 ( .A1(MEM_stage_inst_dmem_n8148), .A2(MEM_stage_inst_dmem_n8147), .ZN(MEM_stage_inst_dmem_n8149) );
NOR2_X1 MEM_stage_inst_dmem_U8263 ( .A1(MEM_stage_inst_dmem_n8146), .A2(MEM_stage_inst_dmem_n8145), .ZN(MEM_stage_inst_dmem_n8147) );
NAND2_X1 MEM_stage_inst_dmem_U8262 ( .A1(MEM_stage_inst_dmem_n8144), .A2(MEM_stage_inst_dmem_n8143), .ZN(MEM_stage_inst_dmem_n8145) );
NOR2_X1 MEM_stage_inst_dmem_U8261 ( .A1(MEM_stage_inst_dmem_n8142), .A2(MEM_stage_inst_dmem_n8141), .ZN(MEM_stage_inst_dmem_n8143) );
NAND2_X1 MEM_stage_inst_dmem_U8260 ( .A1(MEM_stage_inst_dmem_n8140), .A2(MEM_stage_inst_dmem_n8139), .ZN(MEM_stage_inst_dmem_n8141) );
NAND2_X1 MEM_stage_inst_dmem_U8259 ( .A1(MEM_stage_inst_dmem_ram_1183), .A2(MEM_stage_inst_dmem_n44), .ZN(MEM_stage_inst_dmem_n8139) );
NAND2_X1 MEM_stage_inst_dmem_U8258 ( .A1(MEM_stage_inst_dmem_ram_1375), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n8140) );
NAND2_X1 MEM_stage_inst_dmem_U8257 ( .A1(MEM_stage_inst_dmem_n8138), .A2(MEM_stage_inst_dmem_n8137), .ZN(MEM_stage_inst_dmem_n8142) );
NAND2_X1 MEM_stage_inst_dmem_U8256 ( .A1(MEM_stage_inst_dmem_ram_1903), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n8137) );
NAND2_X1 MEM_stage_inst_dmem_U8255 ( .A1(MEM_stage_inst_dmem_ram_1327), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n8138) );
NOR2_X1 MEM_stage_inst_dmem_U8254 ( .A1(MEM_stage_inst_dmem_n8136), .A2(MEM_stage_inst_dmem_n8135), .ZN(MEM_stage_inst_dmem_n8144) );
NAND2_X1 MEM_stage_inst_dmem_U8253 ( .A1(MEM_stage_inst_dmem_n8134), .A2(MEM_stage_inst_dmem_n8133), .ZN(MEM_stage_inst_dmem_n8135) );
NAND2_X1 MEM_stage_inst_dmem_U8252 ( .A1(MEM_stage_inst_dmem_ram_1535), .A2(MEM_stage_inst_dmem_n8535), .ZN(MEM_stage_inst_dmem_n8133) );
NAND2_X1 MEM_stage_inst_dmem_U8251 ( .A1(MEM_stage_inst_dmem_ram_1871), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n8134) );
NAND2_X1 MEM_stage_inst_dmem_U8250 ( .A1(MEM_stage_inst_dmem_n8132), .A2(MEM_stage_inst_dmem_n8131), .ZN(MEM_stage_inst_dmem_n8136) );
NAND2_X1 MEM_stage_inst_dmem_U8249 ( .A1(MEM_stage_inst_dmem_ram_1951), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n8131) );
NAND2_X1 MEM_stage_inst_dmem_U8248 ( .A1(MEM_stage_inst_dmem_ram_1791), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n8132) );
NAND2_X1 MEM_stage_inst_dmem_U8247 ( .A1(MEM_stage_inst_dmem_n8130), .A2(MEM_stage_inst_dmem_n8129), .ZN(MEM_stage_inst_dmem_n8146) );
NOR2_X1 MEM_stage_inst_dmem_U8246 ( .A1(MEM_stage_inst_dmem_n8128), .A2(MEM_stage_inst_dmem_n8127), .ZN(MEM_stage_inst_dmem_n8129) );
NAND2_X1 MEM_stage_inst_dmem_U8245 ( .A1(MEM_stage_inst_dmem_n8126), .A2(MEM_stage_inst_dmem_n8125), .ZN(MEM_stage_inst_dmem_n8127) );
NAND2_X1 MEM_stage_inst_dmem_U8244 ( .A1(MEM_stage_inst_dmem_ram_1471), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n8125) );
NAND2_X1 MEM_stage_inst_dmem_U8243 ( .A1(MEM_stage_inst_dmem_ram_1695), .A2(MEM_stage_inst_dmem_n3076), .ZN(MEM_stage_inst_dmem_n8126) );
NAND2_X1 MEM_stage_inst_dmem_U8242 ( .A1(MEM_stage_inst_dmem_n8124), .A2(MEM_stage_inst_dmem_n8123), .ZN(MEM_stage_inst_dmem_n8128) );
NAND2_X1 MEM_stage_inst_dmem_U8241 ( .A1(MEM_stage_inst_dmem_ram_1071), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n8123) );
NAND2_X1 MEM_stage_inst_dmem_U8240 ( .A1(MEM_stage_inst_dmem_ram_1423), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n8124) );
NOR2_X1 MEM_stage_inst_dmem_U8239 ( .A1(MEM_stage_inst_dmem_n8122), .A2(MEM_stage_inst_dmem_n8121), .ZN(MEM_stage_inst_dmem_n8130) );
NAND2_X1 MEM_stage_inst_dmem_U8238 ( .A1(MEM_stage_inst_dmem_n8120), .A2(MEM_stage_inst_dmem_n8119), .ZN(MEM_stage_inst_dmem_n8121) );
NAND2_X1 MEM_stage_inst_dmem_U8237 ( .A1(MEM_stage_inst_dmem_ram_1087), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n8119) );
NAND2_X1 MEM_stage_inst_dmem_U8236 ( .A1(MEM_stage_inst_dmem_ram_1615), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n8120) );
NAND2_X1 MEM_stage_inst_dmem_U8235 ( .A1(MEM_stage_inst_dmem_n8118), .A2(MEM_stage_inst_dmem_n8117), .ZN(MEM_stage_inst_dmem_n8122) );
NAND2_X1 MEM_stage_inst_dmem_U8234 ( .A1(MEM_stage_inst_dmem_ram_1935), .A2(MEM_stage_inst_dmem_n72), .ZN(MEM_stage_inst_dmem_n8117) );
NAND2_X1 MEM_stage_inst_dmem_U8233 ( .A1(MEM_stage_inst_dmem_ram_1119), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n8118) );
NOR2_X1 MEM_stage_inst_dmem_U8232 ( .A1(MEM_stage_inst_dmem_n8116), .A2(MEM_stage_inst_dmem_n8115), .ZN(MEM_stage_inst_dmem_n8148) );
NAND2_X1 MEM_stage_inst_dmem_U8231 ( .A1(MEM_stage_inst_dmem_n8114), .A2(MEM_stage_inst_dmem_n8113), .ZN(MEM_stage_inst_dmem_n8115) );
NOR2_X1 MEM_stage_inst_dmem_U8230 ( .A1(MEM_stage_inst_dmem_n8112), .A2(MEM_stage_inst_dmem_n8111), .ZN(MEM_stage_inst_dmem_n8113) );
NAND2_X1 MEM_stage_inst_dmem_U8229 ( .A1(MEM_stage_inst_dmem_n8110), .A2(MEM_stage_inst_dmem_n8109), .ZN(MEM_stage_inst_dmem_n8111) );
NAND2_X1 MEM_stage_inst_dmem_U8228 ( .A1(MEM_stage_inst_dmem_ram_1487), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n8109) );
NAND2_X1 MEM_stage_inst_dmem_U8227 ( .A1(MEM_stage_inst_dmem_ram_1823), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n8110) );
NAND2_X1 MEM_stage_inst_dmem_U8226 ( .A1(MEM_stage_inst_dmem_n8108), .A2(MEM_stage_inst_dmem_n8107), .ZN(MEM_stage_inst_dmem_n8112) );
NAND2_X1 MEM_stage_inst_dmem_U8225 ( .A1(MEM_stage_inst_dmem_ram_1055), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n8107) );
NAND2_X1 MEM_stage_inst_dmem_U8224 ( .A1(MEM_stage_inst_dmem_ram_1215), .A2(MEM_stage_inst_dmem_n8434), .ZN(MEM_stage_inst_dmem_n8108) );
NOR2_X1 MEM_stage_inst_dmem_U8223 ( .A1(MEM_stage_inst_dmem_n8106), .A2(MEM_stage_inst_dmem_n8105), .ZN(MEM_stage_inst_dmem_n8114) );
NAND2_X1 MEM_stage_inst_dmem_U8222 ( .A1(MEM_stage_inst_dmem_n8104), .A2(MEM_stage_inst_dmem_n8103), .ZN(MEM_stage_inst_dmem_n8105) );
NAND2_X1 MEM_stage_inst_dmem_U8221 ( .A1(MEM_stage_inst_dmem_ram_2015), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n8103) );
NAND2_X1 MEM_stage_inst_dmem_U8220 ( .A1(MEM_stage_inst_dmem_ram_1039), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n8104) );
NAND2_X1 MEM_stage_inst_dmem_U8219 ( .A1(MEM_stage_inst_dmem_n8102), .A2(MEM_stage_inst_dmem_n8101), .ZN(MEM_stage_inst_dmem_n8106) );
NAND2_X1 MEM_stage_inst_dmem_U8218 ( .A1(MEM_stage_inst_dmem_ram_1263), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n8101) );
NAND2_X1 MEM_stage_inst_dmem_U8217 ( .A1(MEM_stage_inst_dmem_ram_2047), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n8102) );
NAND2_X1 MEM_stage_inst_dmem_U8216 ( .A1(MEM_stage_inst_dmem_n8100), .A2(MEM_stage_inst_dmem_n8099), .ZN(MEM_stage_inst_dmem_n8116) );
NOR2_X1 MEM_stage_inst_dmem_U8215 ( .A1(MEM_stage_inst_dmem_n8098), .A2(MEM_stage_inst_dmem_n8097), .ZN(MEM_stage_inst_dmem_n8099) );
NAND2_X1 MEM_stage_inst_dmem_U8214 ( .A1(MEM_stage_inst_dmem_n8096), .A2(MEM_stage_inst_dmem_n8095), .ZN(MEM_stage_inst_dmem_n8097) );
NAND2_X1 MEM_stage_inst_dmem_U8213 ( .A1(MEM_stage_inst_dmem_n62), .A2(MEM_stage_inst_dmem_ram_1311), .ZN(MEM_stage_inst_dmem_n8095) );
NAND2_X1 MEM_stage_inst_dmem_U8212 ( .A1(MEM_stage_inst_dmem_n8421), .A2(MEM_stage_inst_dmem_ram_1455), .ZN(MEM_stage_inst_dmem_n8096) );
NAND2_X1 MEM_stage_inst_dmem_U8211 ( .A1(MEM_stage_inst_dmem_n8094), .A2(MEM_stage_inst_dmem_n8093), .ZN(MEM_stage_inst_dmem_n8098) );
NAND2_X1 MEM_stage_inst_dmem_U8210 ( .A1(MEM_stage_inst_dmem_ram_1807), .A2(MEM_stage_inst_dmem_n8472), .ZN(MEM_stage_inst_dmem_n8093) );
NAND2_X1 MEM_stage_inst_dmem_U8209 ( .A1(MEM_stage_inst_dmem_ram_1199), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n8094) );
NOR2_X1 MEM_stage_inst_dmem_U8208 ( .A1(MEM_stage_inst_dmem_n8092), .A2(MEM_stage_inst_dmem_n8091), .ZN(MEM_stage_inst_dmem_n8100) );
NAND2_X1 MEM_stage_inst_dmem_U8207 ( .A1(MEM_stage_inst_dmem_n8090), .A2(MEM_stage_inst_dmem_n8089), .ZN(MEM_stage_inst_dmem_n8091) );
NAND2_X1 MEM_stage_inst_dmem_U8206 ( .A1(MEM_stage_inst_dmem_ram_1599), .A2(MEM_stage_inst_dmem_n41), .ZN(MEM_stage_inst_dmem_n8089) );
NAND2_X1 MEM_stage_inst_dmem_U8205 ( .A1(MEM_stage_inst_dmem_ram_1759), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n8090) );
NAND2_X1 MEM_stage_inst_dmem_U8204 ( .A1(MEM_stage_inst_dmem_n8088), .A2(MEM_stage_inst_dmem_n8087), .ZN(MEM_stage_inst_dmem_n8092) );
NAND2_X1 MEM_stage_inst_dmem_U8203 ( .A1(MEM_stage_inst_dmem_n32), .A2(MEM_stage_inst_dmem_ram_1663), .ZN(MEM_stage_inst_dmem_n8087) );
NAND2_X1 MEM_stage_inst_dmem_U8202 ( .A1(MEM_stage_inst_dmem_n52), .A2(MEM_stage_inst_dmem_ram_1151), .ZN(MEM_stage_inst_dmem_n8088) );
NAND2_X1 MEM_stage_inst_dmem_U8201 ( .A1(MEM_stage_inst_dmem_n8086), .A2(MEM_stage_inst_dmem_n8085), .ZN(MEM_stage_inst_dmem_n8150) );
NOR2_X1 MEM_stage_inst_dmem_U8200 ( .A1(MEM_stage_inst_dmem_n8084), .A2(MEM_stage_inst_dmem_n8083), .ZN(MEM_stage_inst_dmem_n8085) );
NAND2_X1 MEM_stage_inst_dmem_U8199 ( .A1(MEM_stage_inst_dmem_n8082), .A2(MEM_stage_inst_dmem_n8081), .ZN(MEM_stage_inst_dmem_n8083) );
NOR2_X1 MEM_stage_inst_dmem_U8198 ( .A1(MEM_stage_inst_dmem_n8080), .A2(MEM_stage_inst_dmem_n8079), .ZN(MEM_stage_inst_dmem_n8081) );
NAND2_X1 MEM_stage_inst_dmem_U8197 ( .A1(MEM_stage_inst_dmem_n8078), .A2(MEM_stage_inst_dmem_n8077), .ZN(MEM_stage_inst_dmem_n8079) );
NAND2_X1 MEM_stage_inst_dmem_U8196 ( .A1(MEM_stage_inst_dmem_ram_1743), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n8077) );
NAND2_X1 MEM_stage_inst_dmem_U8195 ( .A1(MEM_stage_inst_dmem_ram_1295), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n8078) );
NAND2_X1 MEM_stage_inst_dmem_U8194 ( .A1(MEM_stage_inst_dmem_n8076), .A2(MEM_stage_inst_dmem_n8075), .ZN(MEM_stage_inst_dmem_n8080) );
NAND2_X1 MEM_stage_inst_dmem_U8193 ( .A1(MEM_stage_inst_dmem_ram_1231), .A2(MEM_stage_inst_dmem_n36), .ZN(MEM_stage_inst_dmem_n8075) );
NAND2_X1 MEM_stage_inst_dmem_U8192 ( .A1(MEM_stage_inst_dmem_ram_1439), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n8076) );
NOR2_X1 MEM_stage_inst_dmem_U8191 ( .A1(MEM_stage_inst_dmem_n8074), .A2(MEM_stage_inst_dmem_n8073), .ZN(MEM_stage_inst_dmem_n8082) );
NAND2_X1 MEM_stage_inst_dmem_U8190 ( .A1(MEM_stage_inst_dmem_n8072), .A2(MEM_stage_inst_dmem_n8071), .ZN(MEM_stage_inst_dmem_n8073) );
NAND2_X1 MEM_stage_inst_dmem_U8189 ( .A1(MEM_stage_inst_dmem_n39), .A2(MEM_stage_inst_dmem_ram_1279), .ZN(MEM_stage_inst_dmem_n8071) );
NAND2_X1 MEM_stage_inst_dmem_U8188 ( .A1(MEM_stage_inst_dmem_n42), .A2(MEM_stage_inst_dmem_ram_1999), .ZN(MEM_stage_inst_dmem_n8072) );
NAND2_X1 MEM_stage_inst_dmem_U8187 ( .A1(MEM_stage_inst_dmem_n8070), .A2(MEM_stage_inst_dmem_n8069), .ZN(MEM_stage_inst_dmem_n8074) );
NAND2_X1 MEM_stage_inst_dmem_U8186 ( .A1(MEM_stage_inst_dmem_ram_2031), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n8069) );
NAND2_X1 MEM_stage_inst_dmem_U8185 ( .A1(MEM_stage_inst_dmem_ram_1567), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n8070) );
NAND2_X1 MEM_stage_inst_dmem_U8184 ( .A1(MEM_stage_inst_dmem_n8068), .A2(MEM_stage_inst_dmem_n8067), .ZN(MEM_stage_inst_dmem_n8084) );
NOR2_X1 MEM_stage_inst_dmem_U8183 ( .A1(MEM_stage_inst_dmem_n8066), .A2(MEM_stage_inst_dmem_n8065), .ZN(MEM_stage_inst_dmem_n8067) );
NAND2_X1 MEM_stage_inst_dmem_U8182 ( .A1(MEM_stage_inst_dmem_n8064), .A2(MEM_stage_inst_dmem_n8063), .ZN(MEM_stage_inst_dmem_n8065) );
NAND2_X1 MEM_stage_inst_dmem_U8181 ( .A1(MEM_stage_inst_dmem_ram_1919), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n8063) );
NAND2_X1 MEM_stage_inst_dmem_U8180 ( .A1(MEM_stage_inst_dmem_ram_1983), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n8064) );
NAND2_X1 MEM_stage_inst_dmem_U8179 ( .A1(MEM_stage_inst_dmem_n8062), .A2(MEM_stage_inst_dmem_n8061), .ZN(MEM_stage_inst_dmem_n8066) );
NAND2_X1 MEM_stage_inst_dmem_U8178 ( .A1(MEM_stage_inst_dmem_ram_1839), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n8061) );
NAND2_X1 MEM_stage_inst_dmem_U8177 ( .A1(MEM_stage_inst_dmem_ram_1711), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n8062) );
NOR2_X1 MEM_stage_inst_dmem_U8176 ( .A1(MEM_stage_inst_dmem_n8060), .A2(MEM_stage_inst_dmem_n8059), .ZN(MEM_stage_inst_dmem_n8068) );
NAND2_X1 MEM_stage_inst_dmem_U8175 ( .A1(MEM_stage_inst_dmem_n8058), .A2(MEM_stage_inst_dmem_n8057), .ZN(MEM_stage_inst_dmem_n8059) );
NAND2_X1 MEM_stage_inst_dmem_U8174 ( .A1(MEM_stage_inst_dmem_ram_1503), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n8057) );
NAND2_X1 MEM_stage_inst_dmem_U8173 ( .A1(MEM_stage_inst_dmem_ram_1551), .A2(MEM_stage_inst_dmem_n71), .ZN(MEM_stage_inst_dmem_n8058) );
NAND2_X1 MEM_stage_inst_dmem_U8172 ( .A1(MEM_stage_inst_dmem_n8056), .A2(MEM_stage_inst_dmem_n8055), .ZN(MEM_stage_inst_dmem_n8060) );
NAND2_X1 MEM_stage_inst_dmem_U8171 ( .A1(MEM_stage_inst_dmem_n19), .A2(MEM_stage_inst_dmem_ram_1519), .ZN(MEM_stage_inst_dmem_n8055) );
NAND2_X1 MEM_stage_inst_dmem_U8170 ( .A1(MEM_stage_inst_dmem_n22), .A2(MEM_stage_inst_dmem_ram_1775), .ZN(MEM_stage_inst_dmem_n8056) );
NOR2_X1 MEM_stage_inst_dmem_U8169 ( .A1(MEM_stage_inst_dmem_n8054), .A2(MEM_stage_inst_dmem_n8053), .ZN(MEM_stage_inst_dmem_n8086) );
NAND2_X1 MEM_stage_inst_dmem_U8168 ( .A1(MEM_stage_inst_dmem_n8052), .A2(MEM_stage_inst_dmem_n8051), .ZN(MEM_stage_inst_dmem_n8053) );
NOR2_X1 MEM_stage_inst_dmem_U8167 ( .A1(MEM_stage_inst_dmem_n8050), .A2(MEM_stage_inst_dmem_n8049), .ZN(MEM_stage_inst_dmem_n8051) );
NAND2_X1 MEM_stage_inst_dmem_U8166 ( .A1(MEM_stage_inst_dmem_n8048), .A2(MEM_stage_inst_dmem_n8047), .ZN(MEM_stage_inst_dmem_n8049) );
NAND2_X1 MEM_stage_inst_dmem_U8165 ( .A1(MEM_stage_inst_dmem_ram_1391), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n8047) );
NAND2_X1 MEM_stage_inst_dmem_U8164 ( .A1(MEM_stage_inst_dmem_ram_1247), .A2(MEM_stage_inst_dmem_n51), .ZN(MEM_stage_inst_dmem_n8048) );
NAND2_X1 MEM_stage_inst_dmem_U8163 ( .A1(MEM_stage_inst_dmem_n8046), .A2(MEM_stage_inst_dmem_n8045), .ZN(MEM_stage_inst_dmem_n8050) );
NAND2_X1 MEM_stage_inst_dmem_U8162 ( .A1(MEM_stage_inst_dmem_n46), .A2(MEM_stage_inst_dmem_ram_1855), .ZN(MEM_stage_inst_dmem_n8045) );
NAND2_X1 MEM_stage_inst_dmem_U8161 ( .A1(MEM_stage_inst_dmem_n50), .A2(MEM_stage_inst_dmem_ram_1727), .ZN(MEM_stage_inst_dmem_n8046) );
NOR2_X1 MEM_stage_inst_dmem_U8160 ( .A1(MEM_stage_inst_dmem_n8044), .A2(MEM_stage_inst_dmem_n8043), .ZN(MEM_stage_inst_dmem_n8052) );
NAND2_X1 MEM_stage_inst_dmem_U8159 ( .A1(MEM_stage_inst_dmem_n8042), .A2(MEM_stage_inst_dmem_n8041), .ZN(MEM_stage_inst_dmem_n8043) );
NAND2_X1 MEM_stage_inst_dmem_U8158 ( .A1(MEM_stage_inst_dmem_n30), .A2(MEM_stage_inst_dmem_ram_1647), .ZN(MEM_stage_inst_dmem_n8041) );
NAND2_X1 MEM_stage_inst_dmem_U8157 ( .A1(MEM_stage_inst_dmem_n74), .A2(MEM_stage_inst_dmem_ram_1583), .ZN(MEM_stage_inst_dmem_n8042) );
NAND2_X1 MEM_stage_inst_dmem_U8156 ( .A1(MEM_stage_inst_dmem_n8040), .A2(MEM_stage_inst_dmem_n8039), .ZN(MEM_stage_inst_dmem_n8044) );
NAND2_X1 MEM_stage_inst_dmem_U8155 ( .A1(MEM_stage_inst_dmem_ram_1679), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n8039) );
NAND2_X1 MEM_stage_inst_dmem_U8154 ( .A1(MEM_stage_inst_dmem_ram_1631), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n8040) );
NAND2_X1 MEM_stage_inst_dmem_U8153 ( .A1(MEM_stage_inst_dmem_n8038), .A2(MEM_stage_inst_dmem_n8037), .ZN(MEM_stage_inst_dmem_n8054) );
NOR2_X1 MEM_stage_inst_dmem_U8152 ( .A1(MEM_stage_inst_dmem_n8036), .A2(MEM_stage_inst_dmem_n8035), .ZN(MEM_stage_inst_dmem_n8037) );
NAND2_X1 MEM_stage_inst_dmem_U8151 ( .A1(MEM_stage_inst_dmem_n8034), .A2(MEM_stage_inst_dmem_n8033), .ZN(MEM_stage_inst_dmem_n8035) );
NAND2_X1 MEM_stage_inst_dmem_U8150 ( .A1(MEM_stage_inst_dmem_ram_1887), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n8033) );
NAND2_X1 MEM_stage_inst_dmem_U8149 ( .A1(MEM_stage_inst_dmem_ram_1135), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n8034) );
NAND2_X1 MEM_stage_inst_dmem_U8148 ( .A1(MEM_stage_inst_dmem_n8032), .A2(MEM_stage_inst_dmem_n8031), .ZN(MEM_stage_inst_dmem_n8036) );
NAND2_X1 MEM_stage_inst_dmem_U8147 ( .A1(MEM_stage_inst_dmem_n54), .A2(MEM_stage_inst_dmem_ram_1343), .ZN(MEM_stage_inst_dmem_n8031) );
NAND2_X1 MEM_stage_inst_dmem_U8146 ( .A1(MEM_stage_inst_dmem_n66), .A2(MEM_stage_inst_dmem_ram_1359), .ZN(MEM_stage_inst_dmem_n8032) );
NOR2_X1 MEM_stage_inst_dmem_U8145 ( .A1(MEM_stage_inst_dmem_n8030), .A2(MEM_stage_inst_dmem_n8029), .ZN(MEM_stage_inst_dmem_n8038) );
NAND2_X1 MEM_stage_inst_dmem_U8144 ( .A1(MEM_stage_inst_dmem_n8028), .A2(MEM_stage_inst_dmem_n8027), .ZN(MEM_stage_inst_dmem_n8029) );
NAND2_X1 MEM_stage_inst_dmem_U8143 ( .A1(MEM_stage_inst_dmem_ram_1103), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n8027) );
NAND2_X1 MEM_stage_inst_dmem_U8142 ( .A1(MEM_stage_inst_dmem_ram_1167), .A2(MEM_stage_inst_dmem_n61), .ZN(MEM_stage_inst_dmem_n8028) );
NAND2_X1 MEM_stage_inst_dmem_U8141 ( .A1(MEM_stage_inst_dmem_n8026), .A2(MEM_stage_inst_dmem_n8025), .ZN(MEM_stage_inst_dmem_n8030) );
NAND2_X1 MEM_stage_inst_dmem_U8140 ( .A1(MEM_stage_inst_dmem_n76), .A2(MEM_stage_inst_dmem_ram_1967), .ZN(MEM_stage_inst_dmem_n8025) );
NAND2_X1 MEM_stage_inst_dmem_U8139 ( .A1(MEM_stage_inst_dmem_n33), .A2(MEM_stage_inst_dmem_ram_1407), .ZN(MEM_stage_inst_dmem_n8026) );
NAND2_X1 MEM_stage_inst_dmem_U8138 ( .A1(MEM_stage_inst_dmem_n8024), .A2(MEM_stage_inst_dmem_n8023), .ZN(MEM_stage_inst_mem_read_data_14) );
NOR2_X1 MEM_stage_inst_dmem_U8137 ( .A1(MEM_stage_inst_dmem_n8022), .A2(MEM_stage_inst_dmem_n8021), .ZN(MEM_stage_inst_dmem_n8023) );
NOR2_X1 MEM_stage_inst_dmem_U8136 ( .A1(MEM_stage_inst_dmem_n8020), .A2(MEM_stage_inst_dmem_n8286), .ZN(MEM_stage_inst_dmem_n8021) );
NOR2_X1 MEM_stage_inst_dmem_U8135 ( .A1(MEM_stage_inst_dmem_n8019), .A2(MEM_stage_inst_dmem_n8018), .ZN(MEM_stage_inst_dmem_n8020) );
NAND2_X1 MEM_stage_inst_dmem_U8134 ( .A1(MEM_stage_inst_dmem_n8017), .A2(MEM_stage_inst_dmem_n8016), .ZN(MEM_stage_inst_dmem_n8018) );
NOR2_X1 MEM_stage_inst_dmem_U8133 ( .A1(MEM_stage_inst_dmem_n8015), .A2(MEM_stage_inst_dmem_n8014), .ZN(MEM_stage_inst_dmem_n8016) );
NAND2_X1 MEM_stage_inst_dmem_U8132 ( .A1(MEM_stage_inst_dmem_n8013), .A2(MEM_stage_inst_dmem_n8012), .ZN(MEM_stage_inst_dmem_n8014) );
NOR2_X1 MEM_stage_inst_dmem_U8131 ( .A1(MEM_stage_inst_dmem_n8011), .A2(MEM_stage_inst_dmem_n8010), .ZN(MEM_stage_inst_dmem_n8012) );
NAND2_X1 MEM_stage_inst_dmem_U8130 ( .A1(MEM_stage_inst_dmem_n8009), .A2(MEM_stage_inst_dmem_n8008), .ZN(MEM_stage_inst_dmem_n8010) );
NAND2_X1 MEM_stage_inst_dmem_U8129 ( .A1(MEM_stage_inst_dmem_ram_3006), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n8008) );
NAND2_X1 MEM_stage_inst_dmem_U8128 ( .A1(MEM_stage_inst_dmem_ram_2094), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n8009) );
NAND2_X1 MEM_stage_inst_dmem_U8127 ( .A1(MEM_stage_inst_dmem_n8007), .A2(MEM_stage_inst_dmem_n8006), .ZN(MEM_stage_inst_dmem_n8011) );
NAND2_X1 MEM_stage_inst_dmem_U8126 ( .A1(MEM_stage_inst_dmem_ram_2878), .A2(MEM_stage_inst_dmem_n8005), .ZN(MEM_stage_inst_dmem_n8006) );
NAND2_X1 MEM_stage_inst_dmem_U8125 ( .A1(MEM_stage_inst_dmem_ram_2750), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n8007) );
NOR2_X1 MEM_stage_inst_dmem_U8124 ( .A1(MEM_stage_inst_dmem_n8004), .A2(MEM_stage_inst_dmem_n8003), .ZN(MEM_stage_inst_dmem_n8013) );
NAND2_X1 MEM_stage_inst_dmem_U8123 ( .A1(MEM_stage_inst_dmem_n8002), .A2(MEM_stage_inst_dmem_n8001), .ZN(MEM_stage_inst_dmem_n8003) );
NAND2_X1 MEM_stage_inst_dmem_U8122 ( .A1(MEM_stage_inst_dmem_ram_2462), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n8001) );
NAND2_X1 MEM_stage_inst_dmem_U8121 ( .A1(MEM_stage_inst_dmem_ram_2222), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n8002) );
NAND2_X1 MEM_stage_inst_dmem_U8120 ( .A1(MEM_stage_inst_dmem_n8000), .A2(MEM_stage_inst_dmem_n7999), .ZN(MEM_stage_inst_dmem_n8004) );
NAND2_X1 MEM_stage_inst_dmem_U8119 ( .A1(MEM_stage_inst_dmem_ram_2958), .A2(MEM_stage_inst_dmem_n8193), .ZN(MEM_stage_inst_dmem_n7999) );
NAND2_X1 MEM_stage_inst_dmem_U8118 ( .A1(MEM_stage_inst_dmem_ram_2174), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n8000) );
NAND2_X1 MEM_stage_inst_dmem_U8117 ( .A1(MEM_stage_inst_dmem_n7998), .A2(MEM_stage_inst_dmem_n7997), .ZN(MEM_stage_inst_dmem_n8015) );
NOR2_X1 MEM_stage_inst_dmem_U8116 ( .A1(MEM_stage_inst_dmem_n7996), .A2(MEM_stage_inst_dmem_n7995), .ZN(MEM_stage_inst_dmem_n7997) );
NAND2_X1 MEM_stage_inst_dmem_U8115 ( .A1(MEM_stage_inst_dmem_n7994), .A2(MEM_stage_inst_dmem_n7993), .ZN(MEM_stage_inst_dmem_n7995) );
NAND2_X1 MEM_stage_inst_dmem_U8114 ( .A1(MEM_stage_inst_dmem_ram_2830), .A2(MEM_stage_inst_dmem_n7992), .ZN(MEM_stage_inst_dmem_n7993) );
NAND2_X1 MEM_stage_inst_dmem_U8113 ( .A1(MEM_stage_inst_dmem_ram_2686), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n7994) );
NAND2_X1 MEM_stage_inst_dmem_U8112 ( .A1(MEM_stage_inst_dmem_n7991), .A2(MEM_stage_inst_dmem_n7990), .ZN(MEM_stage_inst_dmem_n7996) );
NAND2_X1 MEM_stage_inst_dmem_U8111 ( .A1(MEM_stage_inst_dmem_ram_3022), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n7990) );
NAND2_X1 MEM_stage_inst_dmem_U8110 ( .A1(MEM_stage_inst_dmem_ram_2158), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n7991) );
NOR2_X1 MEM_stage_inst_dmem_U8109 ( .A1(MEM_stage_inst_dmem_n7989), .A2(MEM_stage_inst_dmem_n7988), .ZN(MEM_stage_inst_dmem_n7998) );
NAND2_X1 MEM_stage_inst_dmem_U8108 ( .A1(MEM_stage_inst_dmem_n7987), .A2(MEM_stage_inst_dmem_n7986), .ZN(MEM_stage_inst_dmem_n7988) );
NAND2_X1 MEM_stage_inst_dmem_U8107 ( .A1(MEM_stage_inst_dmem_ram_2846), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n7986) );
NAND2_X1 MEM_stage_inst_dmem_U8106 ( .A1(MEM_stage_inst_dmem_ram_2782), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n7987) );
NAND2_X1 MEM_stage_inst_dmem_U8105 ( .A1(MEM_stage_inst_dmem_n7985), .A2(MEM_stage_inst_dmem_n7984), .ZN(MEM_stage_inst_dmem_n7989) );
NAND2_X1 MEM_stage_inst_dmem_U8104 ( .A1(MEM_stage_inst_dmem_ram_2622), .A2(MEM_stage_inst_dmem_n8169), .ZN(MEM_stage_inst_dmem_n7984) );
NAND2_X1 MEM_stage_inst_dmem_U8103 ( .A1(MEM_stage_inst_dmem_ram_2350), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n7985) );
NOR2_X1 MEM_stage_inst_dmem_U8102 ( .A1(MEM_stage_inst_dmem_n7983), .A2(MEM_stage_inst_dmem_n7982), .ZN(MEM_stage_inst_dmem_n8017) );
NAND2_X1 MEM_stage_inst_dmem_U8101 ( .A1(MEM_stage_inst_dmem_n7981), .A2(MEM_stage_inst_dmem_n7980), .ZN(MEM_stage_inst_dmem_n7982) );
NOR2_X1 MEM_stage_inst_dmem_U8100 ( .A1(MEM_stage_inst_dmem_n7979), .A2(MEM_stage_inst_dmem_n7978), .ZN(MEM_stage_inst_dmem_n7980) );
NAND2_X1 MEM_stage_inst_dmem_U8099 ( .A1(MEM_stage_inst_dmem_n7977), .A2(MEM_stage_inst_dmem_n7976), .ZN(MEM_stage_inst_dmem_n7978) );
NAND2_X1 MEM_stage_inst_dmem_U8098 ( .A1(MEM_stage_inst_dmem_ram_2366), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n7976) );
NAND2_X1 MEM_stage_inst_dmem_U8097 ( .A1(MEM_stage_inst_dmem_ram_2398), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n7977) );
NAND2_X1 MEM_stage_inst_dmem_U8096 ( .A1(MEM_stage_inst_dmem_n7975), .A2(MEM_stage_inst_dmem_n7974), .ZN(MEM_stage_inst_dmem_n7979) );
NAND2_X1 MEM_stage_inst_dmem_U8095 ( .A1(MEM_stage_inst_dmem_ram_2414), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n7974) );
NAND2_X1 MEM_stage_inst_dmem_U8094 ( .A1(MEM_stage_inst_dmem_ram_2638), .A2(MEM_stage_inst_dmem_n7973), .ZN(MEM_stage_inst_dmem_n7975) );
NOR2_X1 MEM_stage_inst_dmem_U8093 ( .A1(MEM_stage_inst_dmem_n7972), .A2(MEM_stage_inst_dmem_n7971), .ZN(MEM_stage_inst_dmem_n7981) );
NAND2_X1 MEM_stage_inst_dmem_U8092 ( .A1(MEM_stage_inst_dmem_n7970), .A2(MEM_stage_inst_dmem_n7969), .ZN(MEM_stage_inst_dmem_n7971) );
NAND2_X1 MEM_stage_inst_dmem_U8091 ( .A1(MEM_stage_inst_dmem_ram_2478), .A2(MEM_stage_inst_dmem_n4772), .ZN(MEM_stage_inst_dmem_n7969) );
NAND2_X1 MEM_stage_inst_dmem_U8090 ( .A1(MEM_stage_inst_dmem_ram_2670), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n7970) );
NAND2_X1 MEM_stage_inst_dmem_U8089 ( .A1(MEM_stage_inst_dmem_n7968), .A2(MEM_stage_inst_dmem_n7967), .ZN(MEM_stage_inst_dmem_n7972) );
NAND2_X1 MEM_stage_inst_dmem_U8088 ( .A1(MEM_stage_inst_dmem_ram_2126), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n7967) );
NAND2_X1 MEM_stage_inst_dmem_U8087 ( .A1(MEM_stage_inst_dmem_ram_2798), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n7968) );
NAND2_X1 MEM_stage_inst_dmem_U8086 ( .A1(MEM_stage_inst_dmem_n7966), .A2(MEM_stage_inst_dmem_n7965), .ZN(MEM_stage_inst_dmem_n7983) );
NOR2_X1 MEM_stage_inst_dmem_U8085 ( .A1(MEM_stage_inst_dmem_n7964), .A2(MEM_stage_inst_dmem_n7963), .ZN(MEM_stage_inst_dmem_n7965) );
NAND2_X1 MEM_stage_inst_dmem_U8084 ( .A1(MEM_stage_inst_dmem_n7962), .A2(MEM_stage_inst_dmem_n7961), .ZN(MEM_stage_inst_dmem_n7963) );
NAND2_X1 MEM_stage_inst_dmem_U8083 ( .A1(MEM_stage_inst_dmem_ram_2702), .A2(MEM_stage_inst_dmem_n7960), .ZN(MEM_stage_inst_dmem_n7961) );
NAND2_X1 MEM_stage_inst_dmem_U8082 ( .A1(MEM_stage_inst_dmem_ram_2190), .A2(MEM_stage_inst_dmem_n8174), .ZN(MEM_stage_inst_dmem_n7962) );
NAND2_X1 MEM_stage_inst_dmem_U8081 ( .A1(MEM_stage_inst_dmem_n7959), .A2(MEM_stage_inst_dmem_n7958), .ZN(MEM_stage_inst_dmem_n7964) );
NAND2_X1 MEM_stage_inst_dmem_U8080 ( .A1(MEM_stage_inst_dmem_ram_2334), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n7958) );
NAND2_X1 MEM_stage_inst_dmem_U8079 ( .A1(MEM_stage_inst_dmem_ram_2430), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n7959) );
NOR2_X1 MEM_stage_inst_dmem_U8078 ( .A1(MEM_stage_inst_dmem_n7957), .A2(MEM_stage_inst_dmem_n7956), .ZN(MEM_stage_inst_dmem_n7966) );
NAND2_X1 MEM_stage_inst_dmem_U8077 ( .A1(MEM_stage_inst_dmem_n7955), .A2(MEM_stage_inst_dmem_n7954), .ZN(MEM_stage_inst_dmem_n7956) );
NAND2_X1 MEM_stage_inst_dmem_U8076 ( .A1(MEM_stage_inst_dmem_ram_2654), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n7954) );
NAND2_X1 MEM_stage_inst_dmem_U8075 ( .A1(MEM_stage_inst_dmem_ram_2062), .A2(MEM_stage_inst_dmem_n7953), .ZN(MEM_stage_inst_dmem_n7955) );
NAND2_X1 MEM_stage_inst_dmem_U8074 ( .A1(MEM_stage_inst_dmem_n7952), .A2(MEM_stage_inst_dmem_n7951), .ZN(MEM_stage_inst_dmem_n7957) );
NAND2_X1 MEM_stage_inst_dmem_U8073 ( .A1(MEM_stage_inst_dmem_ram_2910), .A2(MEM_stage_inst_dmem_n3141), .ZN(MEM_stage_inst_dmem_n7951) );
NAND2_X1 MEM_stage_inst_dmem_U8072 ( .A1(MEM_stage_inst_dmem_ram_3054), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n7952) );
NAND2_X1 MEM_stage_inst_dmem_U8071 ( .A1(MEM_stage_inst_dmem_n7950), .A2(MEM_stage_inst_dmem_n7949), .ZN(MEM_stage_inst_dmem_n8019) );
NOR2_X1 MEM_stage_inst_dmem_U8070 ( .A1(MEM_stage_inst_dmem_n7948), .A2(MEM_stage_inst_dmem_n7947), .ZN(MEM_stage_inst_dmem_n7949) );
NAND2_X1 MEM_stage_inst_dmem_U8069 ( .A1(MEM_stage_inst_dmem_n7946), .A2(MEM_stage_inst_dmem_n7945), .ZN(MEM_stage_inst_dmem_n7947) );
NOR2_X1 MEM_stage_inst_dmem_U8068 ( .A1(MEM_stage_inst_dmem_n7944), .A2(MEM_stage_inst_dmem_n7943), .ZN(MEM_stage_inst_dmem_n7945) );
NAND2_X1 MEM_stage_inst_dmem_U8067 ( .A1(MEM_stage_inst_dmem_n7942), .A2(MEM_stage_inst_dmem_n7941), .ZN(MEM_stage_inst_dmem_n7943) );
NAND2_X1 MEM_stage_inst_dmem_U8066 ( .A1(MEM_stage_inst_dmem_ram_2766), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n7941) );
NAND2_X1 MEM_stage_inst_dmem_U8065 ( .A1(MEM_stage_inst_dmem_ram_2862), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n7942) );
NAND2_X1 MEM_stage_inst_dmem_U8064 ( .A1(MEM_stage_inst_dmem_n7940), .A2(MEM_stage_inst_dmem_n7939), .ZN(MEM_stage_inst_dmem_n7944) );
NAND2_X1 MEM_stage_inst_dmem_U8063 ( .A1(MEM_stage_inst_dmem_ram_2142), .A2(MEM_stage_inst_dmem_n7938), .ZN(MEM_stage_inst_dmem_n7939) );
NAND2_X1 MEM_stage_inst_dmem_U8062 ( .A1(MEM_stage_inst_dmem_ram_2238), .A2(MEM_stage_inst_dmem_n7937), .ZN(MEM_stage_inst_dmem_n7940) );
NOR2_X1 MEM_stage_inst_dmem_U8061 ( .A1(MEM_stage_inst_dmem_n7936), .A2(MEM_stage_inst_dmem_n7935), .ZN(MEM_stage_inst_dmem_n7946) );
NAND2_X1 MEM_stage_inst_dmem_U8060 ( .A1(MEM_stage_inst_dmem_n7934), .A2(MEM_stage_inst_dmem_n7933), .ZN(MEM_stage_inst_dmem_n7935) );
NAND2_X1 MEM_stage_inst_dmem_U8059 ( .A1(MEM_stage_inst_dmem_ram_2558), .A2(MEM_stage_inst_dmem_n64), .ZN(MEM_stage_inst_dmem_n7933) );
NAND2_X1 MEM_stage_inst_dmem_U8058 ( .A1(MEM_stage_inst_dmem_ram_2606), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n7934) );
NAND2_X1 MEM_stage_inst_dmem_U8057 ( .A1(MEM_stage_inst_dmem_n7932), .A2(MEM_stage_inst_dmem_n7931), .ZN(MEM_stage_inst_dmem_n7936) );
NAND2_X1 MEM_stage_inst_dmem_U8056 ( .A1(MEM_stage_inst_dmem_ram_2974), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n7931) );
NAND2_X1 MEM_stage_inst_dmem_U8055 ( .A1(MEM_stage_inst_dmem_ram_2446), .A2(MEM_stage_inst_dmem_n7930), .ZN(MEM_stage_inst_dmem_n7932) );
NAND2_X1 MEM_stage_inst_dmem_U8054 ( .A1(MEM_stage_inst_dmem_n7929), .A2(MEM_stage_inst_dmem_n7928), .ZN(MEM_stage_inst_dmem_n7948) );
NOR2_X1 MEM_stage_inst_dmem_U8053 ( .A1(MEM_stage_inst_dmem_n7927), .A2(MEM_stage_inst_dmem_n7926), .ZN(MEM_stage_inst_dmem_n7928) );
NAND2_X1 MEM_stage_inst_dmem_U8052 ( .A1(MEM_stage_inst_dmem_n7925), .A2(MEM_stage_inst_dmem_n7924), .ZN(MEM_stage_inst_dmem_n7926) );
NAND2_X1 MEM_stage_inst_dmem_U8051 ( .A1(MEM_stage_inst_dmem_ram_2942), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n7924) );
NAND2_X1 MEM_stage_inst_dmem_U8050 ( .A1(MEM_stage_inst_dmem_ram_2926), .A2(MEM_stage_inst_dmem_n7923), .ZN(MEM_stage_inst_dmem_n7925) );
NAND2_X1 MEM_stage_inst_dmem_U8049 ( .A1(MEM_stage_inst_dmem_n7922), .A2(MEM_stage_inst_dmem_n7921), .ZN(MEM_stage_inst_dmem_n7927) );
NAND2_X1 MEM_stage_inst_dmem_U8048 ( .A1(MEM_stage_inst_dmem_ram_2270), .A2(MEM_stage_inst_dmem_n8206), .ZN(MEM_stage_inst_dmem_n7921) );
NAND2_X1 MEM_stage_inst_dmem_U8047 ( .A1(MEM_stage_inst_dmem_ram_3070), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n7922) );
NOR2_X1 MEM_stage_inst_dmem_U8046 ( .A1(MEM_stage_inst_dmem_n7920), .A2(MEM_stage_inst_dmem_n7919), .ZN(MEM_stage_inst_dmem_n7929) );
NAND2_X1 MEM_stage_inst_dmem_U8045 ( .A1(MEM_stage_inst_dmem_n7918), .A2(MEM_stage_inst_dmem_n7917), .ZN(MEM_stage_inst_dmem_n7919) );
NAND2_X1 MEM_stage_inst_dmem_U8044 ( .A1(MEM_stage_inst_dmem_ram_2814), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n7917) );
NAND2_X1 MEM_stage_inst_dmem_U8043 ( .A1(MEM_stage_inst_dmem_ram_2718), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n7918) );
NAND2_X1 MEM_stage_inst_dmem_U8042 ( .A1(MEM_stage_inst_dmem_n7916), .A2(MEM_stage_inst_dmem_n7915), .ZN(MEM_stage_inst_dmem_n7920) );
NAND2_X1 MEM_stage_inst_dmem_U8041 ( .A1(MEM_stage_inst_dmem_ram_2302), .A2(MEM_stage_inst_dmem_n7914), .ZN(MEM_stage_inst_dmem_n7915) );
NAND2_X1 MEM_stage_inst_dmem_U8040 ( .A1(MEM_stage_inst_dmem_ram_2510), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n7916) );
NOR2_X1 MEM_stage_inst_dmem_U8039 ( .A1(MEM_stage_inst_dmem_n7913), .A2(MEM_stage_inst_dmem_n7912), .ZN(MEM_stage_inst_dmem_n7950) );
NAND2_X1 MEM_stage_inst_dmem_U8038 ( .A1(MEM_stage_inst_dmem_n7911), .A2(MEM_stage_inst_dmem_n7910), .ZN(MEM_stage_inst_dmem_n7912) );
NOR2_X1 MEM_stage_inst_dmem_U8037 ( .A1(MEM_stage_inst_dmem_n7909), .A2(MEM_stage_inst_dmem_n7908), .ZN(MEM_stage_inst_dmem_n7910) );
NAND2_X1 MEM_stage_inst_dmem_U8036 ( .A1(MEM_stage_inst_dmem_n7907), .A2(MEM_stage_inst_dmem_n7906), .ZN(MEM_stage_inst_dmem_n7908) );
NAND2_X1 MEM_stage_inst_dmem_U8035 ( .A1(MEM_stage_inst_dmem_ram_2382), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n7906) );
NAND2_X1 MEM_stage_inst_dmem_U8034 ( .A1(MEM_stage_inst_dmem_ram_2542), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n7907) );
NAND2_X1 MEM_stage_inst_dmem_U8033 ( .A1(MEM_stage_inst_dmem_n7905), .A2(MEM_stage_inst_dmem_n7904), .ZN(MEM_stage_inst_dmem_n7909) );
NAND2_X1 MEM_stage_inst_dmem_U8032 ( .A1(MEM_stage_inst_dmem_ram_2526), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n7904) );
NAND2_X1 MEM_stage_inst_dmem_U8031 ( .A1(MEM_stage_inst_dmem_ram_2206), .A2(MEM_stage_inst_dmem_n7903), .ZN(MEM_stage_inst_dmem_n7905) );
NOR2_X1 MEM_stage_inst_dmem_U8030 ( .A1(MEM_stage_inst_dmem_n7902), .A2(MEM_stage_inst_dmem_n7901), .ZN(MEM_stage_inst_dmem_n7911) );
NAND2_X1 MEM_stage_inst_dmem_U8029 ( .A1(MEM_stage_inst_dmem_n7900), .A2(MEM_stage_inst_dmem_n7899), .ZN(MEM_stage_inst_dmem_n7901) );
NAND2_X1 MEM_stage_inst_dmem_U8028 ( .A1(MEM_stage_inst_dmem_ram_2286), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n7899) );
NAND2_X1 MEM_stage_inst_dmem_U8027 ( .A1(MEM_stage_inst_dmem_ram_2318), .A2(MEM_stage_inst_dmem_n7898), .ZN(MEM_stage_inst_dmem_n7900) );
NAND2_X1 MEM_stage_inst_dmem_U8026 ( .A1(MEM_stage_inst_dmem_n7897), .A2(MEM_stage_inst_dmem_n7896), .ZN(MEM_stage_inst_dmem_n7902) );
NAND2_X1 MEM_stage_inst_dmem_U8025 ( .A1(MEM_stage_inst_dmem_ram_3038), .A2(MEM_stage_inst_dmem_n7895), .ZN(MEM_stage_inst_dmem_n7896) );
NAND2_X1 MEM_stage_inst_dmem_U8024 ( .A1(MEM_stage_inst_dmem_ram_2574), .A2(MEM_stage_inst_dmem_n8225), .ZN(MEM_stage_inst_dmem_n7897) );
NAND2_X1 MEM_stage_inst_dmem_U8023 ( .A1(MEM_stage_inst_dmem_n7894), .A2(MEM_stage_inst_dmem_n7893), .ZN(MEM_stage_inst_dmem_n7913) );
NOR2_X1 MEM_stage_inst_dmem_U8022 ( .A1(MEM_stage_inst_dmem_n7892), .A2(MEM_stage_inst_dmem_n7891), .ZN(MEM_stage_inst_dmem_n7893) );
NAND2_X1 MEM_stage_inst_dmem_U8021 ( .A1(MEM_stage_inst_dmem_n7890), .A2(MEM_stage_inst_dmem_n7889), .ZN(MEM_stage_inst_dmem_n7891) );
NAND2_X1 MEM_stage_inst_dmem_U8020 ( .A1(MEM_stage_inst_dmem_ram_2494), .A2(MEM_stage_inst_dmem_n7888), .ZN(MEM_stage_inst_dmem_n7889) );
NAND2_X1 MEM_stage_inst_dmem_U8019 ( .A1(MEM_stage_inst_dmem_ram_2078), .A2(MEM_stage_inst_dmem_n7887), .ZN(MEM_stage_inst_dmem_n7890) );
NAND2_X1 MEM_stage_inst_dmem_U8018 ( .A1(MEM_stage_inst_dmem_n7886), .A2(MEM_stage_inst_dmem_n7885), .ZN(MEM_stage_inst_dmem_n7892) );
NAND2_X1 MEM_stage_inst_dmem_U8017 ( .A1(MEM_stage_inst_dmem_ram_2734), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n7885) );
NAND2_X1 MEM_stage_inst_dmem_U8016 ( .A1(MEM_stage_inst_dmem_ram_2590), .A2(MEM_stage_inst_dmem_n7884), .ZN(MEM_stage_inst_dmem_n7886) );
NOR2_X1 MEM_stage_inst_dmem_U8015 ( .A1(MEM_stage_inst_dmem_n7883), .A2(MEM_stage_inst_dmem_n7882), .ZN(MEM_stage_inst_dmem_n7894) );
NAND2_X1 MEM_stage_inst_dmem_U8014 ( .A1(MEM_stage_inst_dmem_n7881), .A2(MEM_stage_inst_dmem_n7880), .ZN(MEM_stage_inst_dmem_n7882) );
NAND2_X1 MEM_stage_inst_dmem_U8013 ( .A1(MEM_stage_inst_dmem_ram_2110), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n7880) );
NAND2_X1 MEM_stage_inst_dmem_U8012 ( .A1(MEM_stage_inst_dmem_ram_2990), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n7881) );
NAND2_X1 MEM_stage_inst_dmem_U8011 ( .A1(MEM_stage_inst_dmem_n7879), .A2(MEM_stage_inst_dmem_n7878), .ZN(MEM_stage_inst_dmem_n7883) );
NAND2_X1 MEM_stage_inst_dmem_U8010 ( .A1(MEM_stage_inst_dmem_ram_2254), .A2(MEM_stage_inst_dmem_n8256), .ZN(MEM_stage_inst_dmem_n7878) );
NAND2_X1 MEM_stage_inst_dmem_U8009 ( .A1(MEM_stage_inst_dmem_ram_2894), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n7879) );
NOR2_X1 MEM_stage_inst_dmem_U8008 ( .A1(MEM_stage_inst_dmem_n7877), .A2(MEM_stage_inst_dmem_n8551), .ZN(MEM_stage_inst_dmem_n8022) );
NOR2_X1 MEM_stage_inst_dmem_U8007 ( .A1(MEM_stage_inst_dmem_n7876), .A2(MEM_stage_inst_dmem_n7875), .ZN(MEM_stage_inst_dmem_n7877) );
NAND2_X1 MEM_stage_inst_dmem_U8006 ( .A1(MEM_stage_inst_dmem_n7874), .A2(MEM_stage_inst_dmem_n7873), .ZN(MEM_stage_inst_dmem_n7875) );
NOR2_X1 MEM_stage_inst_dmem_U8005 ( .A1(MEM_stage_inst_dmem_n7872), .A2(MEM_stage_inst_dmem_n7871), .ZN(MEM_stage_inst_dmem_n7873) );
NAND2_X1 MEM_stage_inst_dmem_U8004 ( .A1(MEM_stage_inst_dmem_n7870), .A2(MEM_stage_inst_dmem_n7869), .ZN(MEM_stage_inst_dmem_n7871) );
NOR2_X1 MEM_stage_inst_dmem_U8003 ( .A1(MEM_stage_inst_dmem_n7868), .A2(MEM_stage_inst_dmem_n7867), .ZN(MEM_stage_inst_dmem_n7869) );
NAND2_X1 MEM_stage_inst_dmem_U8002 ( .A1(MEM_stage_inst_dmem_n7866), .A2(MEM_stage_inst_dmem_n7865), .ZN(MEM_stage_inst_dmem_n7867) );
NAND2_X1 MEM_stage_inst_dmem_U8001 ( .A1(MEM_stage_inst_dmem_ram_254), .A2(MEM_stage_inst_dmem_n7914), .ZN(MEM_stage_inst_dmem_n7865) );
NAND2_X1 MEM_stage_inst_dmem_U8000 ( .A1(MEM_stage_inst_dmem_ram_542), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n7866) );
NAND2_X1 MEM_stage_inst_dmem_U7999 ( .A1(MEM_stage_inst_dmem_n7864), .A2(MEM_stage_inst_dmem_n7863), .ZN(MEM_stage_inst_dmem_n7868) );
NAND2_X1 MEM_stage_inst_dmem_U7998 ( .A1(MEM_stage_inst_dmem_ram_846), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n7863) );
NAND2_X1 MEM_stage_inst_dmem_U7997 ( .A1(MEM_stage_inst_dmem_ram_478), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n7864) );
NOR2_X1 MEM_stage_inst_dmem_U7996 ( .A1(MEM_stage_inst_dmem_n7862), .A2(MEM_stage_inst_dmem_n7861), .ZN(MEM_stage_inst_dmem_n7870) );
NAND2_X1 MEM_stage_inst_dmem_U7995 ( .A1(MEM_stage_inst_dmem_n7860), .A2(MEM_stage_inst_dmem_n7859), .ZN(MEM_stage_inst_dmem_n7861) );
NAND2_X1 MEM_stage_inst_dmem_U7994 ( .A1(MEM_stage_inst_dmem_ram_238), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n7859) );
NAND2_X1 MEM_stage_inst_dmem_U7993 ( .A1(MEM_stage_inst_dmem_ram_78), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n7860) );
NAND2_X1 MEM_stage_inst_dmem_U7992 ( .A1(MEM_stage_inst_dmem_n7858), .A2(MEM_stage_inst_dmem_n7857), .ZN(MEM_stage_inst_dmem_n7862) );
NAND2_X1 MEM_stage_inst_dmem_U7991 ( .A1(MEM_stage_inst_dmem_ram_1006), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n7857) );
NAND2_X1 MEM_stage_inst_dmem_U7990 ( .A1(MEM_stage_inst_dmem_ram_126), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n7858) );
NAND2_X1 MEM_stage_inst_dmem_U7989 ( .A1(MEM_stage_inst_dmem_n7856), .A2(MEM_stage_inst_dmem_n7855), .ZN(MEM_stage_inst_dmem_n7872) );
NOR2_X1 MEM_stage_inst_dmem_U7988 ( .A1(MEM_stage_inst_dmem_n7854), .A2(MEM_stage_inst_dmem_n7853), .ZN(MEM_stage_inst_dmem_n7855) );
NAND2_X1 MEM_stage_inst_dmem_U7987 ( .A1(MEM_stage_inst_dmem_n7852), .A2(MEM_stage_inst_dmem_n7851), .ZN(MEM_stage_inst_dmem_n7853) );
NAND2_X1 MEM_stage_inst_dmem_U7986 ( .A1(MEM_stage_inst_dmem_ram_878), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n7851) );
NAND2_X1 MEM_stage_inst_dmem_U7985 ( .A1(MEM_stage_inst_dmem_ram_926), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n7852) );
NAND2_X1 MEM_stage_inst_dmem_U7984 ( .A1(MEM_stage_inst_dmem_n7850), .A2(MEM_stage_inst_dmem_n7849), .ZN(MEM_stage_inst_dmem_n7854) );
NAND2_X1 MEM_stage_inst_dmem_U7983 ( .A1(MEM_stage_inst_dmem_ram_222), .A2(MEM_stage_inst_dmem_n51), .ZN(MEM_stage_inst_dmem_n7849) );
NAND2_X1 MEM_stage_inst_dmem_U7982 ( .A1(MEM_stage_inst_dmem_ram_734), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n7850) );
NOR2_X1 MEM_stage_inst_dmem_U7981 ( .A1(MEM_stage_inst_dmem_n7848), .A2(MEM_stage_inst_dmem_n7847), .ZN(MEM_stage_inst_dmem_n7856) );
NAND2_X1 MEM_stage_inst_dmem_U7980 ( .A1(MEM_stage_inst_dmem_n7846), .A2(MEM_stage_inst_dmem_n7845), .ZN(MEM_stage_inst_dmem_n7847) );
NAND2_X1 MEM_stage_inst_dmem_U7979 ( .A1(MEM_stage_inst_dmem_ram_142), .A2(MEM_stage_inst_dmem_n61), .ZN(MEM_stage_inst_dmem_n7845) );
NAND2_X1 MEM_stage_inst_dmem_U7978 ( .A1(MEM_stage_inst_dmem_ram_686), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n7846) );
NAND2_X1 MEM_stage_inst_dmem_U7977 ( .A1(MEM_stage_inst_dmem_n7844), .A2(MEM_stage_inst_dmem_n7843), .ZN(MEM_stage_inst_dmem_n7848) );
NAND2_X1 MEM_stage_inst_dmem_U7976 ( .A1(MEM_stage_inst_dmem_ram_830), .A2(MEM_stage_inst_dmem_n8005), .ZN(MEM_stage_inst_dmem_n7843) );
NAND2_X1 MEM_stage_inst_dmem_U7975 ( .A1(MEM_stage_inst_dmem_ram_750), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n7844) );
NOR2_X1 MEM_stage_inst_dmem_U7974 ( .A1(MEM_stage_inst_dmem_n7842), .A2(MEM_stage_inst_dmem_n7841), .ZN(MEM_stage_inst_dmem_n7874) );
NAND2_X1 MEM_stage_inst_dmem_U7973 ( .A1(MEM_stage_inst_dmem_n7840), .A2(MEM_stage_inst_dmem_n7839), .ZN(MEM_stage_inst_dmem_n7841) );
NOR2_X1 MEM_stage_inst_dmem_U7972 ( .A1(MEM_stage_inst_dmem_n7838), .A2(MEM_stage_inst_dmem_n7837), .ZN(MEM_stage_inst_dmem_n7839) );
NAND2_X1 MEM_stage_inst_dmem_U7971 ( .A1(MEM_stage_inst_dmem_n7836), .A2(MEM_stage_inst_dmem_n7835), .ZN(MEM_stage_inst_dmem_n7837) );
NAND2_X1 MEM_stage_inst_dmem_U7970 ( .A1(MEM_stage_inst_dmem_ram_94), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n7835) );
NAND2_X1 MEM_stage_inst_dmem_U7969 ( .A1(MEM_stage_inst_dmem_ram_270), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n7836) );
NAND2_X1 MEM_stage_inst_dmem_U7968 ( .A1(MEM_stage_inst_dmem_n7834), .A2(MEM_stage_inst_dmem_n7833), .ZN(MEM_stage_inst_dmem_n7838) );
NAND2_X1 MEM_stage_inst_dmem_U7967 ( .A1(MEM_stage_inst_dmem_ram_638), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n7833) );
NAND2_X1 MEM_stage_inst_dmem_U7966 ( .A1(MEM_stage_inst_dmem_ram_606), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n7834) );
NOR2_X1 MEM_stage_inst_dmem_U7965 ( .A1(MEM_stage_inst_dmem_n7832), .A2(MEM_stage_inst_dmem_n7831), .ZN(MEM_stage_inst_dmem_n7840) );
NAND2_X1 MEM_stage_inst_dmem_U7964 ( .A1(MEM_stage_inst_dmem_n7830), .A2(MEM_stage_inst_dmem_n7829), .ZN(MEM_stage_inst_dmem_n7831) );
NAND2_X1 MEM_stage_inst_dmem_U7963 ( .A1(MEM_stage_inst_dmem_ram_62), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n7829) );
NAND2_X1 MEM_stage_inst_dmem_U7962 ( .A1(MEM_stage_inst_dmem_ram_302), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n7830) );
NAND2_X1 MEM_stage_inst_dmem_U7961 ( .A1(MEM_stage_inst_dmem_n7828), .A2(MEM_stage_inst_dmem_n7827), .ZN(MEM_stage_inst_dmem_n7832) );
NAND2_X1 MEM_stage_inst_dmem_U7960 ( .A1(MEM_stage_inst_dmem_ram_494), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n7827) );
NAND2_X1 MEM_stage_inst_dmem_U7959 ( .A1(MEM_stage_inst_dmem_ram_110), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n7828) );
NAND2_X1 MEM_stage_inst_dmem_U7958 ( .A1(MEM_stage_inst_dmem_n7826), .A2(MEM_stage_inst_dmem_n7825), .ZN(MEM_stage_inst_dmem_n7842) );
NOR2_X1 MEM_stage_inst_dmem_U7957 ( .A1(MEM_stage_inst_dmem_n7824), .A2(MEM_stage_inst_dmem_n7823), .ZN(MEM_stage_inst_dmem_n7825) );
NAND2_X1 MEM_stage_inst_dmem_U7956 ( .A1(MEM_stage_inst_dmem_n7822), .A2(MEM_stage_inst_dmem_n7821), .ZN(MEM_stage_inst_dmem_n7823) );
NAND2_X1 MEM_stage_inst_dmem_U7955 ( .A1(MEM_stage_inst_dmem_ram_206), .A2(MEM_stage_inst_dmem_n36), .ZN(MEM_stage_inst_dmem_n7821) );
NAND2_X1 MEM_stage_inst_dmem_U7954 ( .A1(MEM_stage_inst_dmem_ram_14), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n7822) );
NAND2_X1 MEM_stage_inst_dmem_U7953 ( .A1(MEM_stage_inst_dmem_n7820), .A2(MEM_stage_inst_dmem_n7819), .ZN(MEM_stage_inst_dmem_n7824) );
NAND2_X1 MEM_stage_inst_dmem_U7952 ( .A1(MEM_stage_inst_dmem_ram_318), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n7819) );
NAND2_X1 MEM_stage_inst_dmem_U7951 ( .A1(MEM_stage_inst_dmem_ram_942), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n7820) );
NOR2_X1 MEM_stage_inst_dmem_U7950 ( .A1(MEM_stage_inst_dmem_n7818), .A2(MEM_stage_inst_dmem_n7817), .ZN(MEM_stage_inst_dmem_n7826) );
NAND2_X1 MEM_stage_inst_dmem_U7949 ( .A1(MEM_stage_inst_dmem_n7816), .A2(MEM_stage_inst_dmem_n7815), .ZN(MEM_stage_inst_dmem_n7817) );
NAND2_X1 MEM_stage_inst_dmem_U7948 ( .A1(MEM_stage_inst_dmem_ram_446), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n7815) );
NAND2_X1 MEM_stage_inst_dmem_U7947 ( .A1(MEM_stage_inst_dmem_ram_462), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n7816) );
NAND2_X1 MEM_stage_inst_dmem_U7946 ( .A1(MEM_stage_inst_dmem_n7814), .A2(MEM_stage_inst_dmem_n7813), .ZN(MEM_stage_inst_dmem_n7818) );
NAND2_X1 MEM_stage_inst_dmem_U7945 ( .A1(MEM_stage_inst_dmem_ram_910), .A2(MEM_stage_inst_dmem_n72), .ZN(MEM_stage_inst_dmem_n7813) );
NAND2_X1 MEM_stage_inst_dmem_U7944 ( .A1(MEM_stage_inst_dmem_ram_990), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n7814) );
NAND2_X1 MEM_stage_inst_dmem_U7943 ( .A1(MEM_stage_inst_dmem_n7812), .A2(MEM_stage_inst_dmem_n7811), .ZN(MEM_stage_inst_dmem_n7876) );
NOR2_X1 MEM_stage_inst_dmem_U7942 ( .A1(MEM_stage_inst_dmem_n7810), .A2(MEM_stage_inst_dmem_n7809), .ZN(MEM_stage_inst_dmem_n7811) );
NAND2_X1 MEM_stage_inst_dmem_U7941 ( .A1(MEM_stage_inst_dmem_n7808), .A2(MEM_stage_inst_dmem_n7807), .ZN(MEM_stage_inst_dmem_n7809) );
NOR2_X1 MEM_stage_inst_dmem_U7940 ( .A1(MEM_stage_inst_dmem_n7806), .A2(MEM_stage_inst_dmem_n7805), .ZN(MEM_stage_inst_dmem_n7807) );
NAND2_X1 MEM_stage_inst_dmem_U7939 ( .A1(MEM_stage_inst_dmem_n7804), .A2(MEM_stage_inst_dmem_n7803), .ZN(MEM_stage_inst_dmem_n7805) );
NAND2_X1 MEM_stage_inst_dmem_U7938 ( .A1(MEM_stage_inst_dmem_ram_46), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n7803) );
NAND2_X1 MEM_stage_inst_dmem_U7937 ( .A1(MEM_stage_inst_dmem_ram_158), .A2(MEM_stage_inst_dmem_n44), .ZN(MEM_stage_inst_dmem_n7804) );
NAND2_X1 MEM_stage_inst_dmem_U7936 ( .A1(MEM_stage_inst_dmem_n7802), .A2(MEM_stage_inst_dmem_n7801), .ZN(MEM_stage_inst_dmem_n7806) );
NAND2_X1 MEM_stage_inst_dmem_U7935 ( .A1(MEM_stage_inst_dmem_ram_334), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n7801) );
NAND2_X1 MEM_stage_inst_dmem_U7934 ( .A1(MEM_stage_inst_dmem_ram_414), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n7802) );
NOR2_X1 MEM_stage_inst_dmem_U7933 ( .A1(MEM_stage_inst_dmem_n7800), .A2(MEM_stage_inst_dmem_n7799), .ZN(MEM_stage_inst_dmem_n7808) );
NAND2_X1 MEM_stage_inst_dmem_U7932 ( .A1(MEM_stage_inst_dmem_n7798), .A2(MEM_stage_inst_dmem_n7797), .ZN(MEM_stage_inst_dmem_n7799) );
NAND2_X1 MEM_stage_inst_dmem_U7931 ( .A1(MEM_stage_inst_dmem_ram_894), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n7797) );
NAND2_X1 MEM_stage_inst_dmem_U7930 ( .A1(MEM_stage_inst_dmem_ram_766), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n7798) );
NAND2_X1 MEM_stage_inst_dmem_U7929 ( .A1(MEM_stage_inst_dmem_n7796), .A2(MEM_stage_inst_dmem_n7795), .ZN(MEM_stage_inst_dmem_n7800) );
NAND2_X1 MEM_stage_inst_dmem_U7928 ( .A1(MEM_stage_inst_dmem_ram_654), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n7795) );
NAND2_X1 MEM_stage_inst_dmem_U7927 ( .A1(MEM_stage_inst_dmem_ram_30), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n7796) );
NAND2_X1 MEM_stage_inst_dmem_U7926 ( .A1(MEM_stage_inst_dmem_n7794), .A2(MEM_stage_inst_dmem_n7793), .ZN(MEM_stage_inst_dmem_n7810) );
NOR2_X1 MEM_stage_inst_dmem_U7925 ( .A1(MEM_stage_inst_dmem_n7792), .A2(MEM_stage_inst_dmem_n7791), .ZN(MEM_stage_inst_dmem_n7793) );
NAND2_X1 MEM_stage_inst_dmem_U7924 ( .A1(MEM_stage_inst_dmem_n7790), .A2(MEM_stage_inst_dmem_n7789), .ZN(MEM_stage_inst_dmem_n7791) );
NAND2_X1 MEM_stage_inst_dmem_U7923 ( .A1(MEM_stage_inst_dmem_ram_430), .A2(MEM_stage_inst_dmem_n4772), .ZN(MEM_stage_inst_dmem_n7789) );
NAND2_X1 MEM_stage_inst_dmem_U7922 ( .A1(MEM_stage_inst_dmem_ram_174), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n7790) );
NAND2_X1 MEM_stage_inst_dmem_U7921 ( .A1(MEM_stage_inst_dmem_n7788), .A2(MEM_stage_inst_dmem_n7787), .ZN(MEM_stage_inst_dmem_n7792) );
NAND2_X1 MEM_stage_inst_dmem_U7920 ( .A1(MEM_stage_inst_dmem_ram_702), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n7787) );
NAND2_X1 MEM_stage_inst_dmem_U7919 ( .A1(MEM_stage_inst_dmem_ram_1022), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n7788) );
NOR2_X1 MEM_stage_inst_dmem_U7918 ( .A1(MEM_stage_inst_dmem_n7786), .A2(MEM_stage_inst_dmem_n7785), .ZN(MEM_stage_inst_dmem_n7794) );
NAND2_X1 MEM_stage_inst_dmem_U7917 ( .A1(MEM_stage_inst_dmem_n7784), .A2(MEM_stage_inst_dmem_n7783), .ZN(MEM_stage_inst_dmem_n7785) );
NAND2_X1 MEM_stage_inst_dmem_U7916 ( .A1(MEM_stage_inst_dmem_ram_958), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n7783) );
NAND2_X1 MEM_stage_inst_dmem_U7915 ( .A1(MEM_stage_inst_dmem_ram_590), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n7784) );
NAND2_X1 MEM_stage_inst_dmem_U7914 ( .A1(MEM_stage_inst_dmem_n7782), .A2(MEM_stage_inst_dmem_n7781), .ZN(MEM_stage_inst_dmem_n7786) );
NAND2_X1 MEM_stage_inst_dmem_U7913 ( .A1(MEM_stage_inst_dmem_ram_366), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n7781) );
NAND2_X1 MEM_stage_inst_dmem_U7912 ( .A1(MEM_stage_inst_dmem_ram_558), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n7782) );
NOR2_X1 MEM_stage_inst_dmem_U7911 ( .A1(MEM_stage_inst_dmem_n7780), .A2(MEM_stage_inst_dmem_n7779), .ZN(MEM_stage_inst_dmem_n7812) );
NAND2_X1 MEM_stage_inst_dmem_U7910 ( .A1(MEM_stage_inst_dmem_n7778), .A2(MEM_stage_inst_dmem_n7777), .ZN(MEM_stage_inst_dmem_n7779) );
NOR2_X1 MEM_stage_inst_dmem_U7909 ( .A1(MEM_stage_inst_dmem_n7776), .A2(MEM_stage_inst_dmem_n7775), .ZN(MEM_stage_inst_dmem_n7777) );
NAND2_X1 MEM_stage_inst_dmem_U7908 ( .A1(MEM_stage_inst_dmem_n7774), .A2(MEM_stage_inst_dmem_n7773), .ZN(MEM_stage_inst_dmem_n7775) );
NAND2_X1 MEM_stage_inst_dmem_U7907 ( .A1(MEM_stage_inst_dmem_ram_974), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n7773) );
NAND2_X1 MEM_stage_inst_dmem_U7906 ( .A1(MEM_stage_inst_dmem_ram_286), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n7774) );
NAND2_X1 MEM_stage_inst_dmem_U7905 ( .A1(MEM_stage_inst_dmem_n7772), .A2(MEM_stage_inst_dmem_n7771), .ZN(MEM_stage_inst_dmem_n7776) );
NAND2_X1 MEM_stage_inst_dmem_U7904 ( .A1(MEM_stage_inst_dmem_ram_190), .A2(MEM_stage_inst_dmem_n8434), .ZN(MEM_stage_inst_dmem_n7771) );
NAND2_X1 MEM_stage_inst_dmem_U7903 ( .A1(MEM_stage_inst_dmem_ram_670), .A2(MEM_stage_inst_dmem_n3076), .ZN(MEM_stage_inst_dmem_n7772) );
NOR2_X1 MEM_stage_inst_dmem_U7902 ( .A1(MEM_stage_inst_dmem_n7770), .A2(MEM_stage_inst_dmem_n7769), .ZN(MEM_stage_inst_dmem_n7778) );
NAND2_X1 MEM_stage_inst_dmem_U7901 ( .A1(MEM_stage_inst_dmem_n7768), .A2(MEM_stage_inst_dmem_n7767), .ZN(MEM_stage_inst_dmem_n7769) );
NAND2_X1 MEM_stage_inst_dmem_U7900 ( .A1(MEM_stage_inst_dmem_ram_782), .A2(MEM_stage_inst_dmem_n8472), .ZN(MEM_stage_inst_dmem_n7767) );
NAND2_X1 MEM_stage_inst_dmem_U7899 ( .A1(MEM_stage_inst_dmem_ram_574), .A2(MEM_stage_inst_dmem_n41), .ZN(MEM_stage_inst_dmem_n7768) );
NAND2_X1 MEM_stage_inst_dmem_U7898 ( .A1(MEM_stage_inst_dmem_n7766), .A2(MEM_stage_inst_dmem_n7765), .ZN(MEM_stage_inst_dmem_n7770) );
NAND2_X1 MEM_stage_inst_dmem_U7897 ( .A1(MEM_stage_inst_dmem_ram_622), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n7765) );
NAND2_X1 MEM_stage_inst_dmem_U7896 ( .A1(MEM_stage_inst_dmem_ram_526), .A2(MEM_stage_inst_dmem_n71), .ZN(MEM_stage_inst_dmem_n7766) );
NAND2_X1 MEM_stage_inst_dmem_U7895 ( .A1(MEM_stage_inst_dmem_n7764), .A2(MEM_stage_inst_dmem_n7763), .ZN(MEM_stage_inst_dmem_n7780) );
NOR2_X1 MEM_stage_inst_dmem_U7894 ( .A1(MEM_stage_inst_dmem_n7762), .A2(MEM_stage_inst_dmem_n7761), .ZN(MEM_stage_inst_dmem_n7763) );
NAND2_X1 MEM_stage_inst_dmem_U7893 ( .A1(MEM_stage_inst_dmem_n7760), .A2(MEM_stage_inst_dmem_n7759), .ZN(MEM_stage_inst_dmem_n7761) );
NAND2_X1 MEM_stage_inst_dmem_U7892 ( .A1(MEM_stage_inst_dmem_ram_718), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n7759) );
NAND2_X1 MEM_stage_inst_dmem_U7891 ( .A1(MEM_stage_inst_dmem_ram_382), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n7760) );
NAND2_X1 MEM_stage_inst_dmem_U7890 ( .A1(MEM_stage_inst_dmem_n7758), .A2(MEM_stage_inst_dmem_n7757), .ZN(MEM_stage_inst_dmem_n7762) );
NAND2_X1 MEM_stage_inst_dmem_U7889 ( .A1(MEM_stage_inst_dmem_ram_510), .A2(MEM_stage_inst_dmem_n8535), .ZN(MEM_stage_inst_dmem_n7757) );
NAND2_X1 MEM_stage_inst_dmem_U7888 ( .A1(MEM_stage_inst_dmem_ram_798), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n7758) );
NOR2_X1 MEM_stage_inst_dmem_U7887 ( .A1(MEM_stage_inst_dmem_n7756), .A2(MEM_stage_inst_dmem_n7755), .ZN(MEM_stage_inst_dmem_n7764) );
NAND2_X1 MEM_stage_inst_dmem_U7886 ( .A1(MEM_stage_inst_dmem_n7754), .A2(MEM_stage_inst_dmem_n7753), .ZN(MEM_stage_inst_dmem_n7755) );
NAND2_X1 MEM_stage_inst_dmem_U7885 ( .A1(MEM_stage_inst_dmem_ram_862), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n7753) );
NAND2_X1 MEM_stage_inst_dmem_U7884 ( .A1(MEM_stage_inst_dmem_ram_398), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n7754) );
NAND2_X1 MEM_stage_inst_dmem_U7883 ( .A1(MEM_stage_inst_dmem_n7752), .A2(MEM_stage_inst_dmem_n7751), .ZN(MEM_stage_inst_dmem_n7756) );
NAND2_X1 MEM_stage_inst_dmem_U7882 ( .A1(MEM_stage_inst_dmem_ram_814), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n7751) );
NAND2_X1 MEM_stage_inst_dmem_U7881 ( .A1(MEM_stage_inst_dmem_ram_350), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n7752) );
NOR2_X1 MEM_stage_inst_dmem_U7880 ( .A1(MEM_stage_inst_dmem_n7750), .A2(MEM_stage_inst_dmem_n7749), .ZN(MEM_stage_inst_dmem_n8024) );
NOR2_X1 MEM_stage_inst_dmem_U7879 ( .A1(MEM_stage_inst_dmem_n7748), .A2(MEM_stage_inst_dmem_n8152), .ZN(MEM_stage_inst_dmem_n7749) );
NOR2_X1 MEM_stage_inst_dmem_U7878 ( .A1(MEM_stage_inst_dmem_n7747), .A2(MEM_stage_inst_dmem_n7746), .ZN(MEM_stage_inst_dmem_n7748) );
NAND2_X1 MEM_stage_inst_dmem_U7877 ( .A1(MEM_stage_inst_dmem_n7745), .A2(MEM_stage_inst_dmem_n7744), .ZN(MEM_stage_inst_dmem_n7746) );
NOR2_X1 MEM_stage_inst_dmem_U7876 ( .A1(MEM_stage_inst_dmem_n7743), .A2(MEM_stage_inst_dmem_n7742), .ZN(MEM_stage_inst_dmem_n7744) );
NAND2_X1 MEM_stage_inst_dmem_U7875 ( .A1(MEM_stage_inst_dmem_n7741), .A2(MEM_stage_inst_dmem_n7740), .ZN(MEM_stage_inst_dmem_n7742) );
NOR2_X1 MEM_stage_inst_dmem_U7874 ( .A1(MEM_stage_inst_dmem_n7739), .A2(MEM_stage_inst_dmem_n7738), .ZN(MEM_stage_inst_dmem_n7740) );
NAND2_X1 MEM_stage_inst_dmem_U7873 ( .A1(MEM_stage_inst_dmem_n7737), .A2(MEM_stage_inst_dmem_n7736), .ZN(MEM_stage_inst_dmem_n7738) );
NAND2_X1 MEM_stage_inst_dmem_U7872 ( .A1(MEM_stage_inst_dmem_ram_1886), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n7736) );
NAND2_X1 MEM_stage_inst_dmem_U7871 ( .A1(MEM_stage_inst_dmem_ram_2014), .A2(MEM_stage_inst_dmem_n7895), .ZN(MEM_stage_inst_dmem_n7737) );
NAND2_X1 MEM_stage_inst_dmem_U7870 ( .A1(MEM_stage_inst_dmem_n7735), .A2(MEM_stage_inst_dmem_n7734), .ZN(MEM_stage_inst_dmem_n7739) );
NAND2_X1 MEM_stage_inst_dmem_U7869 ( .A1(MEM_stage_inst_dmem_ram_1342), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n7734) );
NAND2_X1 MEM_stage_inst_dmem_U7868 ( .A1(MEM_stage_inst_dmem_ram_1630), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n7735) );
NOR2_X1 MEM_stage_inst_dmem_U7867 ( .A1(MEM_stage_inst_dmem_n7733), .A2(MEM_stage_inst_dmem_n7732), .ZN(MEM_stage_inst_dmem_n7741) );
NAND2_X1 MEM_stage_inst_dmem_U7866 ( .A1(MEM_stage_inst_dmem_n7731), .A2(MEM_stage_inst_dmem_n7730), .ZN(MEM_stage_inst_dmem_n7732) );
NAND2_X1 MEM_stage_inst_dmem_U7865 ( .A1(MEM_stage_inst_dmem_ram_1918), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n7730) );
NAND2_X1 MEM_stage_inst_dmem_U7864 ( .A1(MEM_stage_inst_dmem_ram_1150), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n7731) );
NAND2_X1 MEM_stage_inst_dmem_U7863 ( .A1(MEM_stage_inst_dmem_n7729), .A2(MEM_stage_inst_dmem_n7728), .ZN(MEM_stage_inst_dmem_n7733) );
NAND2_X1 MEM_stage_inst_dmem_U7862 ( .A1(MEM_stage_inst_dmem_ram_1854), .A2(MEM_stage_inst_dmem_n8005), .ZN(MEM_stage_inst_dmem_n7728) );
NAND2_X1 MEM_stage_inst_dmem_U7861 ( .A1(MEM_stage_inst_dmem_ram_1662), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n7729) );
NAND2_X1 MEM_stage_inst_dmem_U7860 ( .A1(MEM_stage_inst_dmem_n7727), .A2(MEM_stage_inst_dmem_n7726), .ZN(MEM_stage_inst_dmem_n7743) );
NOR2_X1 MEM_stage_inst_dmem_U7859 ( .A1(MEM_stage_inst_dmem_n7725), .A2(MEM_stage_inst_dmem_n7724), .ZN(MEM_stage_inst_dmem_n7726) );
NAND2_X1 MEM_stage_inst_dmem_U7858 ( .A1(MEM_stage_inst_dmem_n7723), .A2(MEM_stage_inst_dmem_n7722), .ZN(MEM_stage_inst_dmem_n7724) );
NAND2_X1 MEM_stage_inst_dmem_U7857 ( .A1(MEM_stage_inst_dmem_ram_1502), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n7722) );
NAND2_X1 MEM_stage_inst_dmem_U7856 ( .A1(MEM_stage_inst_dmem_ram_1294), .A2(MEM_stage_inst_dmem_n7898), .ZN(MEM_stage_inst_dmem_n7723) );
NAND2_X1 MEM_stage_inst_dmem_U7855 ( .A1(MEM_stage_inst_dmem_n7721), .A2(MEM_stage_inst_dmem_n7720), .ZN(MEM_stage_inst_dmem_n7725) );
NAND2_X1 MEM_stage_inst_dmem_U7854 ( .A1(MEM_stage_inst_dmem_ram_1246), .A2(MEM_stage_inst_dmem_n51), .ZN(MEM_stage_inst_dmem_n7720) );
NAND2_X1 MEM_stage_inst_dmem_U7853 ( .A1(MEM_stage_inst_dmem_ram_1614), .A2(MEM_stage_inst_dmem_n7973), .ZN(MEM_stage_inst_dmem_n7721) );
NOR2_X1 MEM_stage_inst_dmem_U7852 ( .A1(MEM_stage_inst_dmem_n7719), .A2(MEM_stage_inst_dmem_n7718), .ZN(MEM_stage_inst_dmem_n7727) );
NAND2_X1 MEM_stage_inst_dmem_U7851 ( .A1(MEM_stage_inst_dmem_n7717), .A2(MEM_stage_inst_dmem_n7716), .ZN(MEM_stage_inst_dmem_n7718) );
NAND2_X1 MEM_stage_inst_dmem_U7850 ( .A1(MEM_stage_inst_dmem_ram_1230), .A2(MEM_stage_inst_dmem_n36), .ZN(MEM_stage_inst_dmem_n7716) );
NAND2_X1 MEM_stage_inst_dmem_U7849 ( .A1(MEM_stage_inst_dmem_ram_1982), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n7717) );
NAND2_X1 MEM_stage_inst_dmem_U7848 ( .A1(MEM_stage_inst_dmem_n7715), .A2(MEM_stage_inst_dmem_n7714), .ZN(MEM_stage_inst_dmem_n7719) );
NAND2_X1 MEM_stage_inst_dmem_U7847 ( .A1(MEM_stage_inst_dmem_ram_1486), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n7714) );
NAND2_X1 MEM_stage_inst_dmem_U7846 ( .A1(MEM_stage_inst_dmem_ram_1694), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n7715) );
NOR2_X1 MEM_stage_inst_dmem_U7845 ( .A1(MEM_stage_inst_dmem_n7713), .A2(MEM_stage_inst_dmem_n7712), .ZN(MEM_stage_inst_dmem_n7745) );
NAND2_X1 MEM_stage_inst_dmem_U7844 ( .A1(MEM_stage_inst_dmem_n7711), .A2(MEM_stage_inst_dmem_n7710), .ZN(MEM_stage_inst_dmem_n7712) );
NOR2_X1 MEM_stage_inst_dmem_U7843 ( .A1(MEM_stage_inst_dmem_n7709), .A2(MEM_stage_inst_dmem_n7708), .ZN(MEM_stage_inst_dmem_n7710) );
NAND2_X1 MEM_stage_inst_dmem_U7842 ( .A1(MEM_stage_inst_dmem_n7707), .A2(MEM_stage_inst_dmem_n7706), .ZN(MEM_stage_inst_dmem_n7708) );
NAND2_X1 MEM_stage_inst_dmem_U7841 ( .A1(MEM_stage_inst_dmem_ram_1726), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n7706) );
NAND2_X1 MEM_stage_inst_dmem_U7840 ( .A1(MEM_stage_inst_dmem_ram_1326), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n7707) );
NAND2_X1 MEM_stage_inst_dmem_U7839 ( .A1(MEM_stage_inst_dmem_n7705), .A2(MEM_stage_inst_dmem_n7704), .ZN(MEM_stage_inst_dmem_n7709) );
NAND2_X1 MEM_stage_inst_dmem_U7838 ( .A1(MEM_stage_inst_dmem_ram_1262), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n7704) );
NAND2_X1 MEM_stage_inst_dmem_U7837 ( .A1(MEM_stage_inst_dmem_ram_1118), .A2(MEM_stage_inst_dmem_n7938), .ZN(MEM_stage_inst_dmem_n7705) );
NOR2_X1 MEM_stage_inst_dmem_U7836 ( .A1(MEM_stage_inst_dmem_n7703), .A2(MEM_stage_inst_dmem_n7702), .ZN(MEM_stage_inst_dmem_n7711) );
NAND2_X1 MEM_stage_inst_dmem_U7835 ( .A1(MEM_stage_inst_dmem_n7701), .A2(MEM_stage_inst_dmem_n7700), .ZN(MEM_stage_inst_dmem_n7702) );
NAND2_X1 MEM_stage_inst_dmem_U7834 ( .A1(MEM_stage_inst_dmem_ram_1598), .A2(MEM_stage_inst_dmem_n41), .ZN(MEM_stage_inst_dmem_n7700) );
NAND2_X1 MEM_stage_inst_dmem_U7833 ( .A1(MEM_stage_inst_dmem_ram_1374), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n7701) );
NAND2_X1 MEM_stage_inst_dmem_U7832 ( .A1(MEM_stage_inst_dmem_n7699), .A2(MEM_stage_inst_dmem_n7698), .ZN(MEM_stage_inst_dmem_n7703) );
NAND2_X1 MEM_stage_inst_dmem_U7831 ( .A1(MEM_stage_inst_dmem_ram_1646), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n7698) );
NAND2_X1 MEM_stage_inst_dmem_U7830 ( .A1(MEM_stage_inst_dmem_ram_1966), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n7699) );
NAND2_X1 MEM_stage_inst_dmem_U7829 ( .A1(MEM_stage_inst_dmem_n7697), .A2(MEM_stage_inst_dmem_n7696), .ZN(MEM_stage_inst_dmem_n7713) );
NOR2_X1 MEM_stage_inst_dmem_U7828 ( .A1(MEM_stage_inst_dmem_n7695), .A2(MEM_stage_inst_dmem_n7694), .ZN(MEM_stage_inst_dmem_n7696) );
NAND2_X1 MEM_stage_inst_dmem_U7827 ( .A1(MEM_stage_inst_dmem_n7693), .A2(MEM_stage_inst_dmem_n7692), .ZN(MEM_stage_inst_dmem_n7694) );
NAND2_X1 MEM_stage_inst_dmem_U7826 ( .A1(MEM_stage_inst_dmem_ram_1038), .A2(MEM_stage_inst_dmem_n7953), .ZN(MEM_stage_inst_dmem_n7692) );
NAND2_X1 MEM_stage_inst_dmem_U7825 ( .A1(MEM_stage_inst_dmem_ram_1134), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n7693) );
NAND2_X1 MEM_stage_inst_dmem_U7824 ( .A1(MEM_stage_inst_dmem_n7691), .A2(MEM_stage_inst_dmem_n7690), .ZN(MEM_stage_inst_dmem_n7695) );
NAND2_X1 MEM_stage_inst_dmem_U7823 ( .A1(MEM_stage_inst_dmem_ram_1534), .A2(MEM_stage_inst_dmem_n64), .ZN(MEM_stage_inst_dmem_n7690) );
NAND2_X1 MEM_stage_inst_dmem_U7822 ( .A1(MEM_stage_inst_dmem_ram_1166), .A2(MEM_stage_inst_dmem_n61), .ZN(MEM_stage_inst_dmem_n7691) );
NOR2_X1 MEM_stage_inst_dmem_U7821 ( .A1(MEM_stage_inst_dmem_n7689), .A2(MEM_stage_inst_dmem_n7688), .ZN(MEM_stage_inst_dmem_n7697) );
NAND2_X1 MEM_stage_inst_dmem_U7820 ( .A1(MEM_stage_inst_dmem_n7687), .A2(MEM_stage_inst_dmem_n7686), .ZN(MEM_stage_inst_dmem_n7688) );
NAND2_X1 MEM_stage_inst_dmem_U7819 ( .A1(MEM_stage_inst_dmem_ram_1086), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n7686) );
NAND2_X1 MEM_stage_inst_dmem_U7818 ( .A1(MEM_stage_inst_dmem_ram_1422), .A2(MEM_stage_inst_dmem_n7930), .ZN(MEM_stage_inst_dmem_n7687) );
NAND2_X1 MEM_stage_inst_dmem_U7817 ( .A1(MEM_stage_inst_dmem_n7685), .A2(MEM_stage_inst_dmem_n7684), .ZN(MEM_stage_inst_dmem_n7689) );
NAND2_X1 MEM_stage_inst_dmem_U7816 ( .A1(MEM_stage_inst_dmem_ram_1790), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n7684) );
NAND2_X1 MEM_stage_inst_dmem_U7815 ( .A1(MEM_stage_inst_dmem_ram_1278), .A2(MEM_stage_inst_dmem_n7914), .ZN(MEM_stage_inst_dmem_n7685) );
NAND2_X1 MEM_stage_inst_dmem_U7814 ( .A1(MEM_stage_inst_dmem_n7683), .A2(MEM_stage_inst_dmem_n7682), .ZN(MEM_stage_inst_dmem_n7747) );
NOR2_X1 MEM_stage_inst_dmem_U7813 ( .A1(MEM_stage_inst_dmem_n7681), .A2(MEM_stage_inst_dmem_n7680), .ZN(MEM_stage_inst_dmem_n7682) );
NAND2_X1 MEM_stage_inst_dmem_U7812 ( .A1(MEM_stage_inst_dmem_n7679), .A2(MEM_stage_inst_dmem_n7678), .ZN(MEM_stage_inst_dmem_n7680) );
NOR2_X1 MEM_stage_inst_dmem_U7811 ( .A1(MEM_stage_inst_dmem_n7677), .A2(MEM_stage_inst_dmem_n7676), .ZN(MEM_stage_inst_dmem_n7678) );
NAND2_X1 MEM_stage_inst_dmem_U7810 ( .A1(MEM_stage_inst_dmem_n7675), .A2(MEM_stage_inst_dmem_n7674), .ZN(MEM_stage_inst_dmem_n7676) );
NAND2_X1 MEM_stage_inst_dmem_U7809 ( .A1(MEM_stage_inst_dmem_ram_1310), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n7674) );
NAND2_X1 MEM_stage_inst_dmem_U7808 ( .A1(MEM_stage_inst_dmem_ram_1838), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n7675) );
NAND2_X1 MEM_stage_inst_dmem_U7807 ( .A1(MEM_stage_inst_dmem_n7673), .A2(MEM_stage_inst_dmem_n7672), .ZN(MEM_stage_inst_dmem_n7677) );
NAND2_X1 MEM_stage_inst_dmem_U7806 ( .A1(MEM_stage_inst_dmem_ram_2046), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n7672) );
NAND2_X1 MEM_stage_inst_dmem_U7805 ( .A1(MEM_stage_inst_dmem_ram_1406), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n7673) );
NOR2_X1 MEM_stage_inst_dmem_U7804 ( .A1(MEM_stage_inst_dmem_n7671), .A2(MEM_stage_inst_dmem_n7670), .ZN(MEM_stage_inst_dmem_n7679) );
NAND2_X1 MEM_stage_inst_dmem_U7803 ( .A1(MEM_stage_inst_dmem_n7669), .A2(MEM_stage_inst_dmem_n7668), .ZN(MEM_stage_inst_dmem_n7670) );
NAND2_X1 MEM_stage_inst_dmem_U7802 ( .A1(MEM_stage_inst_dmem_ram_1214), .A2(MEM_stage_inst_dmem_n7937), .ZN(MEM_stage_inst_dmem_n7668) );
NAND2_X1 MEM_stage_inst_dmem_U7801 ( .A1(MEM_stage_inst_dmem_ram_1822), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n7669) );
NAND2_X1 MEM_stage_inst_dmem_U7800 ( .A1(MEM_stage_inst_dmem_n7667), .A2(MEM_stage_inst_dmem_n7666), .ZN(MEM_stage_inst_dmem_n7671) );
NAND2_X1 MEM_stage_inst_dmem_U7799 ( .A1(MEM_stage_inst_dmem_ram_1518), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n7666) );
NAND2_X1 MEM_stage_inst_dmem_U7798 ( .A1(MEM_stage_inst_dmem_ram_1582), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n7667) );
NAND2_X1 MEM_stage_inst_dmem_U7797 ( .A1(MEM_stage_inst_dmem_n7665), .A2(MEM_stage_inst_dmem_n7664), .ZN(MEM_stage_inst_dmem_n7681) );
NOR2_X1 MEM_stage_inst_dmem_U7796 ( .A1(MEM_stage_inst_dmem_n7663), .A2(MEM_stage_inst_dmem_n7662), .ZN(MEM_stage_inst_dmem_n7664) );
NAND2_X1 MEM_stage_inst_dmem_U7795 ( .A1(MEM_stage_inst_dmem_n7661), .A2(MEM_stage_inst_dmem_n7660), .ZN(MEM_stage_inst_dmem_n7662) );
NAND2_X1 MEM_stage_inst_dmem_U7794 ( .A1(MEM_stage_inst_dmem_ram_1742), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n7660) );
NAND2_X1 MEM_stage_inst_dmem_U7793 ( .A1(MEM_stage_inst_dmem_ram_1998), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n7661) );
NAND2_X1 MEM_stage_inst_dmem_U7792 ( .A1(MEM_stage_inst_dmem_n7659), .A2(MEM_stage_inst_dmem_n7658), .ZN(MEM_stage_inst_dmem_n7663) );
NAND2_X1 MEM_stage_inst_dmem_U7791 ( .A1(MEM_stage_inst_dmem_ram_1070), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n7658) );
NAND2_X1 MEM_stage_inst_dmem_U7790 ( .A1(MEM_stage_inst_dmem_ram_1774), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n7659) );
NOR2_X1 MEM_stage_inst_dmem_U7789 ( .A1(MEM_stage_inst_dmem_n7657), .A2(MEM_stage_inst_dmem_n7656), .ZN(MEM_stage_inst_dmem_n7665) );
NAND2_X1 MEM_stage_inst_dmem_U7788 ( .A1(MEM_stage_inst_dmem_n7655), .A2(MEM_stage_inst_dmem_n7654), .ZN(MEM_stage_inst_dmem_n7656) );
NAND2_X1 MEM_stage_inst_dmem_U7787 ( .A1(MEM_stage_inst_dmem_ram_1870), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n7654) );
NAND2_X1 MEM_stage_inst_dmem_U7786 ( .A1(MEM_stage_inst_dmem_ram_1678), .A2(MEM_stage_inst_dmem_n7960), .ZN(MEM_stage_inst_dmem_n7655) );
NAND2_X1 MEM_stage_inst_dmem_U7785 ( .A1(MEM_stage_inst_dmem_n7653), .A2(MEM_stage_inst_dmem_n7652), .ZN(MEM_stage_inst_dmem_n7657) );
NAND2_X1 MEM_stage_inst_dmem_U7784 ( .A1(MEM_stage_inst_dmem_ram_1902), .A2(MEM_stage_inst_dmem_n7923), .ZN(MEM_stage_inst_dmem_n7652) );
NAND2_X1 MEM_stage_inst_dmem_U7783 ( .A1(MEM_stage_inst_dmem_ram_1758), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n7653) );
NOR2_X1 MEM_stage_inst_dmem_U7782 ( .A1(MEM_stage_inst_dmem_n7651), .A2(MEM_stage_inst_dmem_n7650), .ZN(MEM_stage_inst_dmem_n7683) );
NAND2_X1 MEM_stage_inst_dmem_U7781 ( .A1(MEM_stage_inst_dmem_n7649), .A2(MEM_stage_inst_dmem_n7648), .ZN(MEM_stage_inst_dmem_n7650) );
NOR2_X1 MEM_stage_inst_dmem_U7780 ( .A1(MEM_stage_inst_dmem_n7647), .A2(MEM_stage_inst_dmem_n7646), .ZN(MEM_stage_inst_dmem_n7648) );
NAND2_X1 MEM_stage_inst_dmem_U7779 ( .A1(MEM_stage_inst_dmem_n7645), .A2(MEM_stage_inst_dmem_n7644), .ZN(MEM_stage_inst_dmem_n7646) );
NAND2_X1 MEM_stage_inst_dmem_U7778 ( .A1(MEM_stage_inst_dmem_ram_1710), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n7644) );
NAND2_X1 MEM_stage_inst_dmem_U7777 ( .A1(MEM_stage_inst_dmem_ram_1198), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n7645) );
NAND2_X1 MEM_stage_inst_dmem_U7776 ( .A1(MEM_stage_inst_dmem_n7643), .A2(MEM_stage_inst_dmem_n7642), .ZN(MEM_stage_inst_dmem_n7647) );
NAND2_X1 MEM_stage_inst_dmem_U7775 ( .A1(MEM_stage_inst_dmem_ram_1182), .A2(MEM_stage_inst_dmem_n7903), .ZN(MEM_stage_inst_dmem_n7642) );
NAND2_X1 MEM_stage_inst_dmem_U7774 ( .A1(MEM_stage_inst_dmem_ram_1550), .A2(MEM_stage_inst_dmem_n71), .ZN(MEM_stage_inst_dmem_n7643) );
NOR2_X1 MEM_stage_inst_dmem_U7773 ( .A1(MEM_stage_inst_dmem_n7641), .A2(MEM_stage_inst_dmem_n7640), .ZN(MEM_stage_inst_dmem_n7649) );
NAND2_X1 MEM_stage_inst_dmem_U7772 ( .A1(MEM_stage_inst_dmem_n7639), .A2(MEM_stage_inst_dmem_n7638), .ZN(MEM_stage_inst_dmem_n7640) );
NAND2_X1 MEM_stage_inst_dmem_U7771 ( .A1(MEM_stage_inst_dmem_ram_2030), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n7638) );
NAND2_X1 MEM_stage_inst_dmem_U7770 ( .A1(MEM_stage_inst_dmem_ram_1566), .A2(MEM_stage_inst_dmem_n7884), .ZN(MEM_stage_inst_dmem_n7639) );
NAND2_X1 MEM_stage_inst_dmem_U7769 ( .A1(MEM_stage_inst_dmem_n7637), .A2(MEM_stage_inst_dmem_n7636), .ZN(MEM_stage_inst_dmem_n7641) );
NAND2_X1 MEM_stage_inst_dmem_U7768 ( .A1(MEM_stage_inst_dmem_ram_1806), .A2(MEM_stage_inst_dmem_n7992), .ZN(MEM_stage_inst_dmem_n7636) );
NAND2_X1 MEM_stage_inst_dmem_U7767 ( .A1(MEM_stage_inst_dmem_ram_1390), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n7637) );
NAND2_X1 MEM_stage_inst_dmem_U7766 ( .A1(MEM_stage_inst_dmem_n7635), .A2(MEM_stage_inst_dmem_n7634), .ZN(MEM_stage_inst_dmem_n7651) );
NOR2_X1 MEM_stage_inst_dmem_U7765 ( .A1(MEM_stage_inst_dmem_n7633), .A2(MEM_stage_inst_dmem_n7632), .ZN(MEM_stage_inst_dmem_n7634) );
NAND2_X1 MEM_stage_inst_dmem_U7764 ( .A1(MEM_stage_inst_dmem_n7631), .A2(MEM_stage_inst_dmem_n7630), .ZN(MEM_stage_inst_dmem_n7632) );
NAND2_X1 MEM_stage_inst_dmem_U7763 ( .A1(MEM_stage_inst_dmem_ram_1438), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n7630) );
NAND2_X1 MEM_stage_inst_dmem_U7762 ( .A1(MEM_stage_inst_dmem_ram_1454), .A2(MEM_stage_inst_dmem_n4772), .ZN(MEM_stage_inst_dmem_n7631) );
NAND2_X1 MEM_stage_inst_dmem_U7761 ( .A1(MEM_stage_inst_dmem_n7629), .A2(MEM_stage_inst_dmem_n7628), .ZN(MEM_stage_inst_dmem_n7633) );
NAND2_X1 MEM_stage_inst_dmem_U7760 ( .A1(MEM_stage_inst_dmem_ram_1358), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n7628) );
NAND2_X1 MEM_stage_inst_dmem_U7759 ( .A1(MEM_stage_inst_dmem_ram_1054), .A2(MEM_stage_inst_dmem_n7887), .ZN(MEM_stage_inst_dmem_n7629) );
NOR2_X1 MEM_stage_inst_dmem_U7758 ( .A1(MEM_stage_inst_dmem_n7627), .A2(MEM_stage_inst_dmem_n7626), .ZN(MEM_stage_inst_dmem_n7635) );
NAND2_X1 MEM_stage_inst_dmem_U7757 ( .A1(MEM_stage_inst_dmem_n7625), .A2(MEM_stage_inst_dmem_n7624), .ZN(MEM_stage_inst_dmem_n7626) );
NAND2_X1 MEM_stage_inst_dmem_U7756 ( .A1(MEM_stage_inst_dmem_ram_1950), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n7624) );
NAND2_X1 MEM_stage_inst_dmem_U7755 ( .A1(MEM_stage_inst_dmem_ram_1934), .A2(MEM_stage_inst_dmem_n72), .ZN(MEM_stage_inst_dmem_n7625) );
NAND2_X1 MEM_stage_inst_dmem_U7754 ( .A1(MEM_stage_inst_dmem_n7623), .A2(MEM_stage_inst_dmem_n7622), .ZN(MEM_stage_inst_dmem_n7627) );
NAND2_X1 MEM_stage_inst_dmem_U7753 ( .A1(MEM_stage_inst_dmem_ram_1470), .A2(MEM_stage_inst_dmem_n7888), .ZN(MEM_stage_inst_dmem_n7622) );
NAND2_X1 MEM_stage_inst_dmem_U7752 ( .A1(MEM_stage_inst_dmem_ram_1102), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n7623) );
NOR2_X1 MEM_stage_inst_dmem_U7751 ( .A1(MEM_stage_inst_dmem_n7621), .A2(MEM_stage_inst_dmem_n8417), .ZN(MEM_stage_inst_dmem_n7750) );
NOR2_X1 MEM_stage_inst_dmem_U7750 ( .A1(MEM_stage_inst_dmem_n7620), .A2(MEM_stage_inst_dmem_n7619), .ZN(MEM_stage_inst_dmem_n7621) );
NAND2_X1 MEM_stage_inst_dmem_U7749 ( .A1(MEM_stage_inst_dmem_n7618), .A2(MEM_stage_inst_dmem_n7617), .ZN(MEM_stage_inst_dmem_n7619) );
NOR2_X1 MEM_stage_inst_dmem_U7748 ( .A1(MEM_stage_inst_dmem_n7616), .A2(MEM_stage_inst_dmem_n7615), .ZN(MEM_stage_inst_dmem_n7617) );
NAND2_X1 MEM_stage_inst_dmem_U7747 ( .A1(MEM_stage_inst_dmem_n7614), .A2(MEM_stage_inst_dmem_n7613), .ZN(MEM_stage_inst_dmem_n7615) );
NOR2_X1 MEM_stage_inst_dmem_U7746 ( .A1(MEM_stage_inst_dmem_n7612), .A2(MEM_stage_inst_dmem_n7611), .ZN(MEM_stage_inst_dmem_n7613) );
NAND2_X1 MEM_stage_inst_dmem_U7745 ( .A1(MEM_stage_inst_dmem_n7610), .A2(MEM_stage_inst_dmem_n7609), .ZN(MEM_stage_inst_dmem_n7611) );
NAND2_X1 MEM_stage_inst_dmem_U7744 ( .A1(MEM_stage_inst_dmem_ram_3982), .A2(MEM_stage_inst_dmem_n8193), .ZN(MEM_stage_inst_dmem_n7609) );
NAND2_X1 MEM_stage_inst_dmem_U7743 ( .A1(MEM_stage_inst_dmem_ram_3470), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n7610) );
NAND2_X1 MEM_stage_inst_dmem_U7742 ( .A1(MEM_stage_inst_dmem_n7608), .A2(MEM_stage_inst_dmem_n7607), .ZN(MEM_stage_inst_dmem_n7612) );
NAND2_X1 MEM_stage_inst_dmem_U7741 ( .A1(MEM_stage_inst_dmem_ram_3166), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n7607) );
NAND2_X1 MEM_stage_inst_dmem_U7740 ( .A1(MEM_stage_inst_dmem_ram_4094), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n7608) );
NOR2_X1 MEM_stage_inst_dmem_U7739 ( .A1(MEM_stage_inst_dmem_n7606), .A2(MEM_stage_inst_dmem_n7605), .ZN(MEM_stage_inst_dmem_n7614) );
NAND2_X1 MEM_stage_inst_dmem_U7738 ( .A1(MEM_stage_inst_dmem_n7604), .A2(MEM_stage_inst_dmem_n7603), .ZN(MEM_stage_inst_dmem_n7605) );
NAND2_X1 MEM_stage_inst_dmem_U7737 ( .A1(MEM_stage_inst_dmem_ram_3214), .A2(MEM_stage_inst_dmem_n8174), .ZN(MEM_stage_inst_dmem_n7603) );
NAND2_X1 MEM_stage_inst_dmem_U7736 ( .A1(MEM_stage_inst_dmem_ram_3294), .A2(MEM_stage_inst_dmem_n8206), .ZN(MEM_stage_inst_dmem_n7604) );
NAND2_X1 MEM_stage_inst_dmem_U7735 ( .A1(MEM_stage_inst_dmem_n7602), .A2(MEM_stage_inst_dmem_n7601), .ZN(MEM_stage_inst_dmem_n7606) );
NAND2_X1 MEM_stage_inst_dmem_U7734 ( .A1(MEM_stage_inst_dmem_ram_3998), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n7601) );
NAND2_X1 MEM_stage_inst_dmem_U7733 ( .A1(MEM_stage_inst_dmem_ram_4046), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n7602) );
NAND2_X1 MEM_stage_inst_dmem_U7732 ( .A1(MEM_stage_inst_dmem_n7600), .A2(MEM_stage_inst_dmem_n7599), .ZN(MEM_stage_inst_dmem_n7616) );
NOR2_X1 MEM_stage_inst_dmem_U7731 ( .A1(MEM_stage_inst_dmem_n7598), .A2(MEM_stage_inst_dmem_n7597), .ZN(MEM_stage_inst_dmem_n7599) );
NAND2_X1 MEM_stage_inst_dmem_U7730 ( .A1(MEM_stage_inst_dmem_n7596), .A2(MEM_stage_inst_dmem_n7595), .ZN(MEM_stage_inst_dmem_n7597) );
NAND2_X1 MEM_stage_inst_dmem_U7729 ( .A1(MEM_stage_inst_dmem_ram_3646), .A2(MEM_stage_inst_dmem_n8169), .ZN(MEM_stage_inst_dmem_n7595) );
NAND2_X1 MEM_stage_inst_dmem_U7728 ( .A1(MEM_stage_inst_dmem_ram_3614), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n7596) );
NAND2_X1 MEM_stage_inst_dmem_U7727 ( .A1(MEM_stage_inst_dmem_n7594), .A2(MEM_stage_inst_dmem_n7593), .ZN(MEM_stage_inst_dmem_n7598) );
NAND2_X1 MEM_stage_inst_dmem_U7726 ( .A1(MEM_stage_inst_dmem_ram_3310), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n7593) );
NAND2_X1 MEM_stage_inst_dmem_U7725 ( .A1(MEM_stage_inst_dmem_ram_3838), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n7594) );
NOR2_X1 MEM_stage_inst_dmem_U7724 ( .A1(MEM_stage_inst_dmem_n7592), .A2(MEM_stage_inst_dmem_n7591), .ZN(MEM_stage_inst_dmem_n7600) );
NAND2_X1 MEM_stage_inst_dmem_U7723 ( .A1(MEM_stage_inst_dmem_n7590), .A2(MEM_stage_inst_dmem_n7589), .ZN(MEM_stage_inst_dmem_n7591) );
NAND2_X1 MEM_stage_inst_dmem_U7722 ( .A1(MEM_stage_inst_dmem_ram_3774), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n7589) );
NAND2_X1 MEM_stage_inst_dmem_U7721 ( .A1(MEM_stage_inst_dmem_ram_3422), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n7590) );
NAND2_X1 MEM_stage_inst_dmem_U7720 ( .A1(MEM_stage_inst_dmem_n7588), .A2(MEM_stage_inst_dmem_n7587), .ZN(MEM_stage_inst_dmem_n7592) );
NAND2_X1 MEM_stage_inst_dmem_U7719 ( .A1(MEM_stage_inst_dmem_ram_3966), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n7587) );
NAND2_X1 MEM_stage_inst_dmem_U7718 ( .A1(MEM_stage_inst_dmem_ram_3374), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n7588) );
NOR2_X1 MEM_stage_inst_dmem_U7717 ( .A1(MEM_stage_inst_dmem_n7586), .A2(MEM_stage_inst_dmem_n7585), .ZN(MEM_stage_inst_dmem_n7618) );
NAND2_X1 MEM_stage_inst_dmem_U7716 ( .A1(MEM_stage_inst_dmem_n7584), .A2(MEM_stage_inst_dmem_n7583), .ZN(MEM_stage_inst_dmem_n7585) );
NOR2_X1 MEM_stage_inst_dmem_U7715 ( .A1(MEM_stage_inst_dmem_n7582), .A2(MEM_stage_inst_dmem_n7581), .ZN(MEM_stage_inst_dmem_n7583) );
NAND2_X1 MEM_stage_inst_dmem_U7714 ( .A1(MEM_stage_inst_dmem_n7580), .A2(MEM_stage_inst_dmem_n7579), .ZN(MEM_stage_inst_dmem_n7581) );
NAND2_X1 MEM_stage_inst_dmem_U7713 ( .A1(MEM_stage_inst_dmem_ram_3326), .A2(MEM_stage_inst_dmem_n7914), .ZN(MEM_stage_inst_dmem_n7579) );
NAND2_X1 MEM_stage_inst_dmem_U7712 ( .A1(MEM_stage_inst_dmem_ram_3534), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n7580) );
NAND2_X1 MEM_stage_inst_dmem_U7711 ( .A1(MEM_stage_inst_dmem_n7578), .A2(MEM_stage_inst_dmem_n7577), .ZN(MEM_stage_inst_dmem_n7582) );
NAND2_X1 MEM_stage_inst_dmem_U7710 ( .A1(MEM_stage_inst_dmem_ram_3438), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n7577) );
NAND2_X1 MEM_stage_inst_dmem_U7709 ( .A1(MEM_stage_inst_dmem_ram_3230), .A2(MEM_stage_inst_dmem_n44), .ZN(MEM_stage_inst_dmem_n7578) );
NOR2_X1 MEM_stage_inst_dmem_U7708 ( .A1(MEM_stage_inst_dmem_n7576), .A2(MEM_stage_inst_dmem_n7575), .ZN(MEM_stage_inst_dmem_n7584) );
NAND2_X1 MEM_stage_inst_dmem_U7707 ( .A1(MEM_stage_inst_dmem_n7574), .A2(MEM_stage_inst_dmem_n7573), .ZN(MEM_stage_inst_dmem_n7575) );
NAND2_X1 MEM_stage_inst_dmem_U7706 ( .A1(MEM_stage_inst_dmem_ram_3390), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n7573) );
NAND2_X1 MEM_stage_inst_dmem_U7705 ( .A1(MEM_stage_inst_dmem_ram_4030), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n7574) );
NAND2_X1 MEM_stage_inst_dmem_U7704 ( .A1(MEM_stage_inst_dmem_n7572), .A2(MEM_stage_inst_dmem_n7571), .ZN(MEM_stage_inst_dmem_n7576) );
NAND2_X1 MEM_stage_inst_dmem_U7703 ( .A1(MEM_stage_inst_dmem_ram_3934), .A2(MEM_stage_inst_dmem_n3141), .ZN(MEM_stage_inst_dmem_n7571) );
NAND2_X1 MEM_stage_inst_dmem_U7702 ( .A1(MEM_stage_inst_dmem_ram_3726), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n7572) );
NAND2_X1 MEM_stage_inst_dmem_U7701 ( .A1(MEM_stage_inst_dmem_n7570), .A2(MEM_stage_inst_dmem_n7569), .ZN(MEM_stage_inst_dmem_n7586) );
NOR2_X1 MEM_stage_inst_dmem_U7700 ( .A1(MEM_stage_inst_dmem_n7568), .A2(MEM_stage_inst_dmem_n7567), .ZN(MEM_stage_inst_dmem_n7569) );
NAND2_X1 MEM_stage_inst_dmem_U7699 ( .A1(MEM_stage_inst_dmem_n7566), .A2(MEM_stage_inst_dmem_n7565), .ZN(MEM_stage_inst_dmem_n7567) );
NAND2_X1 MEM_stage_inst_dmem_U7698 ( .A1(MEM_stage_inst_dmem_ram_3550), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n7565) );
NAND2_X1 MEM_stage_inst_dmem_U7697 ( .A1(MEM_stage_inst_dmem_ram_3822), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n7566) );
NAND2_X1 MEM_stage_inst_dmem_U7696 ( .A1(MEM_stage_inst_dmem_n7564), .A2(MEM_stage_inst_dmem_n7563), .ZN(MEM_stage_inst_dmem_n7568) );
NAND2_X1 MEM_stage_inst_dmem_U7695 ( .A1(MEM_stage_inst_dmem_ram_3198), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n7563) );
NAND2_X1 MEM_stage_inst_dmem_U7694 ( .A1(MEM_stage_inst_dmem_ram_3678), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n7564) );
NOR2_X1 MEM_stage_inst_dmem_U7693 ( .A1(MEM_stage_inst_dmem_n7562), .A2(MEM_stage_inst_dmem_n7561), .ZN(MEM_stage_inst_dmem_n7570) );
NAND2_X1 MEM_stage_inst_dmem_U7692 ( .A1(MEM_stage_inst_dmem_n7560), .A2(MEM_stage_inst_dmem_n7559), .ZN(MEM_stage_inst_dmem_n7561) );
NAND2_X1 MEM_stage_inst_dmem_U7691 ( .A1(MEM_stage_inst_dmem_ram_3758), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n7559) );
NAND2_X1 MEM_stage_inst_dmem_U7690 ( .A1(MEM_stage_inst_dmem_ram_3342), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n7560) );
NAND2_X1 MEM_stage_inst_dmem_U7689 ( .A1(MEM_stage_inst_dmem_n7558), .A2(MEM_stage_inst_dmem_n7557), .ZN(MEM_stage_inst_dmem_n7562) );
NAND2_X1 MEM_stage_inst_dmem_U7688 ( .A1(MEM_stage_inst_dmem_ram_3950), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n7557) );
NAND2_X1 MEM_stage_inst_dmem_U7687 ( .A1(MEM_stage_inst_dmem_ram_3086), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n7558) );
NAND2_X1 MEM_stage_inst_dmem_U7686 ( .A1(MEM_stage_inst_dmem_n7556), .A2(MEM_stage_inst_dmem_n7555), .ZN(MEM_stage_inst_dmem_n7620) );
NOR2_X1 MEM_stage_inst_dmem_U7685 ( .A1(MEM_stage_inst_dmem_n7554), .A2(MEM_stage_inst_dmem_n7553), .ZN(MEM_stage_inst_dmem_n7555) );
NAND2_X1 MEM_stage_inst_dmem_U7684 ( .A1(MEM_stage_inst_dmem_n7552), .A2(MEM_stage_inst_dmem_n7551), .ZN(MEM_stage_inst_dmem_n7553) );
NOR2_X1 MEM_stage_inst_dmem_U7683 ( .A1(MEM_stage_inst_dmem_n7550), .A2(MEM_stage_inst_dmem_n7549), .ZN(MEM_stage_inst_dmem_n7551) );
NAND2_X1 MEM_stage_inst_dmem_U7682 ( .A1(MEM_stage_inst_dmem_n7548), .A2(MEM_stage_inst_dmem_n7547), .ZN(MEM_stage_inst_dmem_n7549) );
NAND2_X1 MEM_stage_inst_dmem_U7681 ( .A1(MEM_stage_inst_dmem_ram_3710), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n7547) );
NAND2_X1 MEM_stage_inst_dmem_U7680 ( .A1(MEM_stage_inst_dmem_ram_3246), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n7548) );
NAND2_X1 MEM_stage_inst_dmem_U7679 ( .A1(MEM_stage_inst_dmem_n7546), .A2(MEM_stage_inst_dmem_n7545), .ZN(MEM_stage_inst_dmem_n7550) );
NAND2_X1 MEM_stage_inst_dmem_U7678 ( .A1(MEM_stage_inst_dmem_ram_4078), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n7545) );
NAND2_X1 MEM_stage_inst_dmem_U7677 ( .A1(MEM_stage_inst_dmem_ram_3262), .A2(MEM_stage_inst_dmem_n8434), .ZN(MEM_stage_inst_dmem_n7546) );
NOR2_X1 MEM_stage_inst_dmem_U7676 ( .A1(MEM_stage_inst_dmem_n7544), .A2(MEM_stage_inst_dmem_n7543), .ZN(MEM_stage_inst_dmem_n7552) );
NAND2_X1 MEM_stage_inst_dmem_U7675 ( .A1(MEM_stage_inst_dmem_n7542), .A2(MEM_stage_inst_dmem_n7541), .ZN(MEM_stage_inst_dmem_n7543) );
NAND2_X1 MEM_stage_inst_dmem_U7674 ( .A1(MEM_stage_inst_dmem_ram_3134), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n7541) );
NAND2_X1 MEM_stage_inst_dmem_U7673 ( .A1(MEM_stage_inst_dmem_ram_3566), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n7542) );
NAND2_X1 MEM_stage_inst_dmem_U7672 ( .A1(MEM_stage_inst_dmem_n7540), .A2(MEM_stage_inst_dmem_n7539), .ZN(MEM_stage_inst_dmem_n7544) );
NAND2_X1 MEM_stage_inst_dmem_U7671 ( .A1(MEM_stage_inst_dmem_ram_3790), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n7539) );
NAND2_X1 MEM_stage_inst_dmem_U7670 ( .A1(MEM_stage_inst_dmem_ram_3870), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n7540) );
NAND2_X1 MEM_stage_inst_dmem_U7669 ( .A1(MEM_stage_inst_dmem_n7538), .A2(MEM_stage_inst_dmem_n7537), .ZN(MEM_stage_inst_dmem_n7554) );
NOR2_X1 MEM_stage_inst_dmem_U7668 ( .A1(MEM_stage_inst_dmem_n7536), .A2(MEM_stage_inst_dmem_n7535), .ZN(MEM_stage_inst_dmem_n7537) );
NAND2_X1 MEM_stage_inst_dmem_U7667 ( .A1(MEM_stage_inst_dmem_n7534), .A2(MEM_stage_inst_dmem_n7533), .ZN(MEM_stage_inst_dmem_n7535) );
NAND2_X1 MEM_stage_inst_dmem_U7666 ( .A1(MEM_stage_inst_dmem_ram_3918), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n7533) );
NAND2_X1 MEM_stage_inst_dmem_U7665 ( .A1(MEM_stage_inst_dmem_ram_3806), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n7534) );
NAND2_X1 MEM_stage_inst_dmem_U7664 ( .A1(MEM_stage_inst_dmem_n7532), .A2(MEM_stage_inst_dmem_n7531), .ZN(MEM_stage_inst_dmem_n7536) );
NAND2_X1 MEM_stage_inst_dmem_U7663 ( .A1(MEM_stage_inst_dmem_ram_3854), .A2(MEM_stage_inst_dmem_n8472), .ZN(MEM_stage_inst_dmem_n7531) );
NAND2_X1 MEM_stage_inst_dmem_U7662 ( .A1(MEM_stage_inst_dmem_ram_3902), .A2(MEM_stage_inst_dmem_n8005), .ZN(MEM_stage_inst_dmem_n7532) );
NOR2_X1 MEM_stage_inst_dmem_U7661 ( .A1(MEM_stage_inst_dmem_n7530), .A2(MEM_stage_inst_dmem_n7529), .ZN(MEM_stage_inst_dmem_n7538) );
NAND2_X1 MEM_stage_inst_dmem_U7660 ( .A1(MEM_stage_inst_dmem_n7528), .A2(MEM_stage_inst_dmem_n7527), .ZN(MEM_stage_inst_dmem_n7529) );
NAND2_X1 MEM_stage_inst_dmem_U7659 ( .A1(MEM_stage_inst_dmem_ram_3454), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n7527) );
NAND2_X1 MEM_stage_inst_dmem_U7658 ( .A1(MEM_stage_inst_dmem_ram_3662), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n7528) );
NAND2_X1 MEM_stage_inst_dmem_U7657 ( .A1(MEM_stage_inst_dmem_n7526), .A2(MEM_stage_inst_dmem_n7525), .ZN(MEM_stage_inst_dmem_n7530) );
NAND2_X1 MEM_stage_inst_dmem_U7656 ( .A1(MEM_stage_inst_dmem_ram_3518), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n7525) );
NAND2_X1 MEM_stage_inst_dmem_U7655 ( .A1(MEM_stage_inst_dmem_ram_4014), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n7526) );
NOR2_X1 MEM_stage_inst_dmem_U7654 ( .A1(MEM_stage_inst_dmem_n7524), .A2(MEM_stage_inst_dmem_n7523), .ZN(MEM_stage_inst_dmem_n7556) );
NAND2_X1 MEM_stage_inst_dmem_U7653 ( .A1(MEM_stage_inst_dmem_n7522), .A2(MEM_stage_inst_dmem_n7521), .ZN(MEM_stage_inst_dmem_n7523) );
NOR2_X1 MEM_stage_inst_dmem_U7652 ( .A1(MEM_stage_inst_dmem_n7520), .A2(MEM_stage_inst_dmem_n7519), .ZN(MEM_stage_inst_dmem_n7521) );
NAND2_X1 MEM_stage_inst_dmem_U7651 ( .A1(MEM_stage_inst_dmem_n7518), .A2(MEM_stage_inst_dmem_n7517), .ZN(MEM_stage_inst_dmem_n7519) );
NAND2_X1 MEM_stage_inst_dmem_U7650 ( .A1(MEM_stage_inst_dmem_ram_3502), .A2(MEM_stage_inst_dmem_n4772), .ZN(MEM_stage_inst_dmem_n7517) );
NAND2_X1 MEM_stage_inst_dmem_U7649 ( .A1(MEM_stage_inst_dmem_ram_3886), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n7518) );
NAND2_X1 MEM_stage_inst_dmem_U7648 ( .A1(MEM_stage_inst_dmem_n7516), .A2(MEM_stage_inst_dmem_n7515), .ZN(MEM_stage_inst_dmem_n7520) );
NAND2_X1 MEM_stage_inst_dmem_U7647 ( .A1(MEM_stage_inst_dmem_ram_3182), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n7515) );
NAND2_X1 MEM_stage_inst_dmem_U7646 ( .A1(MEM_stage_inst_dmem_ram_3742), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n7516) );
NOR2_X1 MEM_stage_inst_dmem_U7645 ( .A1(MEM_stage_inst_dmem_n7514), .A2(MEM_stage_inst_dmem_n7513), .ZN(MEM_stage_inst_dmem_n7522) );
NAND2_X1 MEM_stage_inst_dmem_U7644 ( .A1(MEM_stage_inst_dmem_n7512), .A2(MEM_stage_inst_dmem_n7511), .ZN(MEM_stage_inst_dmem_n7513) );
NAND2_X1 MEM_stage_inst_dmem_U7643 ( .A1(MEM_stage_inst_dmem_ram_3486), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n7511) );
NAND2_X1 MEM_stage_inst_dmem_U7642 ( .A1(MEM_stage_inst_dmem_ram_3118), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n7512) );
NAND2_X1 MEM_stage_inst_dmem_U7641 ( .A1(MEM_stage_inst_dmem_n7510), .A2(MEM_stage_inst_dmem_n7509), .ZN(MEM_stage_inst_dmem_n7514) );
NAND2_X1 MEM_stage_inst_dmem_U7640 ( .A1(MEM_stage_inst_dmem_ram_3630), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n7509) );
NAND2_X1 MEM_stage_inst_dmem_U7639 ( .A1(MEM_stage_inst_dmem_ram_3694), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n7510) );
NAND2_X1 MEM_stage_inst_dmem_U7638 ( .A1(MEM_stage_inst_dmem_n7508), .A2(MEM_stage_inst_dmem_n7507), .ZN(MEM_stage_inst_dmem_n7524) );
NOR2_X1 MEM_stage_inst_dmem_U7637 ( .A1(MEM_stage_inst_dmem_n7506), .A2(MEM_stage_inst_dmem_n7505), .ZN(MEM_stage_inst_dmem_n7507) );
NAND2_X1 MEM_stage_inst_dmem_U7636 ( .A1(MEM_stage_inst_dmem_n7504), .A2(MEM_stage_inst_dmem_n7503), .ZN(MEM_stage_inst_dmem_n7505) );
NAND2_X1 MEM_stage_inst_dmem_U7635 ( .A1(MEM_stage_inst_dmem_ram_3406), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n7503) );
NAND2_X1 MEM_stage_inst_dmem_U7634 ( .A1(MEM_stage_inst_dmem_ram_3150), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n7504) );
NAND2_X1 MEM_stage_inst_dmem_U7633 ( .A1(MEM_stage_inst_dmem_n7502), .A2(MEM_stage_inst_dmem_n7501), .ZN(MEM_stage_inst_dmem_n7506) );
NAND2_X1 MEM_stage_inst_dmem_U7632 ( .A1(MEM_stage_inst_dmem_ram_3582), .A2(MEM_stage_inst_dmem_n64), .ZN(MEM_stage_inst_dmem_n7501) );
NAND2_X1 MEM_stage_inst_dmem_U7631 ( .A1(MEM_stage_inst_dmem_ram_3358), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n7502) );
NOR2_X1 MEM_stage_inst_dmem_U7630 ( .A1(MEM_stage_inst_dmem_n7500), .A2(MEM_stage_inst_dmem_n7499), .ZN(MEM_stage_inst_dmem_n7508) );
NAND2_X1 MEM_stage_inst_dmem_U7629 ( .A1(MEM_stage_inst_dmem_n7498), .A2(MEM_stage_inst_dmem_n7497), .ZN(MEM_stage_inst_dmem_n7499) );
NAND2_X1 MEM_stage_inst_dmem_U7628 ( .A1(MEM_stage_inst_dmem_ram_3102), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n7497) );
NAND2_X1 MEM_stage_inst_dmem_U7627 ( .A1(MEM_stage_inst_dmem_ram_3598), .A2(MEM_stage_inst_dmem_n8225), .ZN(MEM_stage_inst_dmem_n7498) );
NAND2_X1 MEM_stage_inst_dmem_U7626 ( .A1(MEM_stage_inst_dmem_n7496), .A2(MEM_stage_inst_dmem_n7495), .ZN(MEM_stage_inst_dmem_n7500) );
NAND2_X1 MEM_stage_inst_dmem_U7625 ( .A1(MEM_stage_inst_dmem_ram_3278), .A2(MEM_stage_inst_dmem_n8256), .ZN(MEM_stage_inst_dmem_n7495) );
NAND2_X1 MEM_stage_inst_dmem_U7624 ( .A1(MEM_stage_inst_dmem_ram_4062), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n7496) );
NAND2_X1 MEM_stage_inst_dmem_U7623 ( .A1(MEM_stage_inst_dmem_n7494), .A2(MEM_stage_inst_dmem_n7493), .ZN(MEM_stage_inst_mem_read_data_13) );
NOR2_X1 MEM_stage_inst_dmem_U7622 ( .A1(MEM_stage_inst_dmem_n7492), .A2(MEM_stage_inst_dmem_n7491), .ZN(MEM_stage_inst_dmem_n7493) );
NOR2_X1 MEM_stage_inst_dmem_U7621 ( .A1(MEM_stage_inst_dmem_n7490), .A2(MEM_stage_inst_dmem_n8152), .ZN(MEM_stage_inst_dmem_n7491) );
NOR2_X1 MEM_stage_inst_dmem_U7620 ( .A1(MEM_stage_inst_dmem_n7489), .A2(MEM_stage_inst_dmem_n7488), .ZN(MEM_stage_inst_dmem_n7490) );
NAND2_X1 MEM_stage_inst_dmem_U7619 ( .A1(MEM_stage_inst_dmem_n7487), .A2(MEM_stage_inst_dmem_n7486), .ZN(MEM_stage_inst_dmem_n7488) );
NOR2_X1 MEM_stage_inst_dmem_U7618 ( .A1(MEM_stage_inst_dmem_n7485), .A2(MEM_stage_inst_dmem_n7484), .ZN(MEM_stage_inst_dmem_n7486) );
NAND2_X1 MEM_stage_inst_dmem_U7617 ( .A1(MEM_stage_inst_dmem_n7483), .A2(MEM_stage_inst_dmem_n7482), .ZN(MEM_stage_inst_dmem_n7484) );
NOR2_X1 MEM_stage_inst_dmem_U7616 ( .A1(MEM_stage_inst_dmem_n7481), .A2(MEM_stage_inst_dmem_n7480), .ZN(MEM_stage_inst_dmem_n7482) );
NAND2_X1 MEM_stage_inst_dmem_U7615 ( .A1(MEM_stage_inst_dmem_n7479), .A2(MEM_stage_inst_dmem_n7478), .ZN(MEM_stage_inst_dmem_n7480) );
NAND2_X1 MEM_stage_inst_dmem_U7614 ( .A1(MEM_stage_inst_dmem_ram_1469), .A2(MEM_stage_inst_dmem_n7888), .ZN(MEM_stage_inst_dmem_n7478) );
NAND2_X1 MEM_stage_inst_dmem_U7613 ( .A1(MEM_stage_inst_dmem_ram_1325), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n7479) );
NAND2_X1 MEM_stage_inst_dmem_U7612 ( .A1(MEM_stage_inst_dmem_n7477), .A2(MEM_stage_inst_dmem_n7476), .ZN(MEM_stage_inst_dmem_n7481) );
NAND2_X1 MEM_stage_inst_dmem_U7611 ( .A1(MEM_stage_inst_dmem_ram_1085), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n7476) );
NAND2_X1 MEM_stage_inst_dmem_U7610 ( .A1(MEM_stage_inst_dmem_ram_1741), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n7477) );
NOR2_X1 MEM_stage_inst_dmem_U7609 ( .A1(MEM_stage_inst_dmem_n7475), .A2(MEM_stage_inst_dmem_n7474), .ZN(MEM_stage_inst_dmem_n7483) );
NAND2_X1 MEM_stage_inst_dmem_U7608 ( .A1(MEM_stage_inst_dmem_n7473), .A2(MEM_stage_inst_dmem_n7472), .ZN(MEM_stage_inst_dmem_n7474) );
NAND2_X1 MEM_stage_inst_dmem_U7607 ( .A1(MEM_stage_inst_dmem_ram_1677), .A2(MEM_stage_inst_dmem_n7960), .ZN(MEM_stage_inst_dmem_n7472) );
NAND2_X1 MEM_stage_inst_dmem_U7606 ( .A1(MEM_stage_inst_dmem_ram_1245), .A2(MEM_stage_inst_dmem_n51), .ZN(MEM_stage_inst_dmem_n7473) );
NAND2_X1 MEM_stage_inst_dmem_U7605 ( .A1(MEM_stage_inst_dmem_n7471), .A2(MEM_stage_inst_dmem_n7470), .ZN(MEM_stage_inst_dmem_n7475) );
NAND2_X1 MEM_stage_inst_dmem_U7604 ( .A1(MEM_stage_inst_dmem_ram_1917), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n7470) );
NAND2_X1 MEM_stage_inst_dmem_U7603 ( .A1(MEM_stage_inst_dmem_ram_1661), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n7471) );
NAND2_X1 MEM_stage_inst_dmem_U7602 ( .A1(MEM_stage_inst_dmem_n7469), .A2(MEM_stage_inst_dmem_n7468), .ZN(MEM_stage_inst_dmem_n7485) );
NOR2_X1 MEM_stage_inst_dmem_U7601 ( .A1(MEM_stage_inst_dmem_n7467), .A2(MEM_stage_inst_dmem_n7466), .ZN(MEM_stage_inst_dmem_n7468) );
NAND2_X1 MEM_stage_inst_dmem_U7600 ( .A1(MEM_stage_inst_dmem_n7465), .A2(MEM_stage_inst_dmem_n7464), .ZN(MEM_stage_inst_dmem_n7466) );
NAND2_X1 MEM_stage_inst_dmem_U7599 ( .A1(MEM_stage_inst_dmem_ram_1197), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n7464) );
NAND2_X1 MEM_stage_inst_dmem_U7598 ( .A1(MEM_stage_inst_dmem_ram_1773), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n7465) );
NAND2_X1 MEM_stage_inst_dmem_U7597 ( .A1(MEM_stage_inst_dmem_n7463), .A2(MEM_stage_inst_dmem_n7462), .ZN(MEM_stage_inst_dmem_n7467) );
NAND2_X1 MEM_stage_inst_dmem_U7596 ( .A1(MEM_stage_inst_dmem_ram_1533), .A2(MEM_stage_inst_dmem_n64), .ZN(MEM_stage_inst_dmem_n7462) );
NAND2_X1 MEM_stage_inst_dmem_U7595 ( .A1(MEM_stage_inst_dmem_ram_2013), .A2(MEM_stage_inst_dmem_n7895), .ZN(MEM_stage_inst_dmem_n7463) );
NOR2_X1 MEM_stage_inst_dmem_U7594 ( .A1(MEM_stage_inst_dmem_n7461), .A2(MEM_stage_inst_dmem_n7460), .ZN(MEM_stage_inst_dmem_n7469) );
NAND2_X1 MEM_stage_inst_dmem_U7593 ( .A1(MEM_stage_inst_dmem_n7459), .A2(MEM_stage_inst_dmem_n7458), .ZN(MEM_stage_inst_dmem_n7460) );
NAND2_X1 MEM_stage_inst_dmem_U7592 ( .A1(MEM_stage_inst_dmem_ram_1565), .A2(MEM_stage_inst_dmem_n7884), .ZN(MEM_stage_inst_dmem_n7458) );
NAND2_X1 MEM_stage_inst_dmem_U7591 ( .A1(MEM_stage_inst_dmem_ram_1757), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n7459) );
NAND2_X1 MEM_stage_inst_dmem_U7590 ( .A1(MEM_stage_inst_dmem_n7457), .A2(MEM_stage_inst_dmem_n7456), .ZN(MEM_stage_inst_dmem_n7461) );
NAND2_X1 MEM_stage_inst_dmem_U7589 ( .A1(MEM_stage_inst_dmem_ram_1165), .A2(MEM_stage_inst_dmem_n61), .ZN(MEM_stage_inst_dmem_n7456) );
NAND2_X1 MEM_stage_inst_dmem_U7588 ( .A1(MEM_stage_inst_dmem_ram_1373), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n7457) );
NOR2_X1 MEM_stage_inst_dmem_U7587 ( .A1(MEM_stage_inst_dmem_n7455), .A2(MEM_stage_inst_dmem_n7454), .ZN(MEM_stage_inst_dmem_n7487) );
NAND2_X1 MEM_stage_inst_dmem_U7586 ( .A1(MEM_stage_inst_dmem_n7453), .A2(MEM_stage_inst_dmem_n7452), .ZN(MEM_stage_inst_dmem_n7454) );
NOR2_X1 MEM_stage_inst_dmem_U7585 ( .A1(MEM_stage_inst_dmem_n7451), .A2(MEM_stage_inst_dmem_n7450), .ZN(MEM_stage_inst_dmem_n7452) );
NAND2_X1 MEM_stage_inst_dmem_U7584 ( .A1(MEM_stage_inst_dmem_n7449), .A2(MEM_stage_inst_dmem_n7448), .ZN(MEM_stage_inst_dmem_n7450) );
NAND2_X1 MEM_stage_inst_dmem_U7583 ( .A1(MEM_stage_inst_dmem_ram_2045), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n7448) );
NAND2_X1 MEM_stage_inst_dmem_U7582 ( .A1(MEM_stage_inst_dmem_ram_1293), .A2(MEM_stage_inst_dmem_n7898), .ZN(MEM_stage_inst_dmem_n7449) );
NAND2_X1 MEM_stage_inst_dmem_U7581 ( .A1(MEM_stage_inst_dmem_n7447), .A2(MEM_stage_inst_dmem_n7446), .ZN(MEM_stage_inst_dmem_n7451) );
NAND2_X1 MEM_stage_inst_dmem_U7580 ( .A1(MEM_stage_inst_dmem_ram_1357), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n7446) );
NAND2_X1 MEM_stage_inst_dmem_U7579 ( .A1(MEM_stage_inst_dmem_ram_1405), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n7447) );
NOR2_X1 MEM_stage_inst_dmem_U7578 ( .A1(MEM_stage_inst_dmem_n7445), .A2(MEM_stage_inst_dmem_n7444), .ZN(MEM_stage_inst_dmem_n7453) );
NAND2_X1 MEM_stage_inst_dmem_U7577 ( .A1(MEM_stage_inst_dmem_n7443), .A2(MEM_stage_inst_dmem_n7442), .ZN(MEM_stage_inst_dmem_n7444) );
NAND2_X1 MEM_stage_inst_dmem_U7576 ( .A1(MEM_stage_inst_dmem_ram_1517), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n7442) );
NAND2_X1 MEM_stage_inst_dmem_U7575 ( .A1(MEM_stage_inst_dmem_ram_1181), .A2(MEM_stage_inst_dmem_n7903), .ZN(MEM_stage_inst_dmem_n7443) );
NAND2_X1 MEM_stage_inst_dmem_U7574 ( .A1(MEM_stage_inst_dmem_n7441), .A2(MEM_stage_inst_dmem_n7440), .ZN(MEM_stage_inst_dmem_n7445) );
NAND2_X1 MEM_stage_inst_dmem_U7573 ( .A1(MEM_stage_inst_dmem_ram_1981), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n7440) );
NAND2_X1 MEM_stage_inst_dmem_U7572 ( .A1(MEM_stage_inst_dmem_ram_1581), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n7441) );
NAND2_X1 MEM_stage_inst_dmem_U7571 ( .A1(MEM_stage_inst_dmem_n7439), .A2(MEM_stage_inst_dmem_n7438), .ZN(MEM_stage_inst_dmem_n7455) );
NOR2_X1 MEM_stage_inst_dmem_U7570 ( .A1(MEM_stage_inst_dmem_n7437), .A2(MEM_stage_inst_dmem_n7436), .ZN(MEM_stage_inst_dmem_n7438) );
NAND2_X1 MEM_stage_inst_dmem_U7569 ( .A1(MEM_stage_inst_dmem_n7435), .A2(MEM_stage_inst_dmem_n7434), .ZN(MEM_stage_inst_dmem_n7436) );
NAND2_X1 MEM_stage_inst_dmem_U7568 ( .A1(MEM_stage_inst_dmem_ram_1933), .A2(MEM_stage_inst_dmem_n72), .ZN(MEM_stage_inst_dmem_n7434) );
NAND2_X1 MEM_stage_inst_dmem_U7567 ( .A1(MEM_stage_inst_dmem_ram_1837), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n7435) );
NAND2_X1 MEM_stage_inst_dmem_U7566 ( .A1(MEM_stage_inst_dmem_n7433), .A2(MEM_stage_inst_dmem_n7432), .ZN(MEM_stage_inst_dmem_n7437) );
NAND2_X1 MEM_stage_inst_dmem_U7565 ( .A1(MEM_stage_inst_dmem_ram_1597), .A2(MEM_stage_inst_dmem_n41), .ZN(MEM_stage_inst_dmem_n7432) );
NAND2_X1 MEM_stage_inst_dmem_U7564 ( .A1(MEM_stage_inst_dmem_ram_1309), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n7433) );
NOR2_X1 MEM_stage_inst_dmem_U7563 ( .A1(MEM_stage_inst_dmem_n7431), .A2(MEM_stage_inst_dmem_n7430), .ZN(MEM_stage_inst_dmem_n7439) );
NAND2_X1 MEM_stage_inst_dmem_U7562 ( .A1(MEM_stage_inst_dmem_n7429), .A2(MEM_stage_inst_dmem_n7428), .ZN(MEM_stage_inst_dmem_n7430) );
NAND2_X1 MEM_stage_inst_dmem_U7561 ( .A1(MEM_stage_inst_dmem_ram_1069), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n7428) );
NAND2_X1 MEM_stage_inst_dmem_U7560 ( .A1(MEM_stage_inst_dmem_ram_1853), .A2(MEM_stage_inst_dmem_n8005), .ZN(MEM_stage_inst_dmem_n7429) );
NAND2_X1 MEM_stage_inst_dmem_U7559 ( .A1(MEM_stage_inst_dmem_n7427), .A2(MEM_stage_inst_dmem_n7426), .ZN(MEM_stage_inst_dmem_n7431) );
NAND2_X1 MEM_stage_inst_dmem_U7558 ( .A1(MEM_stage_inst_dmem_ram_1437), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n7426) );
NAND2_X1 MEM_stage_inst_dmem_U7557 ( .A1(MEM_stage_inst_dmem_ram_1997), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n7427) );
NAND2_X1 MEM_stage_inst_dmem_U7556 ( .A1(MEM_stage_inst_dmem_n7425), .A2(MEM_stage_inst_dmem_n7424), .ZN(MEM_stage_inst_dmem_n7489) );
NOR2_X1 MEM_stage_inst_dmem_U7555 ( .A1(MEM_stage_inst_dmem_n7423), .A2(MEM_stage_inst_dmem_n7422), .ZN(MEM_stage_inst_dmem_n7424) );
NAND2_X1 MEM_stage_inst_dmem_U7554 ( .A1(MEM_stage_inst_dmem_n7421), .A2(MEM_stage_inst_dmem_n7420), .ZN(MEM_stage_inst_dmem_n7422) );
NOR2_X1 MEM_stage_inst_dmem_U7553 ( .A1(MEM_stage_inst_dmem_n7419), .A2(MEM_stage_inst_dmem_n7418), .ZN(MEM_stage_inst_dmem_n7420) );
NAND2_X1 MEM_stage_inst_dmem_U7552 ( .A1(MEM_stage_inst_dmem_n7417), .A2(MEM_stage_inst_dmem_n7416), .ZN(MEM_stage_inst_dmem_n7418) );
NAND2_X1 MEM_stage_inst_dmem_U7551 ( .A1(MEM_stage_inst_dmem_ram_1389), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n7416) );
NAND2_X1 MEM_stage_inst_dmem_U7550 ( .A1(MEM_stage_inst_dmem_ram_1421), .A2(MEM_stage_inst_dmem_n7930), .ZN(MEM_stage_inst_dmem_n7417) );
NAND2_X1 MEM_stage_inst_dmem_U7549 ( .A1(MEM_stage_inst_dmem_n7415), .A2(MEM_stage_inst_dmem_n7414), .ZN(MEM_stage_inst_dmem_n7419) );
NAND2_X1 MEM_stage_inst_dmem_U7548 ( .A1(MEM_stage_inst_dmem_ram_1949), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n7414) );
NAND2_X1 MEM_stage_inst_dmem_U7547 ( .A1(MEM_stage_inst_dmem_ram_1645), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n7415) );
NOR2_X1 MEM_stage_inst_dmem_U7546 ( .A1(MEM_stage_inst_dmem_n7413), .A2(MEM_stage_inst_dmem_n7412), .ZN(MEM_stage_inst_dmem_n7421) );
NAND2_X1 MEM_stage_inst_dmem_U7545 ( .A1(MEM_stage_inst_dmem_n7411), .A2(MEM_stage_inst_dmem_n7410), .ZN(MEM_stage_inst_dmem_n7412) );
NAND2_X1 MEM_stage_inst_dmem_U7544 ( .A1(MEM_stage_inst_dmem_ram_1805), .A2(MEM_stage_inst_dmem_n7992), .ZN(MEM_stage_inst_dmem_n7410) );
NAND2_X1 MEM_stage_inst_dmem_U7543 ( .A1(MEM_stage_inst_dmem_ram_1965), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n7411) );
NAND2_X1 MEM_stage_inst_dmem_U7542 ( .A1(MEM_stage_inst_dmem_n7409), .A2(MEM_stage_inst_dmem_n7408), .ZN(MEM_stage_inst_dmem_n7413) );
NAND2_X1 MEM_stage_inst_dmem_U7541 ( .A1(MEM_stage_inst_dmem_ram_1261), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n7408) );
NAND2_X1 MEM_stage_inst_dmem_U7540 ( .A1(MEM_stage_inst_dmem_ram_1133), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n7409) );
NAND2_X1 MEM_stage_inst_dmem_U7539 ( .A1(MEM_stage_inst_dmem_n7407), .A2(MEM_stage_inst_dmem_n7406), .ZN(MEM_stage_inst_dmem_n7423) );
NOR2_X1 MEM_stage_inst_dmem_U7538 ( .A1(MEM_stage_inst_dmem_n7405), .A2(MEM_stage_inst_dmem_n7404), .ZN(MEM_stage_inst_dmem_n7406) );
NAND2_X1 MEM_stage_inst_dmem_U7537 ( .A1(MEM_stage_inst_dmem_n7403), .A2(MEM_stage_inst_dmem_n7402), .ZN(MEM_stage_inst_dmem_n7404) );
NAND2_X1 MEM_stage_inst_dmem_U7536 ( .A1(MEM_stage_inst_dmem_ram_1885), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n7402) );
NAND2_X1 MEM_stage_inst_dmem_U7535 ( .A1(MEM_stage_inst_dmem_ram_1213), .A2(MEM_stage_inst_dmem_n7937), .ZN(MEM_stage_inst_dmem_n7403) );
NAND2_X1 MEM_stage_inst_dmem_U7534 ( .A1(MEM_stage_inst_dmem_n7401), .A2(MEM_stage_inst_dmem_n7400), .ZN(MEM_stage_inst_dmem_n7405) );
NAND2_X1 MEM_stage_inst_dmem_U7533 ( .A1(MEM_stage_inst_dmem_ram_1117), .A2(MEM_stage_inst_dmem_n7938), .ZN(MEM_stage_inst_dmem_n7400) );
NAND2_X1 MEM_stage_inst_dmem_U7532 ( .A1(MEM_stage_inst_dmem_ram_1613), .A2(MEM_stage_inst_dmem_n7973), .ZN(MEM_stage_inst_dmem_n7401) );
NOR2_X1 MEM_stage_inst_dmem_U7531 ( .A1(MEM_stage_inst_dmem_n7399), .A2(MEM_stage_inst_dmem_n7398), .ZN(MEM_stage_inst_dmem_n7407) );
NAND2_X1 MEM_stage_inst_dmem_U7530 ( .A1(MEM_stage_inst_dmem_n7397), .A2(MEM_stage_inst_dmem_n7396), .ZN(MEM_stage_inst_dmem_n7398) );
NAND2_X1 MEM_stage_inst_dmem_U7529 ( .A1(MEM_stage_inst_dmem_ram_1821), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n7396) );
NAND2_X1 MEM_stage_inst_dmem_U7528 ( .A1(MEM_stage_inst_dmem_ram_1037), .A2(MEM_stage_inst_dmem_n7953), .ZN(MEM_stage_inst_dmem_n7397) );
NAND2_X1 MEM_stage_inst_dmem_U7527 ( .A1(MEM_stage_inst_dmem_n7395), .A2(MEM_stage_inst_dmem_n7394), .ZN(MEM_stage_inst_dmem_n7399) );
NAND2_X1 MEM_stage_inst_dmem_U7526 ( .A1(MEM_stage_inst_dmem_ram_1869), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n7394) );
NAND2_X1 MEM_stage_inst_dmem_U7525 ( .A1(MEM_stage_inst_dmem_ram_1549), .A2(MEM_stage_inst_dmem_n71), .ZN(MEM_stage_inst_dmem_n7395) );
NOR2_X1 MEM_stage_inst_dmem_U7524 ( .A1(MEM_stage_inst_dmem_n7393), .A2(MEM_stage_inst_dmem_n7392), .ZN(MEM_stage_inst_dmem_n7425) );
NAND2_X1 MEM_stage_inst_dmem_U7523 ( .A1(MEM_stage_inst_dmem_n7391), .A2(MEM_stage_inst_dmem_n7390), .ZN(MEM_stage_inst_dmem_n7392) );
NOR2_X1 MEM_stage_inst_dmem_U7522 ( .A1(MEM_stage_inst_dmem_n7389), .A2(MEM_stage_inst_dmem_n7388), .ZN(MEM_stage_inst_dmem_n7390) );
NAND2_X1 MEM_stage_inst_dmem_U7521 ( .A1(MEM_stage_inst_dmem_n7387), .A2(MEM_stage_inst_dmem_n7386), .ZN(MEM_stage_inst_dmem_n7388) );
NAND2_X1 MEM_stage_inst_dmem_U7520 ( .A1(MEM_stage_inst_dmem_ram_1901), .A2(MEM_stage_inst_dmem_n7923), .ZN(MEM_stage_inst_dmem_n7386) );
NAND2_X1 MEM_stage_inst_dmem_U7519 ( .A1(MEM_stage_inst_dmem_ram_1485), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n7387) );
NAND2_X1 MEM_stage_inst_dmem_U7518 ( .A1(MEM_stage_inst_dmem_n7385), .A2(MEM_stage_inst_dmem_n7384), .ZN(MEM_stage_inst_dmem_n7389) );
NAND2_X1 MEM_stage_inst_dmem_U7517 ( .A1(MEM_stage_inst_dmem_ram_1341), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n7384) );
NAND2_X1 MEM_stage_inst_dmem_U7516 ( .A1(MEM_stage_inst_dmem_ram_1629), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n7385) );
NOR2_X1 MEM_stage_inst_dmem_U7515 ( .A1(MEM_stage_inst_dmem_n7383), .A2(MEM_stage_inst_dmem_n7382), .ZN(MEM_stage_inst_dmem_n7391) );
NAND2_X1 MEM_stage_inst_dmem_U7514 ( .A1(MEM_stage_inst_dmem_n7381), .A2(MEM_stage_inst_dmem_n7380), .ZN(MEM_stage_inst_dmem_n7382) );
NAND2_X1 MEM_stage_inst_dmem_U7513 ( .A1(MEM_stage_inst_dmem_ram_1277), .A2(MEM_stage_inst_dmem_n7914), .ZN(MEM_stage_inst_dmem_n7380) );
NAND2_X1 MEM_stage_inst_dmem_U7512 ( .A1(MEM_stage_inst_dmem_ram_1709), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n7381) );
NAND2_X1 MEM_stage_inst_dmem_U7511 ( .A1(MEM_stage_inst_dmem_n7379), .A2(MEM_stage_inst_dmem_n7378), .ZN(MEM_stage_inst_dmem_n7383) );
NAND2_X1 MEM_stage_inst_dmem_U7510 ( .A1(MEM_stage_inst_dmem_ram_1053), .A2(MEM_stage_inst_dmem_n7887), .ZN(MEM_stage_inst_dmem_n7378) );
NAND2_X1 MEM_stage_inst_dmem_U7509 ( .A1(MEM_stage_inst_dmem_ram_1693), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n7379) );
NAND2_X1 MEM_stage_inst_dmem_U7508 ( .A1(MEM_stage_inst_dmem_n7377), .A2(MEM_stage_inst_dmem_n7376), .ZN(MEM_stage_inst_dmem_n7393) );
NOR2_X1 MEM_stage_inst_dmem_U7507 ( .A1(MEM_stage_inst_dmem_n7375), .A2(MEM_stage_inst_dmem_n7374), .ZN(MEM_stage_inst_dmem_n7376) );
NAND2_X1 MEM_stage_inst_dmem_U7506 ( .A1(MEM_stage_inst_dmem_n7373), .A2(MEM_stage_inst_dmem_n7372), .ZN(MEM_stage_inst_dmem_n7374) );
NAND2_X1 MEM_stage_inst_dmem_U7505 ( .A1(MEM_stage_inst_dmem_ram_2029), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n7372) );
NAND2_X1 MEM_stage_inst_dmem_U7504 ( .A1(MEM_stage_inst_dmem_ram_1453), .A2(MEM_stage_inst_dmem_n4772), .ZN(MEM_stage_inst_dmem_n7373) );
NAND2_X1 MEM_stage_inst_dmem_U7503 ( .A1(MEM_stage_inst_dmem_n7371), .A2(MEM_stage_inst_dmem_n7370), .ZN(MEM_stage_inst_dmem_n7375) );
NAND2_X1 MEM_stage_inst_dmem_U7502 ( .A1(MEM_stage_inst_dmem_ram_1149), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n7370) );
NAND2_X1 MEM_stage_inst_dmem_U7501 ( .A1(MEM_stage_inst_dmem_ram_1501), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n7371) );
NOR2_X1 MEM_stage_inst_dmem_U7500 ( .A1(MEM_stage_inst_dmem_n7369), .A2(MEM_stage_inst_dmem_n7368), .ZN(MEM_stage_inst_dmem_n7377) );
NAND2_X1 MEM_stage_inst_dmem_U7499 ( .A1(MEM_stage_inst_dmem_n7367), .A2(MEM_stage_inst_dmem_n7366), .ZN(MEM_stage_inst_dmem_n7368) );
NAND2_X1 MEM_stage_inst_dmem_U7498 ( .A1(MEM_stage_inst_dmem_ram_1229), .A2(MEM_stage_inst_dmem_n36), .ZN(MEM_stage_inst_dmem_n7366) );
NAND2_X1 MEM_stage_inst_dmem_U7497 ( .A1(MEM_stage_inst_dmem_ram_1725), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n7367) );
NAND2_X1 MEM_stage_inst_dmem_U7496 ( .A1(MEM_stage_inst_dmem_n7365), .A2(MEM_stage_inst_dmem_n7364), .ZN(MEM_stage_inst_dmem_n7369) );
NAND2_X1 MEM_stage_inst_dmem_U7495 ( .A1(MEM_stage_inst_dmem_ram_1101), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n7364) );
NAND2_X1 MEM_stage_inst_dmem_U7494 ( .A1(MEM_stage_inst_dmem_ram_1789), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n7365) );
NOR2_X1 MEM_stage_inst_dmem_U7493 ( .A1(MEM_stage_inst_dmem_n7363), .A2(MEM_stage_inst_dmem_n8551), .ZN(MEM_stage_inst_dmem_n7492) );
NOR2_X1 MEM_stage_inst_dmem_U7492 ( .A1(MEM_stage_inst_dmem_n7362), .A2(MEM_stage_inst_dmem_n7361), .ZN(MEM_stage_inst_dmem_n7363) );
NAND2_X1 MEM_stage_inst_dmem_U7491 ( .A1(MEM_stage_inst_dmem_n7360), .A2(MEM_stage_inst_dmem_n7359), .ZN(MEM_stage_inst_dmem_n7361) );
NOR2_X1 MEM_stage_inst_dmem_U7490 ( .A1(MEM_stage_inst_dmem_n7358), .A2(MEM_stage_inst_dmem_n7357), .ZN(MEM_stage_inst_dmem_n7359) );
NAND2_X1 MEM_stage_inst_dmem_U7489 ( .A1(MEM_stage_inst_dmem_n7356), .A2(MEM_stage_inst_dmem_n7355), .ZN(MEM_stage_inst_dmem_n7357) );
NOR2_X1 MEM_stage_inst_dmem_U7488 ( .A1(MEM_stage_inst_dmem_n7354), .A2(MEM_stage_inst_dmem_n7353), .ZN(MEM_stage_inst_dmem_n7355) );
NAND2_X1 MEM_stage_inst_dmem_U7487 ( .A1(MEM_stage_inst_dmem_n7352), .A2(MEM_stage_inst_dmem_n7351), .ZN(MEM_stage_inst_dmem_n7353) );
NAND2_X1 MEM_stage_inst_dmem_U7486 ( .A1(MEM_stage_inst_dmem_ram_333), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n7351) );
NAND2_X1 MEM_stage_inst_dmem_U7485 ( .A1(MEM_stage_inst_dmem_ram_589), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n7352) );
NAND2_X1 MEM_stage_inst_dmem_U7484 ( .A1(MEM_stage_inst_dmem_n7350), .A2(MEM_stage_inst_dmem_n7349), .ZN(MEM_stage_inst_dmem_n7354) );
NAND2_X1 MEM_stage_inst_dmem_U7483 ( .A1(MEM_stage_inst_dmem_ram_717), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n7349) );
NAND2_X1 MEM_stage_inst_dmem_U7482 ( .A1(MEM_stage_inst_dmem_ram_621), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n7350) );
NOR2_X1 MEM_stage_inst_dmem_U7481 ( .A1(MEM_stage_inst_dmem_n7348), .A2(MEM_stage_inst_dmem_n7347), .ZN(MEM_stage_inst_dmem_n7356) );
NAND2_X1 MEM_stage_inst_dmem_U7480 ( .A1(MEM_stage_inst_dmem_n7346), .A2(MEM_stage_inst_dmem_n7345), .ZN(MEM_stage_inst_dmem_n7347) );
NAND2_X1 MEM_stage_inst_dmem_U7479 ( .A1(MEM_stage_inst_dmem_ram_525), .A2(MEM_stage_inst_dmem_n8225), .ZN(MEM_stage_inst_dmem_n7345) );
NAND2_X1 MEM_stage_inst_dmem_U7478 ( .A1(MEM_stage_inst_dmem_ram_269), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n7346) );
NAND2_X1 MEM_stage_inst_dmem_U7477 ( .A1(MEM_stage_inst_dmem_n7344), .A2(MEM_stage_inst_dmem_n7343), .ZN(MEM_stage_inst_dmem_n7348) );
NAND2_X1 MEM_stage_inst_dmem_U7476 ( .A1(MEM_stage_inst_dmem_ram_909), .A2(MEM_stage_inst_dmem_n8193), .ZN(MEM_stage_inst_dmem_n7343) );
NAND2_X1 MEM_stage_inst_dmem_U7475 ( .A1(MEM_stage_inst_dmem_ram_461), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n7344) );
NAND2_X1 MEM_stage_inst_dmem_U7474 ( .A1(MEM_stage_inst_dmem_n7342), .A2(MEM_stage_inst_dmem_n7341), .ZN(MEM_stage_inst_dmem_n7358) );
NOR2_X1 MEM_stage_inst_dmem_U7473 ( .A1(MEM_stage_inst_dmem_n7340), .A2(MEM_stage_inst_dmem_n7339), .ZN(MEM_stage_inst_dmem_n7341) );
NAND2_X1 MEM_stage_inst_dmem_U7472 ( .A1(MEM_stage_inst_dmem_n7338), .A2(MEM_stage_inst_dmem_n7337), .ZN(MEM_stage_inst_dmem_n7339) );
NAND2_X1 MEM_stage_inst_dmem_U7471 ( .A1(MEM_stage_inst_dmem_ram_429), .A2(MEM_stage_inst_dmem_n4772), .ZN(MEM_stage_inst_dmem_n7337) );
NAND2_X1 MEM_stage_inst_dmem_U7470 ( .A1(MEM_stage_inst_dmem_ram_813), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n7338) );
NAND2_X1 MEM_stage_inst_dmem_U7469 ( .A1(MEM_stage_inst_dmem_n7336), .A2(MEM_stage_inst_dmem_n7335), .ZN(MEM_stage_inst_dmem_n7340) );
NAND2_X1 MEM_stage_inst_dmem_U7468 ( .A1(MEM_stage_inst_dmem_ram_445), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n7335) );
NAND2_X1 MEM_stage_inst_dmem_U7467 ( .A1(MEM_stage_inst_dmem_ram_173), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n7336) );
NOR2_X1 MEM_stage_inst_dmem_U7466 ( .A1(MEM_stage_inst_dmem_n7334), .A2(MEM_stage_inst_dmem_n7333), .ZN(MEM_stage_inst_dmem_n7342) );
NAND2_X1 MEM_stage_inst_dmem_U7465 ( .A1(MEM_stage_inst_dmem_n7332), .A2(MEM_stage_inst_dmem_n7331), .ZN(MEM_stage_inst_dmem_n7333) );
NAND2_X1 MEM_stage_inst_dmem_U7464 ( .A1(MEM_stage_inst_dmem_ram_573), .A2(MEM_stage_inst_dmem_n8169), .ZN(MEM_stage_inst_dmem_n7331) );
NAND2_X1 MEM_stage_inst_dmem_U7463 ( .A1(MEM_stage_inst_dmem_ram_477), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n7332) );
NAND2_X1 MEM_stage_inst_dmem_U7462 ( .A1(MEM_stage_inst_dmem_n7330), .A2(MEM_stage_inst_dmem_n7329), .ZN(MEM_stage_inst_dmem_n7334) );
NAND2_X1 MEM_stage_inst_dmem_U7461 ( .A1(MEM_stage_inst_dmem_ram_237), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n7329) );
NAND2_X1 MEM_stage_inst_dmem_U7460 ( .A1(MEM_stage_inst_dmem_ram_109), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n7330) );
NOR2_X1 MEM_stage_inst_dmem_U7459 ( .A1(MEM_stage_inst_dmem_n7328), .A2(MEM_stage_inst_dmem_n7327), .ZN(MEM_stage_inst_dmem_n7360) );
NAND2_X1 MEM_stage_inst_dmem_U7458 ( .A1(MEM_stage_inst_dmem_n7326), .A2(MEM_stage_inst_dmem_n7325), .ZN(MEM_stage_inst_dmem_n7327) );
NOR2_X1 MEM_stage_inst_dmem_U7457 ( .A1(MEM_stage_inst_dmem_n7324), .A2(MEM_stage_inst_dmem_n7323), .ZN(MEM_stage_inst_dmem_n7325) );
NAND2_X1 MEM_stage_inst_dmem_U7456 ( .A1(MEM_stage_inst_dmem_n7322), .A2(MEM_stage_inst_dmem_n7321), .ZN(MEM_stage_inst_dmem_n7323) );
NAND2_X1 MEM_stage_inst_dmem_U7455 ( .A1(MEM_stage_inst_dmem_ram_653), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n7321) );
NAND2_X1 MEM_stage_inst_dmem_U7454 ( .A1(MEM_stage_inst_dmem_ram_733), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n7322) );
NAND2_X1 MEM_stage_inst_dmem_U7453 ( .A1(MEM_stage_inst_dmem_n7320), .A2(MEM_stage_inst_dmem_n7319), .ZN(MEM_stage_inst_dmem_n7324) );
NAND2_X1 MEM_stage_inst_dmem_U7452 ( .A1(MEM_stage_inst_dmem_ram_605), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n7319) );
NAND2_X1 MEM_stage_inst_dmem_U7451 ( .A1(MEM_stage_inst_dmem_ram_381), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n7320) );
NOR2_X1 MEM_stage_inst_dmem_U7450 ( .A1(MEM_stage_inst_dmem_n7318), .A2(MEM_stage_inst_dmem_n7317), .ZN(MEM_stage_inst_dmem_n7326) );
NAND2_X1 MEM_stage_inst_dmem_U7449 ( .A1(MEM_stage_inst_dmem_n7316), .A2(MEM_stage_inst_dmem_n7315), .ZN(MEM_stage_inst_dmem_n7317) );
NAND2_X1 MEM_stage_inst_dmem_U7448 ( .A1(MEM_stage_inst_dmem_ram_493), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n7315) );
NAND2_X1 MEM_stage_inst_dmem_U7447 ( .A1(MEM_stage_inst_dmem_ram_829), .A2(MEM_stage_inst_dmem_n8005), .ZN(MEM_stage_inst_dmem_n7316) );
NAND2_X1 MEM_stage_inst_dmem_U7446 ( .A1(MEM_stage_inst_dmem_n7314), .A2(MEM_stage_inst_dmem_n7313), .ZN(MEM_stage_inst_dmem_n7318) );
NAND2_X1 MEM_stage_inst_dmem_U7445 ( .A1(MEM_stage_inst_dmem_ram_93), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n7313) );
NAND2_X1 MEM_stage_inst_dmem_U7444 ( .A1(MEM_stage_inst_dmem_ram_157), .A2(MEM_stage_inst_dmem_n44), .ZN(MEM_stage_inst_dmem_n7314) );
NAND2_X1 MEM_stage_inst_dmem_U7443 ( .A1(MEM_stage_inst_dmem_n7312), .A2(MEM_stage_inst_dmem_n7311), .ZN(MEM_stage_inst_dmem_n7328) );
NOR2_X1 MEM_stage_inst_dmem_U7442 ( .A1(MEM_stage_inst_dmem_n7310), .A2(MEM_stage_inst_dmem_n7309), .ZN(MEM_stage_inst_dmem_n7311) );
NAND2_X1 MEM_stage_inst_dmem_U7441 ( .A1(MEM_stage_inst_dmem_n7308), .A2(MEM_stage_inst_dmem_n7307), .ZN(MEM_stage_inst_dmem_n7309) );
NAND2_X1 MEM_stage_inst_dmem_U7440 ( .A1(MEM_stage_inst_dmem_ram_141), .A2(MEM_stage_inst_dmem_n8174), .ZN(MEM_stage_inst_dmem_n7307) );
NAND2_X1 MEM_stage_inst_dmem_U7439 ( .A1(MEM_stage_inst_dmem_ram_685), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n7308) );
NAND2_X1 MEM_stage_inst_dmem_U7438 ( .A1(MEM_stage_inst_dmem_n7306), .A2(MEM_stage_inst_dmem_n7305), .ZN(MEM_stage_inst_dmem_n7310) );
NAND2_X1 MEM_stage_inst_dmem_U7437 ( .A1(MEM_stage_inst_dmem_ram_317), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n7305) );
NAND2_X1 MEM_stage_inst_dmem_U7436 ( .A1(MEM_stage_inst_dmem_ram_397), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n7306) );
NOR2_X1 MEM_stage_inst_dmem_U7435 ( .A1(MEM_stage_inst_dmem_n7304), .A2(MEM_stage_inst_dmem_n7303), .ZN(MEM_stage_inst_dmem_n7312) );
NAND2_X1 MEM_stage_inst_dmem_U7434 ( .A1(MEM_stage_inst_dmem_n7302), .A2(MEM_stage_inst_dmem_n7301), .ZN(MEM_stage_inst_dmem_n7303) );
NAND2_X1 MEM_stage_inst_dmem_U7433 ( .A1(MEM_stage_inst_dmem_ram_893), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n7301) );
NAND2_X1 MEM_stage_inst_dmem_U7432 ( .A1(MEM_stage_inst_dmem_ram_77), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n7302) );
NAND2_X1 MEM_stage_inst_dmem_U7431 ( .A1(MEM_stage_inst_dmem_n7300), .A2(MEM_stage_inst_dmem_n7299), .ZN(MEM_stage_inst_dmem_n7304) );
NAND2_X1 MEM_stage_inst_dmem_U7430 ( .A1(MEM_stage_inst_dmem_ram_1005), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n7299) );
NAND2_X1 MEM_stage_inst_dmem_U7429 ( .A1(MEM_stage_inst_dmem_ram_941), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n7300) );
NAND2_X1 MEM_stage_inst_dmem_U7428 ( .A1(MEM_stage_inst_dmem_n7298), .A2(MEM_stage_inst_dmem_n7297), .ZN(MEM_stage_inst_dmem_n7362) );
NOR2_X1 MEM_stage_inst_dmem_U7427 ( .A1(MEM_stage_inst_dmem_n7296), .A2(MEM_stage_inst_dmem_n7295), .ZN(MEM_stage_inst_dmem_n7297) );
NAND2_X1 MEM_stage_inst_dmem_U7426 ( .A1(MEM_stage_inst_dmem_n7294), .A2(MEM_stage_inst_dmem_n7293), .ZN(MEM_stage_inst_dmem_n7295) );
NOR2_X1 MEM_stage_inst_dmem_U7425 ( .A1(MEM_stage_inst_dmem_n7292), .A2(MEM_stage_inst_dmem_n7291), .ZN(MEM_stage_inst_dmem_n7293) );
NAND2_X1 MEM_stage_inst_dmem_U7424 ( .A1(MEM_stage_inst_dmem_n7290), .A2(MEM_stage_inst_dmem_n7289), .ZN(MEM_stage_inst_dmem_n7291) );
NAND2_X1 MEM_stage_inst_dmem_U7423 ( .A1(MEM_stage_inst_dmem_ram_29), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n7289) );
NAND2_X1 MEM_stage_inst_dmem_U7422 ( .A1(MEM_stage_inst_dmem_ram_797), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n7290) );
NAND2_X1 MEM_stage_inst_dmem_U7421 ( .A1(MEM_stage_inst_dmem_n7288), .A2(MEM_stage_inst_dmem_n7287), .ZN(MEM_stage_inst_dmem_n7292) );
NAND2_X1 MEM_stage_inst_dmem_U7420 ( .A1(MEM_stage_inst_dmem_ram_61), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n7287) );
NAND2_X1 MEM_stage_inst_dmem_U7419 ( .A1(MEM_stage_inst_dmem_ram_45), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n7288) );
NOR2_X1 MEM_stage_inst_dmem_U7418 ( .A1(MEM_stage_inst_dmem_n7286), .A2(MEM_stage_inst_dmem_n7285), .ZN(MEM_stage_inst_dmem_n7294) );
NAND2_X1 MEM_stage_inst_dmem_U7417 ( .A1(MEM_stage_inst_dmem_n7284), .A2(MEM_stage_inst_dmem_n7283), .ZN(MEM_stage_inst_dmem_n7285) );
NAND2_X1 MEM_stage_inst_dmem_U7416 ( .A1(MEM_stage_inst_dmem_ram_509), .A2(MEM_stage_inst_dmem_n64), .ZN(MEM_stage_inst_dmem_n7283) );
NAND2_X1 MEM_stage_inst_dmem_U7415 ( .A1(MEM_stage_inst_dmem_ram_541), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n7284) );
NAND2_X1 MEM_stage_inst_dmem_U7414 ( .A1(MEM_stage_inst_dmem_n7282), .A2(MEM_stage_inst_dmem_n7281), .ZN(MEM_stage_inst_dmem_n7286) );
NAND2_X1 MEM_stage_inst_dmem_U7413 ( .A1(MEM_stage_inst_dmem_ram_301), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n7281) );
NAND2_X1 MEM_stage_inst_dmem_U7412 ( .A1(MEM_stage_inst_dmem_ram_349), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n7282) );
NAND2_X1 MEM_stage_inst_dmem_U7411 ( .A1(MEM_stage_inst_dmem_n7280), .A2(MEM_stage_inst_dmem_n7279), .ZN(MEM_stage_inst_dmem_n7296) );
NOR2_X1 MEM_stage_inst_dmem_U7410 ( .A1(MEM_stage_inst_dmem_n7278), .A2(MEM_stage_inst_dmem_n7277), .ZN(MEM_stage_inst_dmem_n7279) );
NAND2_X1 MEM_stage_inst_dmem_U7409 ( .A1(MEM_stage_inst_dmem_n7276), .A2(MEM_stage_inst_dmem_n7275), .ZN(MEM_stage_inst_dmem_n7277) );
NAND2_X1 MEM_stage_inst_dmem_U7408 ( .A1(MEM_stage_inst_dmem_ram_925), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n7275) );
NAND2_X1 MEM_stage_inst_dmem_U7407 ( .A1(MEM_stage_inst_dmem_ram_701), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n7276) );
NAND2_X1 MEM_stage_inst_dmem_U7406 ( .A1(MEM_stage_inst_dmem_n7274), .A2(MEM_stage_inst_dmem_n7273), .ZN(MEM_stage_inst_dmem_n7278) );
NAND2_X1 MEM_stage_inst_dmem_U7405 ( .A1(MEM_stage_inst_dmem_ram_877), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n7273) );
NAND2_X1 MEM_stage_inst_dmem_U7404 ( .A1(MEM_stage_inst_dmem_ram_221), .A2(MEM_stage_inst_dmem_n8206), .ZN(MEM_stage_inst_dmem_n7274) );
NOR2_X1 MEM_stage_inst_dmem_U7403 ( .A1(MEM_stage_inst_dmem_n7272), .A2(MEM_stage_inst_dmem_n7271), .ZN(MEM_stage_inst_dmem_n7280) );
NAND2_X1 MEM_stage_inst_dmem_U7402 ( .A1(MEM_stage_inst_dmem_n7270), .A2(MEM_stage_inst_dmem_n7269), .ZN(MEM_stage_inst_dmem_n7271) );
NAND2_X1 MEM_stage_inst_dmem_U7401 ( .A1(MEM_stage_inst_dmem_ram_365), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n7269) );
NAND2_X1 MEM_stage_inst_dmem_U7400 ( .A1(MEM_stage_inst_dmem_ram_1021), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n7270) );
NAND2_X1 MEM_stage_inst_dmem_U7399 ( .A1(MEM_stage_inst_dmem_n7268), .A2(MEM_stage_inst_dmem_n7267), .ZN(MEM_stage_inst_dmem_n7272) );
NAND2_X1 MEM_stage_inst_dmem_U7398 ( .A1(MEM_stage_inst_dmem_ram_957), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n7267) );
NAND2_X1 MEM_stage_inst_dmem_U7397 ( .A1(MEM_stage_inst_dmem_ram_253), .A2(MEM_stage_inst_dmem_n7914), .ZN(MEM_stage_inst_dmem_n7268) );
NOR2_X1 MEM_stage_inst_dmem_U7396 ( .A1(MEM_stage_inst_dmem_n7266), .A2(MEM_stage_inst_dmem_n7265), .ZN(MEM_stage_inst_dmem_n7298) );
NAND2_X1 MEM_stage_inst_dmem_U7395 ( .A1(MEM_stage_inst_dmem_n7264), .A2(MEM_stage_inst_dmem_n7263), .ZN(MEM_stage_inst_dmem_n7265) );
NOR2_X1 MEM_stage_inst_dmem_U7394 ( .A1(MEM_stage_inst_dmem_n7262), .A2(MEM_stage_inst_dmem_n7261), .ZN(MEM_stage_inst_dmem_n7263) );
NAND2_X1 MEM_stage_inst_dmem_U7393 ( .A1(MEM_stage_inst_dmem_n7260), .A2(MEM_stage_inst_dmem_n7259), .ZN(MEM_stage_inst_dmem_n7261) );
NAND2_X1 MEM_stage_inst_dmem_U7392 ( .A1(MEM_stage_inst_dmem_ram_781), .A2(MEM_stage_inst_dmem_n8472), .ZN(MEM_stage_inst_dmem_n7259) );
NAND2_X1 MEM_stage_inst_dmem_U7391 ( .A1(MEM_stage_inst_dmem_ram_861), .A2(MEM_stage_inst_dmem_n3141), .ZN(MEM_stage_inst_dmem_n7260) );
NAND2_X1 MEM_stage_inst_dmem_U7390 ( .A1(MEM_stage_inst_dmem_n7258), .A2(MEM_stage_inst_dmem_n7257), .ZN(MEM_stage_inst_dmem_n7262) );
NAND2_X1 MEM_stage_inst_dmem_U7389 ( .A1(MEM_stage_inst_dmem_ram_973), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n7257) );
NAND2_X1 MEM_stage_inst_dmem_U7388 ( .A1(MEM_stage_inst_dmem_ram_749), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n7258) );
NOR2_X1 MEM_stage_inst_dmem_U7387 ( .A1(MEM_stage_inst_dmem_n7256), .A2(MEM_stage_inst_dmem_n7255), .ZN(MEM_stage_inst_dmem_n7264) );
NAND2_X1 MEM_stage_inst_dmem_U7386 ( .A1(MEM_stage_inst_dmem_n7254), .A2(MEM_stage_inst_dmem_n7253), .ZN(MEM_stage_inst_dmem_n7255) );
NAND2_X1 MEM_stage_inst_dmem_U7385 ( .A1(MEM_stage_inst_dmem_ram_845), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n7253) );
NAND2_X1 MEM_stage_inst_dmem_U7384 ( .A1(MEM_stage_inst_dmem_ram_285), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n7254) );
NAND2_X1 MEM_stage_inst_dmem_U7383 ( .A1(MEM_stage_inst_dmem_n7252), .A2(MEM_stage_inst_dmem_n7251), .ZN(MEM_stage_inst_dmem_n7256) );
NAND2_X1 MEM_stage_inst_dmem_U7382 ( .A1(MEM_stage_inst_dmem_ram_125), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n7251) );
NAND2_X1 MEM_stage_inst_dmem_U7381 ( .A1(MEM_stage_inst_dmem_ram_189), .A2(MEM_stage_inst_dmem_n8434), .ZN(MEM_stage_inst_dmem_n7252) );
NAND2_X1 MEM_stage_inst_dmem_U7380 ( .A1(MEM_stage_inst_dmem_n7250), .A2(MEM_stage_inst_dmem_n7249), .ZN(MEM_stage_inst_dmem_n7266) );
NOR2_X1 MEM_stage_inst_dmem_U7379 ( .A1(MEM_stage_inst_dmem_n7248), .A2(MEM_stage_inst_dmem_n7247), .ZN(MEM_stage_inst_dmem_n7249) );
NAND2_X1 MEM_stage_inst_dmem_U7378 ( .A1(MEM_stage_inst_dmem_n7246), .A2(MEM_stage_inst_dmem_n7245), .ZN(MEM_stage_inst_dmem_n7247) );
NAND2_X1 MEM_stage_inst_dmem_U7377 ( .A1(MEM_stage_inst_dmem_ram_989), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n7245) );
NAND2_X1 MEM_stage_inst_dmem_U7376 ( .A1(MEM_stage_inst_dmem_ram_637), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n7246) );
NAND2_X1 MEM_stage_inst_dmem_U7375 ( .A1(MEM_stage_inst_dmem_n7244), .A2(MEM_stage_inst_dmem_n7243), .ZN(MEM_stage_inst_dmem_n7248) );
NAND2_X1 MEM_stage_inst_dmem_U7374 ( .A1(MEM_stage_inst_dmem_ram_765), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n7243) );
NAND2_X1 MEM_stage_inst_dmem_U7373 ( .A1(MEM_stage_inst_dmem_ram_669), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n7244) );
NOR2_X1 MEM_stage_inst_dmem_U7372 ( .A1(MEM_stage_inst_dmem_n7242), .A2(MEM_stage_inst_dmem_n7241), .ZN(MEM_stage_inst_dmem_n7250) );
NAND2_X1 MEM_stage_inst_dmem_U7371 ( .A1(MEM_stage_inst_dmem_n7240), .A2(MEM_stage_inst_dmem_n7239), .ZN(MEM_stage_inst_dmem_n7241) );
NAND2_X1 MEM_stage_inst_dmem_U7370 ( .A1(MEM_stage_inst_dmem_ram_413), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n7239) );
NAND2_X1 MEM_stage_inst_dmem_U7369 ( .A1(MEM_stage_inst_dmem_ram_557), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n7240) );
NAND2_X1 MEM_stage_inst_dmem_U7368 ( .A1(MEM_stage_inst_dmem_n7238), .A2(MEM_stage_inst_dmem_n7237), .ZN(MEM_stage_inst_dmem_n7242) );
NAND2_X1 MEM_stage_inst_dmem_U7367 ( .A1(MEM_stage_inst_dmem_ram_205), .A2(MEM_stage_inst_dmem_n8256), .ZN(MEM_stage_inst_dmem_n7237) );
NAND2_X1 MEM_stage_inst_dmem_U7366 ( .A1(MEM_stage_inst_dmem_ram_13), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n7238) );
NOR2_X1 MEM_stage_inst_dmem_U7365 ( .A1(MEM_stage_inst_dmem_n7236), .A2(MEM_stage_inst_dmem_n7235), .ZN(MEM_stage_inst_dmem_n7494) );
NOR2_X1 MEM_stage_inst_dmem_U7364 ( .A1(MEM_stage_inst_dmem_n7234), .A2(MEM_stage_inst_dmem_n8286), .ZN(MEM_stage_inst_dmem_n7235) );
NOR2_X1 MEM_stage_inst_dmem_U7363 ( .A1(MEM_stage_inst_dmem_n7233), .A2(MEM_stage_inst_dmem_n7232), .ZN(MEM_stage_inst_dmem_n7234) );
NAND2_X1 MEM_stage_inst_dmem_U7362 ( .A1(MEM_stage_inst_dmem_n7231), .A2(MEM_stage_inst_dmem_n7230), .ZN(MEM_stage_inst_dmem_n7232) );
NOR2_X1 MEM_stage_inst_dmem_U7361 ( .A1(MEM_stage_inst_dmem_n7229), .A2(MEM_stage_inst_dmem_n7228), .ZN(MEM_stage_inst_dmem_n7230) );
NAND2_X1 MEM_stage_inst_dmem_U7360 ( .A1(MEM_stage_inst_dmem_n7227), .A2(MEM_stage_inst_dmem_n7226), .ZN(MEM_stage_inst_dmem_n7228) );
NOR2_X1 MEM_stage_inst_dmem_U7359 ( .A1(MEM_stage_inst_dmem_n7225), .A2(MEM_stage_inst_dmem_n7224), .ZN(MEM_stage_inst_dmem_n7226) );
NAND2_X1 MEM_stage_inst_dmem_U7358 ( .A1(MEM_stage_inst_dmem_n7223), .A2(MEM_stage_inst_dmem_n7222), .ZN(MEM_stage_inst_dmem_n7224) );
NAND2_X1 MEM_stage_inst_dmem_U7357 ( .A1(MEM_stage_inst_dmem_ram_2301), .A2(MEM_stage_inst_dmem_n7914), .ZN(MEM_stage_inst_dmem_n7222) );
NAND2_X1 MEM_stage_inst_dmem_U7356 ( .A1(MEM_stage_inst_dmem_ram_2589), .A2(MEM_stage_inst_dmem_n7884), .ZN(MEM_stage_inst_dmem_n7223) );
NAND2_X1 MEM_stage_inst_dmem_U7355 ( .A1(MEM_stage_inst_dmem_n7221), .A2(MEM_stage_inst_dmem_n7220), .ZN(MEM_stage_inst_dmem_n7225) );
NAND2_X1 MEM_stage_inst_dmem_U7354 ( .A1(MEM_stage_inst_dmem_ram_2861), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n7220) );
NAND2_X1 MEM_stage_inst_dmem_U7353 ( .A1(MEM_stage_inst_dmem_ram_2221), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n7221) );
NOR2_X1 MEM_stage_inst_dmem_U7352 ( .A1(MEM_stage_inst_dmem_n7219), .A2(MEM_stage_inst_dmem_n7218), .ZN(MEM_stage_inst_dmem_n7227) );
NAND2_X1 MEM_stage_inst_dmem_U7351 ( .A1(MEM_stage_inst_dmem_n7217), .A2(MEM_stage_inst_dmem_n7216), .ZN(MEM_stage_inst_dmem_n7218) );
NAND2_X1 MEM_stage_inst_dmem_U7350 ( .A1(MEM_stage_inst_dmem_ram_2173), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n7216) );
NAND2_X1 MEM_stage_inst_dmem_U7349 ( .A1(MEM_stage_inst_dmem_ram_2749), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n7217) );
NAND2_X1 MEM_stage_inst_dmem_U7348 ( .A1(MEM_stage_inst_dmem_n7215), .A2(MEM_stage_inst_dmem_n7214), .ZN(MEM_stage_inst_dmem_n7219) );
NAND2_X1 MEM_stage_inst_dmem_U7347 ( .A1(MEM_stage_inst_dmem_ram_2829), .A2(MEM_stage_inst_dmem_n7992), .ZN(MEM_stage_inst_dmem_n7214) );
NAND2_X1 MEM_stage_inst_dmem_U7346 ( .A1(MEM_stage_inst_dmem_ram_2317), .A2(MEM_stage_inst_dmem_n7898), .ZN(MEM_stage_inst_dmem_n7215) );
NAND2_X1 MEM_stage_inst_dmem_U7345 ( .A1(MEM_stage_inst_dmem_n7213), .A2(MEM_stage_inst_dmem_n7212), .ZN(MEM_stage_inst_dmem_n7229) );
NOR2_X1 MEM_stage_inst_dmem_U7344 ( .A1(MEM_stage_inst_dmem_n7211), .A2(MEM_stage_inst_dmem_n7210), .ZN(MEM_stage_inst_dmem_n7212) );
NAND2_X1 MEM_stage_inst_dmem_U7343 ( .A1(MEM_stage_inst_dmem_n7209), .A2(MEM_stage_inst_dmem_n7208), .ZN(MEM_stage_inst_dmem_n7210) );
NAND2_X1 MEM_stage_inst_dmem_U7342 ( .A1(MEM_stage_inst_dmem_ram_2685), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n7208) );
NAND2_X1 MEM_stage_inst_dmem_U7341 ( .A1(MEM_stage_inst_dmem_ram_2845), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n7209) );
NAND2_X1 MEM_stage_inst_dmem_U7340 ( .A1(MEM_stage_inst_dmem_n7207), .A2(MEM_stage_inst_dmem_n7206), .ZN(MEM_stage_inst_dmem_n7211) );
NAND2_X1 MEM_stage_inst_dmem_U7339 ( .A1(MEM_stage_inst_dmem_ram_2333), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n7206) );
NAND2_X1 MEM_stage_inst_dmem_U7338 ( .A1(MEM_stage_inst_dmem_ram_2269), .A2(MEM_stage_inst_dmem_n51), .ZN(MEM_stage_inst_dmem_n7207) );
NOR2_X1 MEM_stage_inst_dmem_U7337 ( .A1(MEM_stage_inst_dmem_n7205), .A2(MEM_stage_inst_dmem_n7204), .ZN(MEM_stage_inst_dmem_n7213) );
NAND2_X1 MEM_stage_inst_dmem_U7336 ( .A1(MEM_stage_inst_dmem_n7203), .A2(MEM_stage_inst_dmem_n7202), .ZN(MEM_stage_inst_dmem_n7204) );
NAND2_X1 MEM_stage_inst_dmem_U7335 ( .A1(MEM_stage_inst_dmem_ram_2877), .A2(MEM_stage_inst_dmem_n8005), .ZN(MEM_stage_inst_dmem_n7202) );
NAND2_X1 MEM_stage_inst_dmem_U7334 ( .A1(MEM_stage_inst_dmem_ram_3069), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n7203) );
NAND2_X1 MEM_stage_inst_dmem_U7333 ( .A1(MEM_stage_inst_dmem_n7201), .A2(MEM_stage_inst_dmem_n7200), .ZN(MEM_stage_inst_dmem_n7205) );
NAND2_X1 MEM_stage_inst_dmem_U7332 ( .A1(MEM_stage_inst_dmem_ram_2669), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n7200) );
NAND2_X1 MEM_stage_inst_dmem_U7331 ( .A1(MEM_stage_inst_dmem_ram_2637), .A2(MEM_stage_inst_dmem_n7973), .ZN(MEM_stage_inst_dmem_n7201) );
NOR2_X1 MEM_stage_inst_dmem_U7330 ( .A1(MEM_stage_inst_dmem_n7199), .A2(MEM_stage_inst_dmem_n7198), .ZN(MEM_stage_inst_dmem_n7231) );
NAND2_X1 MEM_stage_inst_dmem_U7329 ( .A1(MEM_stage_inst_dmem_n7197), .A2(MEM_stage_inst_dmem_n7196), .ZN(MEM_stage_inst_dmem_n7198) );
NOR2_X1 MEM_stage_inst_dmem_U7328 ( .A1(MEM_stage_inst_dmem_n7195), .A2(MEM_stage_inst_dmem_n7194), .ZN(MEM_stage_inst_dmem_n7196) );
NAND2_X1 MEM_stage_inst_dmem_U7327 ( .A1(MEM_stage_inst_dmem_n7193), .A2(MEM_stage_inst_dmem_n7192), .ZN(MEM_stage_inst_dmem_n7194) );
NAND2_X1 MEM_stage_inst_dmem_U7326 ( .A1(MEM_stage_inst_dmem_ram_2253), .A2(MEM_stage_inst_dmem_n36), .ZN(MEM_stage_inst_dmem_n7192) );
NAND2_X1 MEM_stage_inst_dmem_U7325 ( .A1(MEM_stage_inst_dmem_ram_3021), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n7193) );
NAND2_X1 MEM_stage_inst_dmem_U7324 ( .A1(MEM_stage_inst_dmem_n7191), .A2(MEM_stage_inst_dmem_n7190), .ZN(MEM_stage_inst_dmem_n7195) );
NAND2_X1 MEM_stage_inst_dmem_U7323 ( .A1(MEM_stage_inst_dmem_ram_2381), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n7190) );
NAND2_X1 MEM_stage_inst_dmem_U7322 ( .A1(MEM_stage_inst_dmem_ram_2973), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n7191) );
NOR2_X1 MEM_stage_inst_dmem_U7321 ( .A1(MEM_stage_inst_dmem_n7189), .A2(MEM_stage_inst_dmem_n7188), .ZN(MEM_stage_inst_dmem_n7197) );
NAND2_X1 MEM_stage_inst_dmem_U7320 ( .A1(MEM_stage_inst_dmem_n7187), .A2(MEM_stage_inst_dmem_n7186), .ZN(MEM_stage_inst_dmem_n7188) );
NAND2_X1 MEM_stage_inst_dmem_U7319 ( .A1(MEM_stage_inst_dmem_ram_2621), .A2(MEM_stage_inst_dmem_n41), .ZN(MEM_stage_inst_dmem_n7186) );
NAND2_X1 MEM_stage_inst_dmem_U7318 ( .A1(MEM_stage_inst_dmem_ram_2189), .A2(MEM_stage_inst_dmem_n61), .ZN(MEM_stage_inst_dmem_n7187) );
NAND2_X1 MEM_stage_inst_dmem_U7317 ( .A1(MEM_stage_inst_dmem_n7185), .A2(MEM_stage_inst_dmem_n7184), .ZN(MEM_stage_inst_dmem_n7189) );
NAND2_X1 MEM_stage_inst_dmem_U7316 ( .A1(MEM_stage_inst_dmem_ram_2477), .A2(MEM_stage_inst_dmem_n4772), .ZN(MEM_stage_inst_dmem_n7184) );
NAND2_X1 MEM_stage_inst_dmem_U7315 ( .A1(MEM_stage_inst_dmem_ram_3037), .A2(MEM_stage_inst_dmem_n7895), .ZN(MEM_stage_inst_dmem_n7185) );
NAND2_X1 MEM_stage_inst_dmem_U7314 ( .A1(MEM_stage_inst_dmem_n7183), .A2(MEM_stage_inst_dmem_n7182), .ZN(MEM_stage_inst_dmem_n7199) );
NOR2_X1 MEM_stage_inst_dmem_U7313 ( .A1(MEM_stage_inst_dmem_n7181), .A2(MEM_stage_inst_dmem_n7180), .ZN(MEM_stage_inst_dmem_n7182) );
NAND2_X1 MEM_stage_inst_dmem_U7312 ( .A1(MEM_stage_inst_dmem_n7179), .A2(MEM_stage_inst_dmem_n7178), .ZN(MEM_stage_inst_dmem_n7180) );
NAND2_X1 MEM_stage_inst_dmem_U7311 ( .A1(MEM_stage_inst_dmem_ram_2413), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n7178) );
NAND2_X1 MEM_stage_inst_dmem_U7310 ( .A1(MEM_stage_inst_dmem_ram_2701), .A2(MEM_stage_inst_dmem_n7960), .ZN(MEM_stage_inst_dmem_n7179) );
NAND2_X1 MEM_stage_inst_dmem_U7309 ( .A1(MEM_stage_inst_dmem_n7177), .A2(MEM_stage_inst_dmem_n7176), .ZN(MEM_stage_inst_dmem_n7181) );
NAND2_X1 MEM_stage_inst_dmem_U7308 ( .A1(MEM_stage_inst_dmem_ram_2285), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n7176) );
NAND2_X1 MEM_stage_inst_dmem_U7307 ( .A1(MEM_stage_inst_dmem_ram_2397), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n7177) );
NOR2_X1 MEM_stage_inst_dmem_U7306 ( .A1(MEM_stage_inst_dmem_n7175), .A2(MEM_stage_inst_dmem_n7174), .ZN(MEM_stage_inst_dmem_n7183) );
NAND2_X1 MEM_stage_inst_dmem_U7305 ( .A1(MEM_stage_inst_dmem_n7173), .A2(MEM_stage_inst_dmem_n7172), .ZN(MEM_stage_inst_dmem_n7174) );
NAND2_X1 MEM_stage_inst_dmem_U7304 ( .A1(MEM_stage_inst_dmem_ram_2061), .A2(MEM_stage_inst_dmem_n7953), .ZN(MEM_stage_inst_dmem_n7172) );
NAND2_X1 MEM_stage_inst_dmem_U7303 ( .A1(MEM_stage_inst_dmem_ram_2717), .A2(MEM_stage_inst_dmem_n3076), .ZN(MEM_stage_inst_dmem_n7173) );
NAND2_X1 MEM_stage_inst_dmem_U7302 ( .A1(MEM_stage_inst_dmem_n7171), .A2(MEM_stage_inst_dmem_n7170), .ZN(MEM_stage_inst_dmem_n7175) );
NAND2_X1 MEM_stage_inst_dmem_U7301 ( .A1(MEM_stage_inst_dmem_ram_2909), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n7170) );
NAND2_X1 MEM_stage_inst_dmem_U7300 ( .A1(MEM_stage_inst_dmem_ram_2781), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n7171) );
NAND2_X1 MEM_stage_inst_dmem_U7299 ( .A1(MEM_stage_inst_dmem_n7169), .A2(MEM_stage_inst_dmem_n7168), .ZN(MEM_stage_inst_dmem_n7233) );
NOR2_X1 MEM_stage_inst_dmem_U7298 ( .A1(MEM_stage_inst_dmem_n7167), .A2(MEM_stage_inst_dmem_n7166), .ZN(MEM_stage_inst_dmem_n7168) );
NAND2_X1 MEM_stage_inst_dmem_U7297 ( .A1(MEM_stage_inst_dmem_n7165), .A2(MEM_stage_inst_dmem_n7164), .ZN(MEM_stage_inst_dmem_n7166) );
NOR2_X1 MEM_stage_inst_dmem_U7296 ( .A1(MEM_stage_inst_dmem_n7163), .A2(MEM_stage_inst_dmem_n7162), .ZN(MEM_stage_inst_dmem_n7164) );
NAND2_X1 MEM_stage_inst_dmem_U7295 ( .A1(MEM_stage_inst_dmem_n7161), .A2(MEM_stage_inst_dmem_n7160), .ZN(MEM_stage_inst_dmem_n7162) );
NAND2_X1 MEM_stage_inst_dmem_U7294 ( .A1(MEM_stage_inst_dmem_ram_2957), .A2(MEM_stage_inst_dmem_n72), .ZN(MEM_stage_inst_dmem_n7160) );
NAND2_X1 MEM_stage_inst_dmem_U7293 ( .A1(MEM_stage_inst_dmem_ram_2077), .A2(MEM_stage_inst_dmem_n7887), .ZN(MEM_stage_inst_dmem_n7161) );
NAND2_X1 MEM_stage_inst_dmem_U7292 ( .A1(MEM_stage_inst_dmem_n7159), .A2(MEM_stage_inst_dmem_n7158), .ZN(MEM_stage_inst_dmem_n7163) );
NAND2_X1 MEM_stage_inst_dmem_U7291 ( .A1(MEM_stage_inst_dmem_ram_2557), .A2(MEM_stage_inst_dmem_n8535), .ZN(MEM_stage_inst_dmem_n7158) );
NAND2_X1 MEM_stage_inst_dmem_U7290 ( .A1(MEM_stage_inst_dmem_ram_2237), .A2(MEM_stage_inst_dmem_n7937), .ZN(MEM_stage_inst_dmem_n7159) );
NOR2_X1 MEM_stage_inst_dmem_U7289 ( .A1(MEM_stage_inst_dmem_n7157), .A2(MEM_stage_inst_dmem_n7156), .ZN(MEM_stage_inst_dmem_n7165) );
NAND2_X1 MEM_stage_inst_dmem_U7288 ( .A1(MEM_stage_inst_dmem_n7155), .A2(MEM_stage_inst_dmem_n7154), .ZN(MEM_stage_inst_dmem_n7156) );
NAND2_X1 MEM_stage_inst_dmem_U7287 ( .A1(MEM_stage_inst_dmem_ram_2941), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n7154) );
NAND2_X1 MEM_stage_inst_dmem_U7286 ( .A1(MEM_stage_inst_dmem_ram_3053), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n7155) );
NAND2_X1 MEM_stage_inst_dmem_U7285 ( .A1(MEM_stage_inst_dmem_n7153), .A2(MEM_stage_inst_dmem_n7152), .ZN(MEM_stage_inst_dmem_n7157) );
NAND2_X1 MEM_stage_inst_dmem_U7284 ( .A1(MEM_stage_inst_dmem_ram_2109), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n7152) );
NAND2_X1 MEM_stage_inst_dmem_U7283 ( .A1(MEM_stage_inst_dmem_ram_2989), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n7153) );
NAND2_X1 MEM_stage_inst_dmem_U7282 ( .A1(MEM_stage_inst_dmem_n7151), .A2(MEM_stage_inst_dmem_n7150), .ZN(MEM_stage_inst_dmem_n7167) );
NOR2_X1 MEM_stage_inst_dmem_U7281 ( .A1(MEM_stage_inst_dmem_n7149), .A2(MEM_stage_inst_dmem_n7148), .ZN(MEM_stage_inst_dmem_n7150) );
NAND2_X1 MEM_stage_inst_dmem_U7280 ( .A1(MEM_stage_inst_dmem_n7147), .A2(MEM_stage_inst_dmem_n7146), .ZN(MEM_stage_inst_dmem_n7148) );
NAND2_X1 MEM_stage_inst_dmem_U7279 ( .A1(MEM_stage_inst_dmem_ram_2365), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n7146) );
NAND2_X1 MEM_stage_inst_dmem_U7278 ( .A1(MEM_stage_inst_dmem_ram_2573), .A2(MEM_stage_inst_dmem_n71), .ZN(MEM_stage_inst_dmem_n7147) );
NAND2_X1 MEM_stage_inst_dmem_U7277 ( .A1(MEM_stage_inst_dmem_n7145), .A2(MEM_stage_inst_dmem_n7144), .ZN(MEM_stage_inst_dmem_n7149) );
NAND2_X1 MEM_stage_inst_dmem_U7276 ( .A1(MEM_stage_inst_dmem_ram_2925), .A2(MEM_stage_inst_dmem_n7923), .ZN(MEM_stage_inst_dmem_n7144) );
NAND2_X1 MEM_stage_inst_dmem_U7275 ( .A1(MEM_stage_inst_dmem_ram_2141), .A2(MEM_stage_inst_dmem_n7938), .ZN(MEM_stage_inst_dmem_n7145) );
NOR2_X1 MEM_stage_inst_dmem_U7274 ( .A1(MEM_stage_inst_dmem_n7143), .A2(MEM_stage_inst_dmem_n7142), .ZN(MEM_stage_inst_dmem_n7151) );
NAND2_X1 MEM_stage_inst_dmem_U7273 ( .A1(MEM_stage_inst_dmem_n7141), .A2(MEM_stage_inst_dmem_n7140), .ZN(MEM_stage_inst_dmem_n7142) );
NAND2_X1 MEM_stage_inst_dmem_U7272 ( .A1(MEM_stage_inst_dmem_ram_2525), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n7140) );
NAND2_X1 MEM_stage_inst_dmem_U7271 ( .A1(MEM_stage_inst_dmem_ram_2429), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n7141) );
NAND2_X1 MEM_stage_inst_dmem_U7270 ( .A1(MEM_stage_inst_dmem_n7139), .A2(MEM_stage_inst_dmem_n7138), .ZN(MEM_stage_inst_dmem_n7143) );
NAND2_X1 MEM_stage_inst_dmem_U7269 ( .A1(MEM_stage_inst_dmem_ram_2605), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n7138) );
NAND2_X1 MEM_stage_inst_dmem_U7268 ( .A1(MEM_stage_inst_dmem_ram_2205), .A2(MEM_stage_inst_dmem_n7903), .ZN(MEM_stage_inst_dmem_n7139) );
NOR2_X1 MEM_stage_inst_dmem_U7267 ( .A1(MEM_stage_inst_dmem_n7137), .A2(MEM_stage_inst_dmem_n7136), .ZN(MEM_stage_inst_dmem_n7169) );
NAND2_X1 MEM_stage_inst_dmem_U7266 ( .A1(MEM_stage_inst_dmem_n7135), .A2(MEM_stage_inst_dmem_n7134), .ZN(MEM_stage_inst_dmem_n7136) );
NOR2_X1 MEM_stage_inst_dmem_U7265 ( .A1(MEM_stage_inst_dmem_n7133), .A2(MEM_stage_inst_dmem_n7132), .ZN(MEM_stage_inst_dmem_n7134) );
NAND2_X1 MEM_stage_inst_dmem_U7264 ( .A1(MEM_stage_inst_dmem_n7131), .A2(MEM_stage_inst_dmem_n7130), .ZN(MEM_stage_inst_dmem_n7132) );
NAND2_X1 MEM_stage_inst_dmem_U7263 ( .A1(MEM_stage_inst_dmem_ram_2893), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n7130) );
NAND2_X1 MEM_stage_inst_dmem_U7262 ( .A1(MEM_stage_inst_dmem_ram_3005), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n7131) );
NAND2_X1 MEM_stage_inst_dmem_U7261 ( .A1(MEM_stage_inst_dmem_n7129), .A2(MEM_stage_inst_dmem_n7128), .ZN(MEM_stage_inst_dmem_n7133) );
NAND2_X1 MEM_stage_inst_dmem_U7260 ( .A1(MEM_stage_inst_dmem_ram_2813), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n7128) );
NAND2_X1 MEM_stage_inst_dmem_U7259 ( .A1(MEM_stage_inst_dmem_ram_2733), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n7129) );
NOR2_X1 MEM_stage_inst_dmem_U7258 ( .A1(MEM_stage_inst_dmem_n7127), .A2(MEM_stage_inst_dmem_n7126), .ZN(MEM_stage_inst_dmem_n7135) );
NAND2_X1 MEM_stage_inst_dmem_U7257 ( .A1(MEM_stage_inst_dmem_n7125), .A2(MEM_stage_inst_dmem_n7124), .ZN(MEM_stage_inst_dmem_n7126) );
NAND2_X1 MEM_stage_inst_dmem_U7256 ( .A1(MEM_stage_inst_dmem_ram_2349), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n7124) );
NAND2_X1 MEM_stage_inst_dmem_U7255 ( .A1(MEM_stage_inst_dmem_ram_2797), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n7125) );
NAND2_X1 MEM_stage_inst_dmem_U7254 ( .A1(MEM_stage_inst_dmem_n7123), .A2(MEM_stage_inst_dmem_n7122), .ZN(MEM_stage_inst_dmem_n7127) );
NAND2_X1 MEM_stage_inst_dmem_U7253 ( .A1(MEM_stage_inst_dmem_ram_2541), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n7122) );
NAND2_X1 MEM_stage_inst_dmem_U7252 ( .A1(MEM_stage_inst_dmem_ram_2093), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n7123) );
NAND2_X1 MEM_stage_inst_dmem_U7251 ( .A1(MEM_stage_inst_dmem_n7121), .A2(MEM_stage_inst_dmem_n7120), .ZN(MEM_stage_inst_dmem_n7137) );
NOR2_X1 MEM_stage_inst_dmem_U7250 ( .A1(MEM_stage_inst_dmem_n7119), .A2(MEM_stage_inst_dmem_n7118), .ZN(MEM_stage_inst_dmem_n7120) );
NAND2_X1 MEM_stage_inst_dmem_U7249 ( .A1(MEM_stage_inst_dmem_n7117), .A2(MEM_stage_inst_dmem_n7116), .ZN(MEM_stage_inst_dmem_n7118) );
NAND2_X1 MEM_stage_inst_dmem_U7248 ( .A1(MEM_stage_inst_dmem_ram_2493), .A2(MEM_stage_inst_dmem_n7888), .ZN(MEM_stage_inst_dmem_n7116) );
NAND2_X1 MEM_stage_inst_dmem_U7247 ( .A1(MEM_stage_inst_dmem_ram_2509), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n7117) );
NAND2_X1 MEM_stage_inst_dmem_U7246 ( .A1(MEM_stage_inst_dmem_n7115), .A2(MEM_stage_inst_dmem_n7114), .ZN(MEM_stage_inst_dmem_n7119) );
NAND2_X1 MEM_stage_inst_dmem_U7245 ( .A1(MEM_stage_inst_dmem_ram_2765), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n7114) );
NAND2_X1 MEM_stage_inst_dmem_U7244 ( .A1(MEM_stage_inst_dmem_ram_2157), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n7115) );
NOR2_X1 MEM_stage_inst_dmem_U7243 ( .A1(MEM_stage_inst_dmem_n7113), .A2(MEM_stage_inst_dmem_n7112), .ZN(MEM_stage_inst_dmem_n7121) );
NAND2_X1 MEM_stage_inst_dmem_U7242 ( .A1(MEM_stage_inst_dmem_n7111), .A2(MEM_stage_inst_dmem_n7110), .ZN(MEM_stage_inst_dmem_n7112) );
NAND2_X1 MEM_stage_inst_dmem_U7241 ( .A1(MEM_stage_inst_dmem_ram_2125), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n7110) );
NAND2_X1 MEM_stage_inst_dmem_U7240 ( .A1(MEM_stage_inst_dmem_ram_2445), .A2(MEM_stage_inst_dmem_n7930), .ZN(MEM_stage_inst_dmem_n7111) );
NAND2_X1 MEM_stage_inst_dmem_U7239 ( .A1(MEM_stage_inst_dmem_n7109), .A2(MEM_stage_inst_dmem_n7108), .ZN(MEM_stage_inst_dmem_n7113) );
NAND2_X1 MEM_stage_inst_dmem_U7238 ( .A1(MEM_stage_inst_dmem_ram_2461), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n7108) );
NAND2_X1 MEM_stage_inst_dmem_U7237 ( .A1(MEM_stage_inst_dmem_ram_2653), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n7109) );
NOR2_X1 MEM_stage_inst_dmem_U7236 ( .A1(MEM_stage_inst_dmem_n7107), .A2(MEM_stage_inst_dmem_n8417), .ZN(MEM_stage_inst_dmem_n7236) );
NOR2_X1 MEM_stage_inst_dmem_U7235 ( .A1(MEM_stage_inst_dmem_n7106), .A2(MEM_stage_inst_dmem_n7105), .ZN(MEM_stage_inst_dmem_n7107) );
NAND2_X1 MEM_stage_inst_dmem_U7234 ( .A1(MEM_stage_inst_dmem_n7104), .A2(MEM_stage_inst_dmem_n7103), .ZN(MEM_stage_inst_dmem_n7105) );
NOR2_X1 MEM_stage_inst_dmem_U7233 ( .A1(MEM_stage_inst_dmem_n7102), .A2(MEM_stage_inst_dmem_n7101), .ZN(MEM_stage_inst_dmem_n7103) );
NAND2_X1 MEM_stage_inst_dmem_U7232 ( .A1(MEM_stage_inst_dmem_n7100), .A2(MEM_stage_inst_dmem_n7099), .ZN(MEM_stage_inst_dmem_n7101) );
NOR2_X1 MEM_stage_inst_dmem_U7231 ( .A1(MEM_stage_inst_dmem_n7098), .A2(MEM_stage_inst_dmem_n7097), .ZN(MEM_stage_inst_dmem_n7099) );
NAND2_X1 MEM_stage_inst_dmem_U7230 ( .A1(MEM_stage_inst_dmem_n7096), .A2(MEM_stage_inst_dmem_n7095), .ZN(MEM_stage_inst_dmem_n7097) );
NAND2_X1 MEM_stage_inst_dmem_U7229 ( .A1(MEM_stage_inst_dmem_ram_4013), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n7095) );
NAND2_X1 MEM_stage_inst_dmem_U7228 ( .A1(MEM_stage_inst_dmem_ram_3805), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n7096) );
NAND2_X1 MEM_stage_inst_dmem_U7227 ( .A1(MEM_stage_inst_dmem_n7094), .A2(MEM_stage_inst_dmem_n7093), .ZN(MEM_stage_inst_dmem_n7098) );
NAND2_X1 MEM_stage_inst_dmem_U7226 ( .A1(MEM_stage_inst_dmem_ram_3277), .A2(MEM_stage_inst_dmem_n36), .ZN(MEM_stage_inst_dmem_n7093) );
NAND2_X1 MEM_stage_inst_dmem_U7225 ( .A1(MEM_stage_inst_dmem_ram_3933), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n7094) );
NOR2_X1 MEM_stage_inst_dmem_U7224 ( .A1(MEM_stage_inst_dmem_n7092), .A2(MEM_stage_inst_dmem_n7091), .ZN(MEM_stage_inst_dmem_n7100) );
NAND2_X1 MEM_stage_inst_dmem_U7223 ( .A1(MEM_stage_inst_dmem_n7090), .A2(MEM_stage_inst_dmem_n7089), .ZN(MEM_stage_inst_dmem_n7091) );
NAND2_X1 MEM_stage_inst_dmem_U7222 ( .A1(MEM_stage_inst_dmem_ram_3965), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n7089) );
NAND2_X1 MEM_stage_inst_dmem_U7221 ( .A1(MEM_stage_inst_dmem_ram_4045), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n7090) );
NAND2_X1 MEM_stage_inst_dmem_U7220 ( .A1(MEM_stage_inst_dmem_n7088), .A2(MEM_stage_inst_dmem_n7087), .ZN(MEM_stage_inst_dmem_n7092) );
NAND2_X1 MEM_stage_inst_dmem_U7219 ( .A1(MEM_stage_inst_dmem_ram_3517), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n7087) );
NAND2_X1 MEM_stage_inst_dmem_U7218 ( .A1(MEM_stage_inst_dmem_ram_3437), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n7088) );
NAND2_X1 MEM_stage_inst_dmem_U7217 ( .A1(MEM_stage_inst_dmem_n7086), .A2(MEM_stage_inst_dmem_n7085), .ZN(MEM_stage_inst_dmem_n7102) );
NOR2_X1 MEM_stage_inst_dmem_U7216 ( .A1(MEM_stage_inst_dmem_n7084), .A2(MEM_stage_inst_dmem_n7083), .ZN(MEM_stage_inst_dmem_n7085) );
NAND2_X1 MEM_stage_inst_dmem_U7215 ( .A1(MEM_stage_inst_dmem_n7082), .A2(MEM_stage_inst_dmem_n7081), .ZN(MEM_stage_inst_dmem_n7083) );
NAND2_X1 MEM_stage_inst_dmem_U7214 ( .A1(MEM_stage_inst_dmem_ram_3117), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n7081) );
NAND2_X1 MEM_stage_inst_dmem_U7213 ( .A1(MEM_stage_inst_dmem_ram_3885), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n7082) );
NAND2_X1 MEM_stage_inst_dmem_U7212 ( .A1(MEM_stage_inst_dmem_n7080), .A2(MEM_stage_inst_dmem_n7079), .ZN(MEM_stage_inst_dmem_n7084) );
NAND2_X1 MEM_stage_inst_dmem_U7211 ( .A1(MEM_stage_inst_dmem_ram_3133), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n7079) );
NAND2_X1 MEM_stage_inst_dmem_U7210 ( .A1(MEM_stage_inst_dmem_ram_3981), .A2(MEM_stage_inst_dmem_n72), .ZN(MEM_stage_inst_dmem_n7080) );
NOR2_X1 MEM_stage_inst_dmem_U7209 ( .A1(MEM_stage_inst_dmem_n7078), .A2(MEM_stage_inst_dmem_n7077), .ZN(MEM_stage_inst_dmem_n7086) );
NAND2_X1 MEM_stage_inst_dmem_U7208 ( .A1(MEM_stage_inst_dmem_n7076), .A2(MEM_stage_inst_dmem_n7075), .ZN(MEM_stage_inst_dmem_n7077) );
NAND2_X1 MEM_stage_inst_dmem_U7207 ( .A1(MEM_stage_inst_dmem_ram_4077), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n7075) );
NAND2_X1 MEM_stage_inst_dmem_U7206 ( .A1(MEM_stage_inst_dmem_ram_3533), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n7076) );
NAND2_X1 MEM_stage_inst_dmem_U7205 ( .A1(MEM_stage_inst_dmem_n7074), .A2(MEM_stage_inst_dmem_n7073), .ZN(MEM_stage_inst_dmem_n7078) );
NAND2_X1 MEM_stage_inst_dmem_U7204 ( .A1(MEM_stage_inst_dmem_ram_3917), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n7073) );
NAND2_X1 MEM_stage_inst_dmem_U7203 ( .A1(MEM_stage_inst_dmem_ram_3213), .A2(MEM_stage_inst_dmem_n61), .ZN(MEM_stage_inst_dmem_n7074) );
NOR2_X1 MEM_stage_inst_dmem_U7202 ( .A1(MEM_stage_inst_dmem_n7072), .A2(MEM_stage_inst_dmem_n7071), .ZN(MEM_stage_inst_dmem_n7104) );
NAND2_X1 MEM_stage_inst_dmem_U7201 ( .A1(MEM_stage_inst_dmem_n7070), .A2(MEM_stage_inst_dmem_n7069), .ZN(MEM_stage_inst_dmem_n7071) );
NOR2_X1 MEM_stage_inst_dmem_U7200 ( .A1(MEM_stage_inst_dmem_n7068), .A2(MEM_stage_inst_dmem_n7067), .ZN(MEM_stage_inst_dmem_n7069) );
NAND2_X1 MEM_stage_inst_dmem_U7199 ( .A1(MEM_stage_inst_dmem_n7066), .A2(MEM_stage_inst_dmem_n7065), .ZN(MEM_stage_inst_dmem_n7067) );
NAND2_X1 MEM_stage_inst_dmem_U7198 ( .A1(MEM_stage_inst_dmem_ram_3485), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n7065) );
NAND2_X1 MEM_stage_inst_dmem_U7197 ( .A1(MEM_stage_inst_dmem_ram_3101), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n7066) );
NAND2_X1 MEM_stage_inst_dmem_U7196 ( .A1(MEM_stage_inst_dmem_n7064), .A2(MEM_stage_inst_dmem_n7063), .ZN(MEM_stage_inst_dmem_n7068) );
NAND2_X1 MEM_stage_inst_dmem_U7195 ( .A1(MEM_stage_inst_dmem_ram_3309), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n7063) );
NAND2_X1 MEM_stage_inst_dmem_U7194 ( .A1(MEM_stage_inst_dmem_ram_3821), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n7064) );
NOR2_X1 MEM_stage_inst_dmem_U7193 ( .A1(MEM_stage_inst_dmem_n7062), .A2(MEM_stage_inst_dmem_n7061), .ZN(MEM_stage_inst_dmem_n7070) );
NAND2_X1 MEM_stage_inst_dmem_U7192 ( .A1(MEM_stage_inst_dmem_n7060), .A2(MEM_stage_inst_dmem_n7059), .ZN(MEM_stage_inst_dmem_n7061) );
NAND2_X1 MEM_stage_inst_dmem_U7191 ( .A1(MEM_stage_inst_dmem_ram_3405), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n7059) );
NAND2_X1 MEM_stage_inst_dmem_U7190 ( .A1(MEM_stage_inst_dmem_ram_3469), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n7060) );
NAND2_X1 MEM_stage_inst_dmem_U7189 ( .A1(MEM_stage_inst_dmem_n7058), .A2(MEM_stage_inst_dmem_n7057), .ZN(MEM_stage_inst_dmem_n7062) );
NAND2_X1 MEM_stage_inst_dmem_U7188 ( .A1(MEM_stage_inst_dmem_ram_3693), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n7057) );
NAND2_X1 MEM_stage_inst_dmem_U7187 ( .A1(MEM_stage_inst_dmem_ram_3261), .A2(MEM_stage_inst_dmem_n8434), .ZN(MEM_stage_inst_dmem_n7058) );
NAND2_X1 MEM_stage_inst_dmem_U7186 ( .A1(MEM_stage_inst_dmem_n7056), .A2(MEM_stage_inst_dmem_n7055), .ZN(MEM_stage_inst_dmem_n7072) );
NOR2_X1 MEM_stage_inst_dmem_U7185 ( .A1(MEM_stage_inst_dmem_n7054), .A2(MEM_stage_inst_dmem_n7053), .ZN(MEM_stage_inst_dmem_n7055) );
NAND2_X1 MEM_stage_inst_dmem_U7184 ( .A1(MEM_stage_inst_dmem_n7052), .A2(MEM_stage_inst_dmem_n7051), .ZN(MEM_stage_inst_dmem_n7053) );
NAND2_X1 MEM_stage_inst_dmem_U7183 ( .A1(MEM_stage_inst_dmem_ram_3549), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n7051) );
NAND2_X1 MEM_stage_inst_dmem_U7182 ( .A1(MEM_stage_inst_dmem_ram_3709), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n7052) );
NAND2_X1 MEM_stage_inst_dmem_U7181 ( .A1(MEM_stage_inst_dmem_n7050), .A2(MEM_stage_inst_dmem_n7049), .ZN(MEM_stage_inst_dmem_n7054) );
NAND2_X1 MEM_stage_inst_dmem_U7180 ( .A1(MEM_stage_inst_dmem_ram_3757), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n7049) );
NAND2_X1 MEM_stage_inst_dmem_U7179 ( .A1(MEM_stage_inst_dmem_ram_3181), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n7050) );
NOR2_X1 MEM_stage_inst_dmem_U7178 ( .A1(MEM_stage_inst_dmem_n7048), .A2(MEM_stage_inst_dmem_n7047), .ZN(MEM_stage_inst_dmem_n7056) );
NAND2_X1 MEM_stage_inst_dmem_U7177 ( .A1(MEM_stage_inst_dmem_n7046), .A2(MEM_stage_inst_dmem_n7045), .ZN(MEM_stage_inst_dmem_n7047) );
NAND2_X1 MEM_stage_inst_dmem_U7176 ( .A1(MEM_stage_inst_dmem_ram_3149), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n7045) );
NAND2_X1 MEM_stage_inst_dmem_U7175 ( .A1(MEM_stage_inst_dmem_ram_4093), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n7046) );
NAND2_X1 MEM_stage_inst_dmem_U7174 ( .A1(MEM_stage_inst_dmem_n7044), .A2(MEM_stage_inst_dmem_n7043), .ZN(MEM_stage_inst_dmem_n7048) );
NAND2_X1 MEM_stage_inst_dmem_U7173 ( .A1(MEM_stage_inst_dmem_ram_3773), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n7043) );
NAND2_X1 MEM_stage_inst_dmem_U7172 ( .A1(MEM_stage_inst_dmem_ram_3613), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n7044) );
NAND2_X1 MEM_stage_inst_dmem_U7171 ( .A1(MEM_stage_inst_dmem_n7042), .A2(MEM_stage_inst_dmem_n7041), .ZN(MEM_stage_inst_dmem_n7106) );
NOR2_X1 MEM_stage_inst_dmem_U7170 ( .A1(MEM_stage_inst_dmem_n7040), .A2(MEM_stage_inst_dmem_n7039), .ZN(MEM_stage_inst_dmem_n7041) );
NAND2_X1 MEM_stage_inst_dmem_U7169 ( .A1(MEM_stage_inst_dmem_n7038), .A2(MEM_stage_inst_dmem_n7037), .ZN(MEM_stage_inst_dmem_n7039) );
NOR2_X1 MEM_stage_inst_dmem_U7168 ( .A1(MEM_stage_inst_dmem_n7036), .A2(MEM_stage_inst_dmem_n7035), .ZN(MEM_stage_inst_dmem_n7037) );
NAND2_X1 MEM_stage_inst_dmem_U7167 ( .A1(MEM_stage_inst_dmem_n7034), .A2(MEM_stage_inst_dmem_n7033), .ZN(MEM_stage_inst_dmem_n7035) );
NAND2_X1 MEM_stage_inst_dmem_U7166 ( .A1(MEM_stage_inst_dmem_ram_3389), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n7033) );
NAND2_X1 MEM_stage_inst_dmem_U7165 ( .A1(MEM_stage_inst_dmem_ram_3421), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n7034) );
NAND2_X1 MEM_stage_inst_dmem_U7164 ( .A1(MEM_stage_inst_dmem_n7032), .A2(MEM_stage_inst_dmem_n7031), .ZN(MEM_stage_inst_dmem_n7036) );
NAND2_X1 MEM_stage_inst_dmem_U7163 ( .A1(MEM_stage_inst_dmem_ram_3325), .A2(MEM_stage_inst_dmem_n7914), .ZN(MEM_stage_inst_dmem_n7031) );
NAND2_X1 MEM_stage_inst_dmem_U7162 ( .A1(MEM_stage_inst_dmem_ram_3341), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n7032) );
NOR2_X1 MEM_stage_inst_dmem_U7161 ( .A1(MEM_stage_inst_dmem_n7030), .A2(MEM_stage_inst_dmem_n7029), .ZN(MEM_stage_inst_dmem_n7038) );
NAND2_X1 MEM_stage_inst_dmem_U7160 ( .A1(MEM_stage_inst_dmem_n7028), .A2(MEM_stage_inst_dmem_n7027), .ZN(MEM_stage_inst_dmem_n7029) );
NAND2_X1 MEM_stage_inst_dmem_U7159 ( .A1(MEM_stage_inst_dmem_ram_3949), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n7027) );
NAND2_X1 MEM_stage_inst_dmem_U7158 ( .A1(MEM_stage_inst_dmem_ram_3869), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n7028) );
NAND2_X1 MEM_stage_inst_dmem_U7157 ( .A1(MEM_stage_inst_dmem_n7026), .A2(MEM_stage_inst_dmem_n7025), .ZN(MEM_stage_inst_dmem_n7030) );
NAND2_X1 MEM_stage_inst_dmem_U7156 ( .A1(MEM_stage_inst_dmem_ram_4029), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n7025) );
NAND2_X1 MEM_stage_inst_dmem_U7155 ( .A1(MEM_stage_inst_dmem_ram_3597), .A2(MEM_stage_inst_dmem_n71), .ZN(MEM_stage_inst_dmem_n7026) );
NAND2_X1 MEM_stage_inst_dmem_U7154 ( .A1(MEM_stage_inst_dmem_n7024), .A2(MEM_stage_inst_dmem_n7023), .ZN(MEM_stage_inst_dmem_n7040) );
NOR2_X1 MEM_stage_inst_dmem_U7153 ( .A1(MEM_stage_inst_dmem_n7022), .A2(MEM_stage_inst_dmem_n7021), .ZN(MEM_stage_inst_dmem_n7023) );
NAND2_X1 MEM_stage_inst_dmem_U7152 ( .A1(MEM_stage_inst_dmem_n7020), .A2(MEM_stage_inst_dmem_n7019), .ZN(MEM_stage_inst_dmem_n7021) );
NAND2_X1 MEM_stage_inst_dmem_U7151 ( .A1(MEM_stage_inst_dmem_ram_3997), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n7019) );
NAND2_X1 MEM_stage_inst_dmem_U7150 ( .A1(MEM_stage_inst_dmem_ram_3357), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n7020) );
NAND2_X1 MEM_stage_inst_dmem_U7149 ( .A1(MEM_stage_inst_dmem_n7018), .A2(MEM_stage_inst_dmem_n7017), .ZN(MEM_stage_inst_dmem_n7022) );
NAND2_X1 MEM_stage_inst_dmem_U7148 ( .A1(MEM_stage_inst_dmem_ram_3789), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n7017) );
NAND2_X1 MEM_stage_inst_dmem_U7147 ( .A1(MEM_stage_inst_dmem_ram_3629), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n7018) );
NOR2_X1 MEM_stage_inst_dmem_U7146 ( .A1(MEM_stage_inst_dmem_n7016), .A2(MEM_stage_inst_dmem_n7015), .ZN(MEM_stage_inst_dmem_n7024) );
NAND2_X1 MEM_stage_inst_dmem_U7145 ( .A1(MEM_stage_inst_dmem_n7014), .A2(MEM_stage_inst_dmem_n7013), .ZN(MEM_stage_inst_dmem_n7015) );
NAND2_X1 MEM_stage_inst_dmem_U7144 ( .A1(MEM_stage_inst_dmem_ram_3245), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n7013) );
NAND2_X1 MEM_stage_inst_dmem_U7143 ( .A1(MEM_stage_inst_dmem_ram_3085), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n7014) );
NAND2_X1 MEM_stage_inst_dmem_U7142 ( .A1(MEM_stage_inst_dmem_n7012), .A2(MEM_stage_inst_dmem_n7011), .ZN(MEM_stage_inst_dmem_n7016) );
NAND2_X1 MEM_stage_inst_dmem_U7141 ( .A1(MEM_stage_inst_dmem_ram_3229), .A2(MEM_stage_inst_dmem_n44), .ZN(MEM_stage_inst_dmem_n7011) );
NAND2_X1 MEM_stage_inst_dmem_U7140 ( .A1(MEM_stage_inst_dmem_ram_3741), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n7012) );
NOR2_X1 MEM_stage_inst_dmem_U7139 ( .A1(MEM_stage_inst_dmem_n7010), .A2(MEM_stage_inst_dmem_n7009), .ZN(MEM_stage_inst_dmem_n7042) );
NAND2_X1 MEM_stage_inst_dmem_U7138 ( .A1(MEM_stage_inst_dmem_n7008), .A2(MEM_stage_inst_dmem_n7007), .ZN(MEM_stage_inst_dmem_n7009) );
NOR2_X1 MEM_stage_inst_dmem_U7137 ( .A1(MEM_stage_inst_dmem_n7006), .A2(MEM_stage_inst_dmem_n7005), .ZN(MEM_stage_inst_dmem_n7007) );
NAND2_X1 MEM_stage_inst_dmem_U7136 ( .A1(MEM_stage_inst_dmem_n7004), .A2(MEM_stage_inst_dmem_n7003), .ZN(MEM_stage_inst_dmem_n7005) );
NAND2_X1 MEM_stage_inst_dmem_U7135 ( .A1(MEM_stage_inst_dmem_ram_3645), .A2(MEM_stage_inst_dmem_n41), .ZN(MEM_stage_inst_dmem_n7003) );
NAND2_X1 MEM_stage_inst_dmem_U7134 ( .A1(MEM_stage_inst_dmem_ram_3453), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n7004) );
NAND2_X1 MEM_stage_inst_dmem_U7133 ( .A1(MEM_stage_inst_dmem_n7002), .A2(MEM_stage_inst_dmem_n7001), .ZN(MEM_stage_inst_dmem_n7006) );
NAND2_X1 MEM_stage_inst_dmem_U7132 ( .A1(MEM_stage_inst_dmem_ram_3853), .A2(MEM_stage_inst_dmem_n8472), .ZN(MEM_stage_inst_dmem_n7001) );
NAND2_X1 MEM_stage_inst_dmem_U7131 ( .A1(MEM_stage_inst_dmem_ram_3197), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n7002) );
NOR2_X1 MEM_stage_inst_dmem_U7130 ( .A1(MEM_stage_inst_dmem_n7000), .A2(MEM_stage_inst_dmem_n6999), .ZN(MEM_stage_inst_dmem_n7008) );
NAND2_X1 MEM_stage_inst_dmem_U7129 ( .A1(MEM_stage_inst_dmem_n6998), .A2(MEM_stage_inst_dmem_n6997), .ZN(MEM_stage_inst_dmem_n6999) );
NAND2_X1 MEM_stage_inst_dmem_U7128 ( .A1(MEM_stage_inst_dmem_ram_3165), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n6997) );
NAND2_X1 MEM_stage_inst_dmem_U7127 ( .A1(MEM_stage_inst_dmem_ram_3293), .A2(MEM_stage_inst_dmem_n51), .ZN(MEM_stage_inst_dmem_n6998) );
NAND2_X1 MEM_stage_inst_dmem_U7126 ( .A1(MEM_stage_inst_dmem_n6996), .A2(MEM_stage_inst_dmem_n6995), .ZN(MEM_stage_inst_dmem_n7000) );
NAND2_X1 MEM_stage_inst_dmem_U7125 ( .A1(MEM_stage_inst_dmem_ram_3837), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n6995) );
NAND2_X1 MEM_stage_inst_dmem_U7124 ( .A1(MEM_stage_inst_dmem_ram_3901), .A2(MEM_stage_inst_dmem_n8005), .ZN(MEM_stage_inst_dmem_n6996) );
NAND2_X1 MEM_stage_inst_dmem_U7123 ( .A1(MEM_stage_inst_dmem_n6994), .A2(MEM_stage_inst_dmem_n6993), .ZN(MEM_stage_inst_dmem_n7010) );
NOR2_X1 MEM_stage_inst_dmem_U7122 ( .A1(MEM_stage_inst_dmem_n6992), .A2(MEM_stage_inst_dmem_n6991), .ZN(MEM_stage_inst_dmem_n6993) );
NAND2_X1 MEM_stage_inst_dmem_U7121 ( .A1(MEM_stage_inst_dmem_n6990), .A2(MEM_stage_inst_dmem_n6989), .ZN(MEM_stage_inst_dmem_n6991) );
NAND2_X1 MEM_stage_inst_dmem_U7120 ( .A1(MEM_stage_inst_dmem_ram_3501), .A2(MEM_stage_inst_dmem_n4772), .ZN(MEM_stage_inst_dmem_n6989) );
NAND2_X1 MEM_stage_inst_dmem_U7119 ( .A1(MEM_stage_inst_dmem_ram_3677), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n6990) );
NAND2_X1 MEM_stage_inst_dmem_U7118 ( .A1(MEM_stage_inst_dmem_n6988), .A2(MEM_stage_inst_dmem_n6987), .ZN(MEM_stage_inst_dmem_n6992) );
NAND2_X1 MEM_stage_inst_dmem_U7117 ( .A1(MEM_stage_inst_dmem_ram_3565), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n6987) );
NAND2_X1 MEM_stage_inst_dmem_U7116 ( .A1(MEM_stage_inst_dmem_ram_3373), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n6988) );
NOR2_X1 MEM_stage_inst_dmem_U7115 ( .A1(MEM_stage_inst_dmem_n6986), .A2(MEM_stage_inst_dmem_n6985), .ZN(MEM_stage_inst_dmem_n6994) );
NAND2_X1 MEM_stage_inst_dmem_U7114 ( .A1(MEM_stage_inst_dmem_n6984), .A2(MEM_stage_inst_dmem_n6983), .ZN(MEM_stage_inst_dmem_n6985) );
NAND2_X1 MEM_stage_inst_dmem_U7113 ( .A1(MEM_stage_inst_dmem_ram_3725), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n6983) );
NAND2_X1 MEM_stage_inst_dmem_U7112 ( .A1(MEM_stage_inst_dmem_ram_4061), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n6984) );
NAND2_X1 MEM_stage_inst_dmem_U7111 ( .A1(MEM_stage_inst_dmem_n6982), .A2(MEM_stage_inst_dmem_n6981), .ZN(MEM_stage_inst_dmem_n6986) );
NAND2_X1 MEM_stage_inst_dmem_U7110 ( .A1(MEM_stage_inst_dmem_ram_3581), .A2(MEM_stage_inst_dmem_n64), .ZN(MEM_stage_inst_dmem_n6981) );
NAND2_X1 MEM_stage_inst_dmem_U7109 ( .A1(MEM_stage_inst_dmem_ram_3661), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n6982) );
NAND2_X1 MEM_stage_inst_dmem_U7108 ( .A1(MEM_stage_inst_dmem_n6980), .A2(MEM_stage_inst_dmem_n6979), .ZN(MEM_stage_inst_mem_read_data_12) );
NOR2_X1 MEM_stage_inst_dmem_U7107 ( .A1(MEM_stage_inst_dmem_n6978), .A2(MEM_stage_inst_dmem_n6977), .ZN(MEM_stage_inst_dmem_n6979) );
NOR2_X1 MEM_stage_inst_dmem_U7106 ( .A1(MEM_stage_inst_dmem_n6976), .A2(MEM_stage_inst_dmem_n8286), .ZN(MEM_stage_inst_dmem_n6977) );
NOR2_X1 MEM_stage_inst_dmem_U7105 ( .A1(MEM_stage_inst_dmem_n6975), .A2(MEM_stage_inst_dmem_n6974), .ZN(MEM_stage_inst_dmem_n6976) );
NAND2_X1 MEM_stage_inst_dmem_U7104 ( .A1(MEM_stage_inst_dmem_n6973), .A2(MEM_stage_inst_dmem_n6972), .ZN(MEM_stage_inst_dmem_n6974) );
NOR2_X1 MEM_stage_inst_dmem_U7103 ( .A1(MEM_stage_inst_dmem_n6971), .A2(MEM_stage_inst_dmem_n6970), .ZN(MEM_stage_inst_dmem_n6972) );
NAND2_X1 MEM_stage_inst_dmem_U7102 ( .A1(MEM_stage_inst_dmem_n6969), .A2(MEM_stage_inst_dmem_n6968), .ZN(MEM_stage_inst_dmem_n6970) );
NOR2_X1 MEM_stage_inst_dmem_U7101 ( .A1(MEM_stage_inst_dmem_n6967), .A2(MEM_stage_inst_dmem_n6966), .ZN(MEM_stage_inst_dmem_n6968) );
NAND2_X1 MEM_stage_inst_dmem_U7100 ( .A1(MEM_stage_inst_dmem_n6965), .A2(MEM_stage_inst_dmem_n6964), .ZN(MEM_stage_inst_dmem_n6966) );
NAND2_X1 MEM_stage_inst_dmem_U7099 ( .A1(MEM_stage_inst_dmem_ram_2476), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n6964) );
NAND2_X1 MEM_stage_inst_dmem_U7098 ( .A1(MEM_stage_inst_dmem_ram_2156), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n6965) );
NAND2_X1 MEM_stage_inst_dmem_U7097 ( .A1(MEM_stage_inst_dmem_n6963), .A2(MEM_stage_inst_dmem_n6962), .ZN(MEM_stage_inst_dmem_n6967) );
NAND2_X1 MEM_stage_inst_dmem_U7096 ( .A1(MEM_stage_inst_dmem_ram_2460), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n6962) );
NAND2_X1 MEM_stage_inst_dmem_U7095 ( .A1(MEM_stage_inst_dmem_ram_3004), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n6963) );
NOR2_X1 MEM_stage_inst_dmem_U7094 ( .A1(MEM_stage_inst_dmem_n6961), .A2(MEM_stage_inst_dmem_n6960), .ZN(MEM_stage_inst_dmem_n6969) );
NAND2_X1 MEM_stage_inst_dmem_U7093 ( .A1(MEM_stage_inst_dmem_n6959), .A2(MEM_stage_inst_dmem_n6958), .ZN(MEM_stage_inst_dmem_n6960) );
NAND2_X1 MEM_stage_inst_dmem_U7092 ( .A1(MEM_stage_inst_dmem_ram_2972), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n6958) );
NAND2_X1 MEM_stage_inst_dmem_U7091 ( .A1(MEM_stage_inst_dmem_ram_3020), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n6959) );
NAND2_X1 MEM_stage_inst_dmem_U7090 ( .A1(MEM_stage_inst_dmem_n6957), .A2(MEM_stage_inst_dmem_n6956), .ZN(MEM_stage_inst_dmem_n6961) );
NAND2_X1 MEM_stage_inst_dmem_U7089 ( .A1(MEM_stage_inst_dmem_ram_2172), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n6956) );
NAND2_X1 MEM_stage_inst_dmem_U7088 ( .A1(MEM_stage_inst_dmem_ram_2684), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n6957) );
NAND2_X1 MEM_stage_inst_dmem_U7087 ( .A1(MEM_stage_inst_dmem_n6955), .A2(MEM_stage_inst_dmem_n6954), .ZN(MEM_stage_inst_dmem_n6971) );
NOR2_X1 MEM_stage_inst_dmem_U7086 ( .A1(MEM_stage_inst_dmem_n6953), .A2(MEM_stage_inst_dmem_n6952), .ZN(MEM_stage_inst_dmem_n6954) );
NAND2_X1 MEM_stage_inst_dmem_U7085 ( .A1(MEM_stage_inst_dmem_n6951), .A2(MEM_stage_inst_dmem_n6950), .ZN(MEM_stage_inst_dmem_n6952) );
NAND2_X1 MEM_stage_inst_dmem_U7084 ( .A1(MEM_stage_inst_dmem_ram_2188), .A2(MEM_stage_inst_dmem_n8174), .ZN(MEM_stage_inst_dmem_n6950) );
NAND2_X1 MEM_stage_inst_dmem_U7083 ( .A1(MEM_stage_inst_dmem_ram_2748), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n6951) );
NAND2_X1 MEM_stage_inst_dmem_U7082 ( .A1(MEM_stage_inst_dmem_n6949), .A2(MEM_stage_inst_dmem_n6948), .ZN(MEM_stage_inst_dmem_n6953) );
NAND2_X1 MEM_stage_inst_dmem_U7081 ( .A1(MEM_stage_inst_dmem_ram_2924), .A2(MEM_stage_inst_dmem_n7923), .ZN(MEM_stage_inst_dmem_n6948) );
NAND2_X1 MEM_stage_inst_dmem_U7080 ( .A1(MEM_stage_inst_dmem_ram_2396), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n6949) );
NOR2_X1 MEM_stage_inst_dmem_U7079 ( .A1(MEM_stage_inst_dmem_n6947), .A2(MEM_stage_inst_dmem_n6946), .ZN(MEM_stage_inst_dmem_n6955) );
NAND2_X1 MEM_stage_inst_dmem_U7078 ( .A1(MEM_stage_inst_dmem_n6945), .A2(MEM_stage_inst_dmem_n6944), .ZN(MEM_stage_inst_dmem_n6946) );
NAND2_X1 MEM_stage_inst_dmem_U7077 ( .A1(MEM_stage_inst_dmem_ram_2412), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n6944) );
NAND2_X1 MEM_stage_inst_dmem_U7076 ( .A1(MEM_stage_inst_dmem_ram_2332), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n6945) );
NAND2_X1 MEM_stage_inst_dmem_U7075 ( .A1(MEM_stage_inst_dmem_n6943), .A2(MEM_stage_inst_dmem_n6942), .ZN(MEM_stage_inst_dmem_n6947) );
NAND2_X1 MEM_stage_inst_dmem_U7074 ( .A1(MEM_stage_inst_dmem_ram_2300), .A2(MEM_stage_inst_dmem_n7914), .ZN(MEM_stage_inst_dmem_n6942) );
NAND2_X1 MEM_stage_inst_dmem_U7073 ( .A1(MEM_stage_inst_dmem_ram_2876), .A2(MEM_stage_inst_dmem_n8005), .ZN(MEM_stage_inst_dmem_n6943) );
NOR2_X1 MEM_stage_inst_dmem_U7072 ( .A1(MEM_stage_inst_dmem_n6941), .A2(MEM_stage_inst_dmem_n6940), .ZN(MEM_stage_inst_dmem_n6973) );
NAND2_X1 MEM_stage_inst_dmem_U7071 ( .A1(MEM_stage_inst_dmem_n6939), .A2(MEM_stage_inst_dmem_n6938), .ZN(MEM_stage_inst_dmem_n6940) );
NOR2_X1 MEM_stage_inst_dmem_U7070 ( .A1(MEM_stage_inst_dmem_n6937), .A2(MEM_stage_inst_dmem_n6936), .ZN(MEM_stage_inst_dmem_n6938) );
NAND2_X1 MEM_stage_inst_dmem_U7069 ( .A1(MEM_stage_inst_dmem_n6935), .A2(MEM_stage_inst_dmem_n6934), .ZN(MEM_stage_inst_dmem_n6936) );
NAND2_X1 MEM_stage_inst_dmem_U7068 ( .A1(MEM_stage_inst_dmem_ram_2124), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n6934) );
NAND2_X1 MEM_stage_inst_dmem_U7067 ( .A1(MEM_stage_inst_dmem_ram_2732), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n6935) );
NAND2_X1 MEM_stage_inst_dmem_U7066 ( .A1(MEM_stage_inst_dmem_n6933), .A2(MEM_stage_inst_dmem_n6932), .ZN(MEM_stage_inst_dmem_n6937) );
NAND2_X1 MEM_stage_inst_dmem_U7065 ( .A1(MEM_stage_inst_dmem_ram_2364), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n6932) );
NAND2_X1 MEM_stage_inst_dmem_U7064 ( .A1(MEM_stage_inst_dmem_ram_2444), .A2(MEM_stage_inst_dmem_n7930), .ZN(MEM_stage_inst_dmem_n6933) );
NOR2_X1 MEM_stage_inst_dmem_U7063 ( .A1(MEM_stage_inst_dmem_n6931), .A2(MEM_stage_inst_dmem_n6930), .ZN(MEM_stage_inst_dmem_n6939) );
NAND2_X1 MEM_stage_inst_dmem_U7062 ( .A1(MEM_stage_inst_dmem_n6929), .A2(MEM_stage_inst_dmem_n6928), .ZN(MEM_stage_inst_dmem_n6930) );
NAND2_X1 MEM_stage_inst_dmem_U7061 ( .A1(MEM_stage_inst_dmem_ram_2348), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n6928) );
NAND2_X1 MEM_stage_inst_dmem_U7060 ( .A1(MEM_stage_inst_dmem_ram_2220), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n6929) );
NAND2_X1 MEM_stage_inst_dmem_U7059 ( .A1(MEM_stage_inst_dmem_n6927), .A2(MEM_stage_inst_dmem_n6926), .ZN(MEM_stage_inst_dmem_n6931) );
NAND2_X1 MEM_stage_inst_dmem_U7058 ( .A1(MEM_stage_inst_dmem_ram_2540), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n6926) );
NAND2_X1 MEM_stage_inst_dmem_U7057 ( .A1(MEM_stage_inst_dmem_ram_3036), .A2(MEM_stage_inst_dmem_n7895), .ZN(MEM_stage_inst_dmem_n6927) );
NAND2_X1 MEM_stage_inst_dmem_U7056 ( .A1(MEM_stage_inst_dmem_n6925), .A2(MEM_stage_inst_dmem_n6924), .ZN(MEM_stage_inst_dmem_n6941) );
NOR2_X1 MEM_stage_inst_dmem_U7055 ( .A1(MEM_stage_inst_dmem_n6923), .A2(MEM_stage_inst_dmem_n6922), .ZN(MEM_stage_inst_dmem_n6924) );
NAND2_X1 MEM_stage_inst_dmem_U7054 ( .A1(MEM_stage_inst_dmem_n6921), .A2(MEM_stage_inst_dmem_n6920), .ZN(MEM_stage_inst_dmem_n6922) );
NAND2_X1 MEM_stage_inst_dmem_U7053 ( .A1(MEM_stage_inst_dmem_ram_2620), .A2(MEM_stage_inst_dmem_n8169), .ZN(MEM_stage_inst_dmem_n6920) );
NAND2_X1 MEM_stage_inst_dmem_U7052 ( .A1(MEM_stage_inst_dmem_ram_2812), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n6921) );
NAND2_X1 MEM_stage_inst_dmem_U7051 ( .A1(MEM_stage_inst_dmem_n6919), .A2(MEM_stage_inst_dmem_n6918), .ZN(MEM_stage_inst_dmem_n6923) );
NAND2_X1 MEM_stage_inst_dmem_U7050 ( .A1(MEM_stage_inst_dmem_ram_2236), .A2(MEM_stage_inst_dmem_n7937), .ZN(MEM_stage_inst_dmem_n6918) );
NAND2_X1 MEM_stage_inst_dmem_U7049 ( .A1(MEM_stage_inst_dmem_ram_2796), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n6919) );
NOR2_X1 MEM_stage_inst_dmem_U7048 ( .A1(MEM_stage_inst_dmem_n6917), .A2(MEM_stage_inst_dmem_n6916), .ZN(MEM_stage_inst_dmem_n6925) );
NAND2_X1 MEM_stage_inst_dmem_U7047 ( .A1(MEM_stage_inst_dmem_n6915), .A2(MEM_stage_inst_dmem_n6914), .ZN(MEM_stage_inst_dmem_n6916) );
NAND2_X1 MEM_stage_inst_dmem_U7046 ( .A1(MEM_stage_inst_dmem_ram_2140), .A2(MEM_stage_inst_dmem_n7938), .ZN(MEM_stage_inst_dmem_n6914) );
NAND2_X1 MEM_stage_inst_dmem_U7045 ( .A1(MEM_stage_inst_dmem_ram_3068), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n6915) );
NAND2_X1 MEM_stage_inst_dmem_U7044 ( .A1(MEM_stage_inst_dmem_n6913), .A2(MEM_stage_inst_dmem_n6912), .ZN(MEM_stage_inst_dmem_n6917) );
NAND2_X1 MEM_stage_inst_dmem_U7043 ( .A1(MEM_stage_inst_dmem_ram_3052), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n6912) );
NAND2_X1 MEM_stage_inst_dmem_U7042 ( .A1(MEM_stage_inst_dmem_ram_2636), .A2(MEM_stage_inst_dmem_n7973), .ZN(MEM_stage_inst_dmem_n6913) );
NAND2_X1 MEM_stage_inst_dmem_U7041 ( .A1(MEM_stage_inst_dmem_n6911), .A2(MEM_stage_inst_dmem_n6910), .ZN(MEM_stage_inst_dmem_n6975) );
NOR2_X1 MEM_stage_inst_dmem_U7040 ( .A1(MEM_stage_inst_dmem_n6909), .A2(MEM_stage_inst_dmem_n6908), .ZN(MEM_stage_inst_dmem_n6910) );
NAND2_X1 MEM_stage_inst_dmem_U7039 ( .A1(MEM_stage_inst_dmem_n6907), .A2(MEM_stage_inst_dmem_n6906), .ZN(MEM_stage_inst_dmem_n6908) );
NOR2_X1 MEM_stage_inst_dmem_U7038 ( .A1(MEM_stage_inst_dmem_n6905), .A2(MEM_stage_inst_dmem_n6904), .ZN(MEM_stage_inst_dmem_n6906) );
NAND2_X1 MEM_stage_inst_dmem_U7037 ( .A1(MEM_stage_inst_dmem_n6903), .A2(MEM_stage_inst_dmem_n6902), .ZN(MEM_stage_inst_dmem_n6904) );
NAND2_X1 MEM_stage_inst_dmem_U7036 ( .A1(MEM_stage_inst_dmem_ram_2828), .A2(MEM_stage_inst_dmem_n7992), .ZN(MEM_stage_inst_dmem_n6902) );
NAND2_X1 MEM_stage_inst_dmem_U7035 ( .A1(MEM_stage_inst_dmem_ram_2076), .A2(MEM_stage_inst_dmem_n7887), .ZN(MEM_stage_inst_dmem_n6903) );
NAND2_X1 MEM_stage_inst_dmem_U7034 ( .A1(MEM_stage_inst_dmem_n6901), .A2(MEM_stage_inst_dmem_n6900), .ZN(MEM_stage_inst_dmem_n6905) );
NAND2_X1 MEM_stage_inst_dmem_U7033 ( .A1(MEM_stage_inst_dmem_ram_2764), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n6900) );
NAND2_X1 MEM_stage_inst_dmem_U7032 ( .A1(MEM_stage_inst_dmem_ram_2604), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n6901) );
NOR2_X1 MEM_stage_inst_dmem_U7031 ( .A1(MEM_stage_inst_dmem_n6899), .A2(MEM_stage_inst_dmem_n6898), .ZN(MEM_stage_inst_dmem_n6907) );
NAND2_X1 MEM_stage_inst_dmem_U7030 ( .A1(MEM_stage_inst_dmem_n6897), .A2(MEM_stage_inst_dmem_n6896), .ZN(MEM_stage_inst_dmem_n6898) );
NAND2_X1 MEM_stage_inst_dmem_U7029 ( .A1(MEM_stage_inst_dmem_ram_2524), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n6896) );
NAND2_X1 MEM_stage_inst_dmem_U7028 ( .A1(MEM_stage_inst_dmem_ram_2204), .A2(MEM_stage_inst_dmem_n7903), .ZN(MEM_stage_inst_dmem_n6897) );
NAND2_X1 MEM_stage_inst_dmem_U7027 ( .A1(MEM_stage_inst_dmem_n6895), .A2(MEM_stage_inst_dmem_n6894), .ZN(MEM_stage_inst_dmem_n6899) );
NAND2_X1 MEM_stage_inst_dmem_U7026 ( .A1(MEM_stage_inst_dmem_ram_2380), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n6894) );
NAND2_X1 MEM_stage_inst_dmem_U7025 ( .A1(MEM_stage_inst_dmem_ram_2668), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n6895) );
NAND2_X1 MEM_stage_inst_dmem_U7024 ( .A1(MEM_stage_inst_dmem_n6893), .A2(MEM_stage_inst_dmem_n6892), .ZN(MEM_stage_inst_dmem_n6909) );
NOR2_X1 MEM_stage_inst_dmem_U7023 ( .A1(MEM_stage_inst_dmem_n6891), .A2(MEM_stage_inst_dmem_n6890), .ZN(MEM_stage_inst_dmem_n6892) );
NAND2_X1 MEM_stage_inst_dmem_U7022 ( .A1(MEM_stage_inst_dmem_n6889), .A2(MEM_stage_inst_dmem_n6888), .ZN(MEM_stage_inst_dmem_n6890) );
NAND2_X1 MEM_stage_inst_dmem_U7021 ( .A1(MEM_stage_inst_dmem_ram_2508), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n6888) );
NAND2_X1 MEM_stage_inst_dmem_U7020 ( .A1(MEM_stage_inst_dmem_ram_2844), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n6889) );
NAND2_X1 MEM_stage_inst_dmem_U7019 ( .A1(MEM_stage_inst_dmem_n6887), .A2(MEM_stage_inst_dmem_n6886), .ZN(MEM_stage_inst_dmem_n6891) );
NAND2_X1 MEM_stage_inst_dmem_U7018 ( .A1(MEM_stage_inst_dmem_ram_2572), .A2(MEM_stage_inst_dmem_n8225), .ZN(MEM_stage_inst_dmem_n6886) );
NAND2_X1 MEM_stage_inst_dmem_U7017 ( .A1(MEM_stage_inst_dmem_ram_2316), .A2(MEM_stage_inst_dmem_n7898), .ZN(MEM_stage_inst_dmem_n6887) );
NOR2_X1 MEM_stage_inst_dmem_U7016 ( .A1(MEM_stage_inst_dmem_n6885), .A2(MEM_stage_inst_dmem_n6884), .ZN(MEM_stage_inst_dmem_n6893) );
NAND2_X1 MEM_stage_inst_dmem_U7015 ( .A1(MEM_stage_inst_dmem_n6883), .A2(MEM_stage_inst_dmem_n6882), .ZN(MEM_stage_inst_dmem_n6884) );
NAND2_X1 MEM_stage_inst_dmem_U7014 ( .A1(MEM_stage_inst_dmem_ram_2652), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n6882) );
NAND2_X1 MEM_stage_inst_dmem_U7013 ( .A1(MEM_stage_inst_dmem_ram_2780), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n6883) );
NAND2_X1 MEM_stage_inst_dmem_U7012 ( .A1(MEM_stage_inst_dmem_n6881), .A2(MEM_stage_inst_dmem_n6880), .ZN(MEM_stage_inst_dmem_n6885) );
NAND2_X1 MEM_stage_inst_dmem_U7011 ( .A1(MEM_stage_inst_dmem_ram_2588), .A2(MEM_stage_inst_dmem_n7884), .ZN(MEM_stage_inst_dmem_n6880) );
NAND2_X1 MEM_stage_inst_dmem_U7010 ( .A1(MEM_stage_inst_dmem_ram_2060), .A2(MEM_stage_inst_dmem_n7953), .ZN(MEM_stage_inst_dmem_n6881) );
NOR2_X1 MEM_stage_inst_dmem_U7009 ( .A1(MEM_stage_inst_dmem_n6879), .A2(MEM_stage_inst_dmem_n6878), .ZN(MEM_stage_inst_dmem_n6911) );
NAND2_X1 MEM_stage_inst_dmem_U7008 ( .A1(MEM_stage_inst_dmem_n6877), .A2(MEM_stage_inst_dmem_n6876), .ZN(MEM_stage_inst_dmem_n6878) );
NOR2_X1 MEM_stage_inst_dmem_U7007 ( .A1(MEM_stage_inst_dmem_n6875), .A2(MEM_stage_inst_dmem_n6874), .ZN(MEM_stage_inst_dmem_n6876) );
NAND2_X1 MEM_stage_inst_dmem_U7006 ( .A1(MEM_stage_inst_dmem_n6873), .A2(MEM_stage_inst_dmem_n6872), .ZN(MEM_stage_inst_dmem_n6874) );
NAND2_X1 MEM_stage_inst_dmem_U7005 ( .A1(MEM_stage_inst_dmem_ram_2988), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n6872) );
NAND2_X1 MEM_stage_inst_dmem_U7004 ( .A1(MEM_stage_inst_dmem_ram_2716), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n6873) );
NAND2_X1 MEM_stage_inst_dmem_U7003 ( .A1(MEM_stage_inst_dmem_n6871), .A2(MEM_stage_inst_dmem_n6870), .ZN(MEM_stage_inst_dmem_n6875) );
NAND2_X1 MEM_stage_inst_dmem_U7002 ( .A1(MEM_stage_inst_dmem_ram_2700), .A2(MEM_stage_inst_dmem_n7960), .ZN(MEM_stage_inst_dmem_n6870) );
NAND2_X1 MEM_stage_inst_dmem_U7001 ( .A1(MEM_stage_inst_dmem_ram_2268), .A2(MEM_stage_inst_dmem_n8206), .ZN(MEM_stage_inst_dmem_n6871) );
NOR2_X1 MEM_stage_inst_dmem_U7000 ( .A1(MEM_stage_inst_dmem_n6869), .A2(MEM_stage_inst_dmem_n6868), .ZN(MEM_stage_inst_dmem_n6877) );
NAND2_X1 MEM_stage_inst_dmem_U6999 ( .A1(MEM_stage_inst_dmem_n6867), .A2(MEM_stage_inst_dmem_n6866), .ZN(MEM_stage_inst_dmem_n6868) );
NAND2_X1 MEM_stage_inst_dmem_U6998 ( .A1(MEM_stage_inst_dmem_ram_2252), .A2(MEM_stage_inst_dmem_n8256), .ZN(MEM_stage_inst_dmem_n6866) );
NAND2_X1 MEM_stage_inst_dmem_U6997 ( .A1(MEM_stage_inst_dmem_ram_2556), .A2(MEM_stage_inst_dmem_n64), .ZN(MEM_stage_inst_dmem_n6867) );
NAND2_X1 MEM_stage_inst_dmem_U6996 ( .A1(MEM_stage_inst_dmem_n6865), .A2(MEM_stage_inst_dmem_n6864), .ZN(MEM_stage_inst_dmem_n6869) );
NAND2_X1 MEM_stage_inst_dmem_U6995 ( .A1(MEM_stage_inst_dmem_ram_2908), .A2(MEM_stage_inst_dmem_n3141), .ZN(MEM_stage_inst_dmem_n6864) );
NAND2_X1 MEM_stage_inst_dmem_U6994 ( .A1(MEM_stage_inst_dmem_ram_2284), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n6865) );
NAND2_X1 MEM_stage_inst_dmem_U6993 ( .A1(MEM_stage_inst_dmem_n6863), .A2(MEM_stage_inst_dmem_n6862), .ZN(MEM_stage_inst_dmem_n6879) );
NOR2_X1 MEM_stage_inst_dmem_U6992 ( .A1(MEM_stage_inst_dmem_n6861), .A2(MEM_stage_inst_dmem_n6860), .ZN(MEM_stage_inst_dmem_n6862) );
NAND2_X1 MEM_stage_inst_dmem_U6991 ( .A1(MEM_stage_inst_dmem_n6859), .A2(MEM_stage_inst_dmem_n6858), .ZN(MEM_stage_inst_dmem_n6860) );
NAND2_X1 MEM_stage_inst_dmem_U6990 ( .A1(MEM_stage_inst_dmem_ram_2892), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n6858) );
NAND2_X1 MEM_stage_inst_dmem_U6989 ( .A1(MEM_stage_inst_dmem_ram_2860), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n6859) );
NAND2_X1 MEM_stage_inst_dmem_U6988 ( .A1(MEM_stage_inst_dmem_n6857), .A2(MEM_stage_inst_dmem_n6856), .ZN(MEM_stage_inst_dmem_n6861) );
NAND2_X1 MEM_stage_inst_dmem_U6987 ( .A1(MEM_stage_inst_dmem_ram_2940), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n6856) );
NAND2_X1 MEM_stage_inst_dmem_U6986 ( .A1(MEM_stage_inst_dmem_ram_2108), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n6857) );
NOR2_X1 MEM_stage_inst_dmem_U6985 ( .A1(MEM_stage_inst_dmem_n6855), .A2(MEM_stage_inst_dmem_n6854), .ZN(MEM_stage_inst_dmem_n6863) );
NAND2_X1 MEM_stage_inst_dmem_U6984 ( .A1(MEM_stage_inst_dmem_n6853), .A2(MEM_stage_inst_dmem_n6852), .ZN(MEM_stage_inst_dmem_n6854) );
NAND2_X1 MEM_stage_inst_dmem_U6983 ( .A1(MEM_stage_inst_dmem_ram_2492), .A2(MEM_stage_inst_dmem_n7888), .ZN(MEM_stage_inst_dmem_n6852) );
NAND2_X1 MEM_stage_inst_dmem_U6982 ( .A1(MEM_stage_inst_dmem_ram_2092), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n6853) );
NAND2_X1 MEM_stage_inst_dmem_U6981 ( .A1(MEM_stage_inst_dmem_n6851), .A2(MEM_stage_inst_dmem_n6850), .ZN(MEM_stage_inst_dmem_n6855) );
NAND2_X1 MEM_stage_inst_dmem_U6980 ( .A1(MEM_stage_inst_dmem_ram_2956), .A2(MEM_stage_inst_dmem_n8193), .ZN(MEM_stage_inst_dmem_n6850) );
NAND2_X1 MEM_stage_inst_dmem_U6979 ( .A1(MEM_stage_inst_dmem_ram_2428), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n6851) );
NOR2_X1 MEM_stage_inst_dmem_U6978 ( .A1(MEM_stage_inst_dmem_n6849), .A2(MEM_stage_inst_dmem_n8152), .ZN(MEM_stage_inst_dmem_n6978) );
NOR2_X1 MEM_stage_inst_dmem_U6977 ( .A1(MEM_stage_inst_dmem_n6848), .A2(MEM_stage_inst_dmem_n6847), .ZN(MEM_stage_inst_dmem_n6849) );
NAND2_X1 MEM_stage_inst_dmem_U6976 ( .A1(MEM_stage_inst_dmem_n6846), .A2(MEM_stage_inst_dmem_n6845), .ZN(MEM_stage_inst_dmem_n6847) );
NOR2_X1 MEM_stage_inst_dmem_U6975 ( .A1(MEM_stage_inst_dmem_n6844), .A2(MEM_stage_inst_dmem_n6843), .ZN(MEM_stage_inst_dmem_n6845) );
NAND2_X1 MEM_stage_inst_dmem_U6974 ( .A1(MEM_stage_inst_dmem_n6842), .A2(MEM_stage_inst_dmem_n6841), .ZN(MEM_stage_inst_dmem_n6843) );
NOR2_X1 MEM_stage_inst_dmem_U6973 ( .A1(MEM_stage_inst_dmem_n6840), .A2(MEM_stage_inst_dmem_n6839), .ZN(MEM_stage_inst_dmem_n6841) );
NAND2_X1 MEM_stage_inst_dmem_U6972 ( .A1(MEM_stage_inst_dmem_n6838), .A2(MEM_stage_inst_dmem_n6837), .ZN(MEM_stage_inst_dmem_n6839) );
NAND2_X1 MEM_stage_inst_dmem_U6971 ( .A1(MEM_stage_inst_dmem_ram_1804), .A2(MEM_stage_inst_dmem_n8472), .ZN(MEM_stage_inst_dmem_n6837) );
NAND2_X1 MEM_stage_inst_dmem_U6970 ( .A1(MEM_stage_inst_dmem_ram_1756), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n6838) );
NAND2_X1 MEM_stage_inst_dmem_U6969 ( .A1(MEM_stage_inst_dmem_n6836), .A2(MEM_stage_inst_dmem_n6835), .ZN(MEM_stage_inst_dmem_n6840) );
NAND2_X1 MEM_stage_inst_dmem_U6968 ( .A1(MEM_stage_inst_dmem_ram_1708), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n6835) );
NAND2_X1 MEM_stage_inst_dmem_U6967 ( .A1(MEM_stage_inst_dmem_ram_1196), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n6836) );
NOR2_X1 MEM_stage_inst_dmem_U6966 ( .A1(MEM_stage_inst_dmem_n6834), .A2(MEM_stage_inst_dmem_n6833), .ZN(MEM_stage_inst_dmem_n6842) );
NAND2_X1 MEM_stage_inst_dmem_U6965 ( .A1(MEM_stage_inst_dmem_n6832), .A2(MEM_stage_inst_dmem_n6831), .ZN(MEM_stage_inst_dmem_n6833) );
NAND2_X1 MEM_stage_inst_dmem_U6964 ( .A1(MEM_stage_inst_dmem_ram_1788), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n6831) );
NAND2_X1 MEM_stage_inst_dmem_U6963 ( .A1(MEM_stage_inst_dmem_ram_1180), .A2(MEM_stage_inst_dmem_n44), .ZN(MEM_stage_inst_dmem_n6832) );
NAND2_X1 MEM_stage_inst_dmem_U6962 ( .A1(MEM_stage_inst_dmem_n6830), .A2(MEM_stage_inst_dmem_n6829), .ZN(MEM_stage_inst_dmem_n6834) );
NAND2_X1 MEM_stage_inst_dmem_U6961 ( .A1(MEM_stage_inst_dmem_ram_1916), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n6829) );
NAND2_X1 MEM_stage_inst_dmem_U6960 ( .A1(MEM_stage_inst_dmem_ram_1868), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n6830) );
NAND2_X1 MEM_stage_inst_dmem_U6959 ( .A1(MEM_stage_inst_dmem_n6828), .A2(MEM_stage_inst_dmem_n6827), .ZN(MEM_stage_inst_dmem_n6844) );
NOR2_X1 MEM_stage_inst_dmem_U6958 ( .A1(MEM_stage_inst_dmem_n6826), .A2(MEM_stage_inst_dmem_n6825), .ZN(MEM_stage_inst_dmem_n6827) );
NAND2_X1 MEM_stage_inst_dmem_U6957 ( .A1(MEM_stage_inst_dmem_n6824), .A2(MEM_stage_inst_dmem_n6823), .ZN(MEM_stage_inst_dmem_n6825) );
NAND2_X1 MEM_stage_inst_dmem_U6956 ( .A1(MEM_stage_inst_dmem_ram_1660), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n6823) );
NAND2_X1 MEM_stage_inst_dmem_U6955 ( .A1(MEM_stage_inst_dmem_ram_1628), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n6824) );
NAND2_X1 MEM_stage_inst_dmem_U6954 ( .A1(MEM_stage_inst_dmem_n6822), .A2(MEM_stage_inst_dmem_n6821), .ZN(MEM_stage_inst_dmem_n6826) );
NAND2_X1 MEM_stage_inst_dmem_U6953 ( .A1(MEM_stage_inst_dmem_ram_1116), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n6821) );
NAND2_X1 MEM_stage_inst_dmem_U6952 ( .A1(MEM_stage_inst_dmem_ram_2044), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n6822) );
NOR2_X1 MEM_stage_inst_dmem_U6951 ( .A1(MEM_stage_inst_dmem_n6820), .A2(MEM_stage_inst_dmem_n6819), .ZN(MEM_stage_inst_dmem_n6828) );
NAND2_X1 MEM_stage_inst_dmem_U6950 ( .A1(MEM_stage_inst_dmem_n6818), .A2(MEM_stage_inst_dmem_n6817), .ZN(MEM_stage_inst_dmem_n6819) );
NAND2_X1 MEM_stage_inst_dmem_U6949 ( .A1(MEM_stage_inst_dmem_ram_1980), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n6817) );
NAND2_X1 MEM_stage_inst_dmem_U6948 ( .A1(MEM_stage_inst_dmem_ram_1852), .A2(MEM_stage_inst_dmem_n8005), .ZN(MEM_stage_inst_dmem_n6818) );
NAND2_X1 MEM_stage_inst_dmem_U6947 ( .A1(MEM_stage_inst_dmem_n6816), .A2(MEM_stage_inst_dmem_n6815), .ZN(MEM_stage_inst_dmem_n6820) );
NAND2_X1 MEM_stage_inst_dmem_U6946 ( .A1(MEM_stage_inst_dmem_ram_1388), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n6815) );
NAND2_X1 MEM_stage_inst_dmem_U6945 ( .A1(MEM_stage_inst_dmem_ram_1148), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n6816) );
NOR2_X1 MEM_stage_inst_dmem_U6944 ( .A1(MEM_stage_inst_dmem_n6814), .A2(MEM_stage_inst_dmem_n6813), .ZN(MEM_stage_inst_dmem_n6846) );
NAND2_X1 MEM_stage_inst_dmem_U6943 ( .A1(MEM_stage_inst_dmem_n6812), .A2(MEM_stage_inst_dmem_n6811), .ZN(MEM_stage_inst_dmem_n6813) );
NOR2_X1 MEM_stage_inst_dmem_U6942 ( .A1(MEM_stage_inst_dmem_n6810), .A2(MEM_stage_inst_dmem_n6809), .ZN(MEM_stage_inst_dmem_n6811) );
NAND2_X1 MEM_stage_inst_dmem_U6941 ( .A1(MEM_stage_inst_dmem_n6808), .A2(MEM_stage_inst_dmem_n6807), .ZN(MEM_stage_inst_dmem_n6809) );
NAND2_X1 MEM_stage_inst_dmem_U6940 ( .A1(MEM_stage_inst_dmem_ram_1516), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n6807) );
NAND2_X1 MEM_stage_inst_dmem_U6939 ( .A1(MEM_stage_inst_dmem_ram_1548), .A2(MEM_stage_inst_dmem_n8225), .ZN(MEM_stage_inst_dmem_n6808) );
NAND2_X1 MEM_stage_inst_dmem_U6938 ( .A1(MEM_stage_inst_dmem_n6806), .A2(MEM_stage_inst_dmem_n6805), .ZN(MEM_stage_inst_dmem_n6810) );
NAND2_X1 MEM_stage_inst_dmem_U6937 ( .A1(MEM_stage_inst_dmem_ram_1324), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n6805) );
NAND2_X1 MEM_stage_inst_dmem_U6936 ( .A1(MEM_stage_inst_dmem_ram_1404), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n6806) );
NOR2_X1 MEM_stage_inst_dmem_U6935 ( .A1(MEM_stage_inst_dmem_n6804), .A2(MEM_stage_inst_dmem_n6803), .ZN(MEM_stage_inst_dmem_n6812) );
NAND2_X1 MEM_stage_inst_dmem_U6934 ( .A1(MEM_stage_inst_dmem_n6802), .A2(MEM_stage_inst_dmem_n6801), .ZN(MEM_stage_inst_dmem_n6803) );
NAND2_X1 MEM_stage_inst_dmem_U6933 ( .A1(MEM_stage_inst_dmem_ram_1884), .A2(MEM_stage_inst_dmem_n3141), .ZN(MEM_stage_inst_dmem_n6801) );
NAND2_X1 MEM_stage_inst_dmem_U6932 ( .A1(MEM_stage_inst_dmem_ram_1292), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n6802) );
NAND2_X1 MEM_stage_inst_dmem_U6931 ( .A1(MEM_stage_inst_dmem_n6800), .A2(MEM_stage_inst_dmem_n6799), .ZN(MEM_stage_inst_dmem_n6804) );
NAND2_X1 MEM_stage_inst_dmem_U6930 ( .A1(MEM_stage_inst_dmem_ram_1532), .A2(MEM_stage_inst_dmem_n64), .ZN(MEM_stage_inst_dmem_n6799) );
NAND2_X1 MEM_stage_inst_dmem_U6929 ( .A1(MEM_stage_inst_dmem_ram_1484), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n6800) );
NAND2_X1 MEM_stage_inst_dmem_U6928 ( .A1(MEM_stage_inst_dmem_n6798), .A2(MEM_stage_inst_dmem_n6797), .ZN(MEM_stage_inst_dmem_n6814) );
NOR2_X1 MEM_stage_inst_dmem_U6927 ( .A1(MEM_stage_inst_dmem_n6796), .A2(MEM_stage_inst_dmem_n6795), .ZN(MEM_stage_inst_dmem_n6797) );
NAND2_X1 MEM_stage_inst_dmem_U6926 ( .A1(MEM_stage_inst_dmem_n6794), .A2(MEM_stage_inst_dmem_n6793), .ZN(MEM_stage_inst_dmem_n6795) );
NAND2_X1 MEM_stage_inst_dmem_U6925 ( .A1(MEM_stage_inst_dmem_ram_1340), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n6793) );
NAND2_X1 MEM_stage_inst_dmem_U6924 ( .A1(MEM_stage_inst_dmem_ram_1580), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n6794) );
NAND2_X1 MEM_stage_inst_dmem_U6923 ( .A1(MEM_stage_inst_dmem_n6792), .A2(MEM_stage_inst_dmem_n6791), .ZN(MEM_stage_inst_dmem_n6796) );
NAND2_X1 MEM_stage_inst_dmem_U6922 ( .A1(MEM_stage_inst_dmem_ram_2012), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n6791) );
NAND2_X1 MEM_stage_inst_dmem_U6921 ( .A1(MEM_stage_inst_dmem_ram_1836), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n6792) );
NOR2_X1 MEM_stage_inst_dmem_U6920 ( .A1(MEM_stage_inst_dmem_n6790), .A2(MEM_stage_inst_dmem_n6789), .ZN(MEM_stage_inst_dmem_n6798) );
NAND2_X1 MEM_stage_inst_dmem_U6919 ( .A1(MEM_stage_inst_dmem_n6788), .A2(MEM_stage_inst_dmem_n6787), .ZN(MEM_stage_inst_dmem_n6789) );
NAND2_X1 MEM_stage_inst_dmem_U6918 ( .A1(MEM_stage_inst_dmem_ram_1468), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n6787) );
NAND2_X1 MEM_stage_inst_dmem_U6917 ( .A1(MEM_stage_inst_dmem_ram_1964), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n6788) );
NAND2_X1 MEM_stage_inst_dmem_U6916 ( .A1(MEM_stage_inst_dmem_n6786), .A2(MEM_stage_inst_dmem_n6785), .ZN(MEM_stage_inst_dmem_n6790) );
NAND2_X1 MEM_stage_inst_dmem_U6915 ( .A1(MEM_stage_inst_dmem_ram_1724), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n6785) );
NAND2_X1 MEM_stage_inst_dmem_U6914 ( .A1(MEM_stage_inst_dmem_ram_1612), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n6786) );
NAND2_X1 MEM_stage_inst_dmem_U6913 ( .A1(MEM_stage_inst_dmem_n6784), .A2(MEM_stage_inst_dmem_n6783), .ZN(MEM_stage_inst_dmem_n6848) );
NOR2_X1 MEM_stage_inst_dmem_U6912 ( .A1(MEM_stage_inst_dmem_n6782), .A2(MEM_stage_inst_dmem_n6781), .ZN(MEM_stage_inst_dmem_n6783) );
NAND2_X1 MEM_stage_inst_dmem_U6911 ( .A1(MEM_stage_inst_dmem_n6780), .A2(MEM_stage_inst_dmem_n6779), .ZN(MEM_stage_inst_dmem_n6781) );
NOR2_X1 MEM_stage_inst_dmem_U6910 ( .A1(MEM_stage_inst_dmem_n6778), .A2(MEM_stage_inst_dmem_n6777), .ZN(MEM_stage_inst_dmem_n6779) );
NAND2_X1 MEM_stage_inst_dmem_U6909 ( .A1(MEM_stage_inst_dmem_n6776), .A2(MEM_stage_inst_dmem_n6775), .ZN(MEM_stage_inst_dmem_n6777) );
NAND2_X1 MEM_stage_inst_dmem_U6908 ( .A1(MEM_stage_inst_dmem_ram_1900), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n6775) );
NAND2_X1 MEM_stage_inst_dmem_U6907 ( .A1(MEM_stage_inst_dmem_ram_1164), .A2(MEM_stage_inst_dmem_n8174), .ZN(MEM_stage_inst_dmem_n6776) );
NAND2_X1 MEM_stage_inst_dmem_U6906 ( .A1(MEM_stage_inst_dmem_n6774), .A2(MEM_stage_inst_dmem_n6773), .ZN(MEM_stage_inst_dmem_n6778) );
NAND2_X1 MEM_stage_inst_dmem_U6905 ( .A1(MEM_stage_inst_dmem_ram_1996), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n6773) );
NAND2_X1 MEM_stage_inst_dmem_U6904 ( .A1(MEM_stage_inst_dmem_ram_1932), .A2(MEM_stage_inst_dmem_n8193), .ZN(MEM_stage_inst_dmem_n6774) );
NOR2_X1 MEM_stage_inst_dmem_U6903 ( .A1(MEM_stage_inst_dmem_n6772), .A2(MEM_stage_inst_dmem_n6771), .ZN(MEM_stage_inst_dmem_n6780) );
NAND2_X1 MEM_stage_inst_dmem_U6902 ( .A1(MEM_stage_inst_dmem_n6770), .A2(MEM_stage_inst_dmem_n6769), .ZN(MEM_stage_inst_dmem_n6771) );
NAND2_X1 MEM_stage_inst_dmem_U6901 ( .A1(MEM_stage_inst_dmem_ram_1068), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n6769) );
NAND2_X1 MEM_stage_inst_dmem_U6900 ( .A1(MEM_stage_inst_dmem_ram_1212), .A2(MEM_stage_inst_dmem_n8434), .ZN(MEM_stage_inst_dmem_n6770) );
NAND2_X1 MEM_stage_inst_dmem_U6899 ( .A1(MEM_stage_inst_dmem_n6768), .A2(MEM_stage_inst_dmem_n6767), .ZN(MEM_stage_inst_dmem_n6772) );
NAND2_X1 MEM_stage_inst_dmem_U6898 ( .A1(MEM_stage_inst_dmem_ram_1052), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n6767) );
NAND2_X1 MEM_stage_inst_dmem_U6897 ( .A1(MEM_stage_inst_dmem_ram_1644), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n6768) );
NAND2_X1 MEM_stage_inst_dmem_U6896 ( .A1(MEM_stage_inst_dmem_n6766), .A2(MEM_stage_inst_dmem_n6765), .ZN(MEM_stage_inst_dmem_n6782) );
NOR2_X1 MEM_stage_inst_dmem_U6895 ( .A1(MEM_stage_inst_dmem_n6764), .A2(MEM_stage_inst_dmem_n6763), .ZN(MEM_stage_inst_dmem_n6765) );
NAND2_X1 MEM_stage_inst_dmem_U6894 ( .A1(MEM_stage_inst_dmem_n6762), .A2(MEM_stage_inst_dmem_n6761), .ZN(MEM_stage_inst_dmem_n6763) );
NAND2_X1 MEM_stage_inst_dmem_U6893 ( .A1(MEM_stage_inst_dmem_ram_1260), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n6761) );
NAND2_X1 MEM_stage_inst_dmem_U6892 ( .A1(MEM_stage_inst_dmem_ram_1036), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n6762) );
NAND2_X1 MEM_stage_inst_dmem_U6891 ( .A1(MEM_stage_inst_dmem_n6760), .A2(MEM_stage_inst_dmem_n6759), .ZN(MEM_stage_inst_dmem_n6764) );
NAND2_X1 MEM_stage_inst_dmem_U6890 ( .A1(MEM_stage_inst_dmem_ram_1436), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n6759) );
NAND2_X1 MEM_stage_inst_dmem_U6889 ( .A1(MEM_stage_inst_dmem_ram_1372), .A2(MEM_stage_inst_dmem_n3216), .ZN(MEM_stage_inst_dmem_n6760) );
NOR2_X1 MEM_stage_inst_dmem_U6888 ( .A1(MEM_stage_inst_dmem_n6758), .A2(MEM_stage_inst_dmem_n6757), .ZN(MEM_stage_inst_dmem_n6766) );
NAND2_X1 MEM_stage_inst_dmem_U6887 ( .A1(MEM_stage_inst_dmem_n6756), .A2(MEM_stage_inst_dmem_n6755), .ZN(MEM_stage_inst_dmem_n6757) );
NAND2_X1 MEM_stage_inst_dmem_U6886 ( .A1(MEM_stage_inst_dmem_ram_1452), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n6755) );
NAND2_X1 MEM_stage_inst_dmem_U6885 ( .A1(MEM_stage_inst_dmem_ram_1692), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n6756) );
NAND2_X1 MEM_stage_inst_dmem_U6884 ( .A1(MEM_stage_inst_dmem_n6754), .A2(MEM_stage_inst_dmem_n6753), .ZN(MEM_stage_inst_dmem_n6758) );
NAND2_X1 MEM_stage_inst_dmem_U6883 ( .A1(MEM_stage_inst_dmem_ram_1084), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n6753) );
NAND2_X1 MEM_stage_inst_dmem_U6882 ( .A1(MEM_stage_inst_dmem_ram_1100), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n6754) );
NOR2_X1 MEM_stage_inst_dmem_U6881 ( .A1(MEM_stage_inst_dmem_n6752), .A2(MEM_stage_inst_dmem_n6751), .ZN(MEM_stage_inst_dmem_n6784) );
NAND2_X1 MEM_stage_inst_dmem_U6880 ( .A1(MEM_stage_inst_dmem_n6750), .A2(MEM_stage_inst_dmem_n6749), .ZN(MEM_stage_inst_dmem_n6751) );
NOR2_X1 MEM_stage_inst_dmem_U6879 ( .A1(MEM_stage_inst_dmem_n6748), .A2(MEM_stage_inst_dmem_n6747), .ZN(MEM_stage_inst_dmem_n6749) );
NAND2_X1 MEM_stage_inst_dmem_U6878 ( .A1(MEM_stage_inst_dmem_n6746), .A2(MEM_stage_inst_dmem_n6745), .ZN(MEM_stage_inst_dmem_n6747) );
NAND2_X1 MEM_stage_inst_dmem_U6877 ( .A1(MEM_stage_inst_dmem_ram_1820), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n6745) );
NAND2_X1 MEM_stage_inst_dmem_U6876 ( .A1(MEM_stage_inst_dmem_ram_1564), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n6746) );
NAND2_X1 MEM_stage_inst_dmem_U6875 ( .A1(MEM_stage_inst_dmem_n6744), .A2(MEM_stage_inst_dmem_n6743), .ZN(MEM_stage_inst_dmem_n6748) );
NAND2_X1 MEM_stage_inst_dmem_U6874 ( .A1(MEM_stage_inst_dmem_ram_1228), .A2(MEM_stage_inst_dmem_n8256), .ZN(MEM_stage_inst_dmem_n6743) );
NAND2_X1 MEM_stage_inst_dmem_U6873 ( .A1(MEM_stage_inst_dmem_ram_1308), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n6744) );
NOR2_X1 MEM_stage_inst_dmem_U6872 ( .A1(MEM_stage_inst_dmem_n6742), .A2(MEM_stage_inst_dmem_n6741), .ZN(MEM_stage_inst_dmem_n6750) );
NAND2_X1 MEM_stage_inst_dmem_U6871 ( .A1(MEM_stage_inst_dmem_n6740), .A2(MEM_stage_inst_dmem_n6739), .ZN(MEM_stage_inst_dmem_n6741) );
NAND2_X1 MEM_stage_inst_dmem_U6870 ( .A1(MEM_stage_inst_dmem_ram_1676), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n6739) );
NAND2_X1 MEM_stage_inst_dmem_U6869 ( .A1(MEM_stage_inst_dmem_ram_1500), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n6740) );
NAND2_X1 MEM_stage_inst_dmem_U6868 ( .A1(MEM_stage_inst_dmem_n6738), .A2(MEM_stage_inst_dmem_n6737), .ZN(MEM_stage_inst_dmem_n6742) );
NAND2_X1 MEM_stage_inst_dmem_U6867 ( .A1(MEM_stage_inst_dmem_ram_1356), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n6737) );
NAND2_X1 MEM_stage_inst_dmem_U6866 ( .A1(MEM_stage_inst_dmem_ram_1740), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n6738) );
NAND2_X1 MEM_stage_inst_dmem_U6865 ( .A1(MEM_stage_inst_dmem_n6736), .A2(MEM_stage_inst_dmem_n6735), .ZN(MEM_stage_inst_dmem_n6752) );
NOR2_X1 MEM_stage_inst_dmem_U6864 ( .A1(MEM_stage_inst_dmem_n6734), .A2(MEM_stage_inst_dmem_n6733), .ZN(MEM_stage_inst_dmem_n6735) );
NAND2_X1 MEM_stage_inst_dmem_U6863 ( .A1(MEM_stage_inst_dmem_n6732), .A2(MEM_stage_inst_dmem_n6731), .ZN(MEM_stage_inst_dmem_n6733) );
NAND2_X1 MEM_stage_inst_dmem_U6862 ( .A1(MEM_stage_inst_dmem_ram_1596), .A2(MEM_stage_inst_dmem_n8169), .ZN(MEM_stage_inst_dmem_n6731) );
NAND2_X1 MEM_stage_inst_dmem_U6861 ( .A1(MEM_stage_inst_dmem_ram_1772), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n6732) );
NAND2_X1 MEM_stage_inst_dmem_U6860 ( .A1(MEM_stage_inst_dmem_n6730), .A2(MEM_stage_inst_dmem_n6729), .ZN(MEM_stage_inst_dmem_n6734) );
NAND2_X1 MEM_stage_inst_dmem_U6859 ( .A1(MEM_stage_inst_dmem_ram_1948), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n6729) );
NAND2_X1 MEM_stage_inst_dmem_U6858 ( .A1(MEM_stage_inst_dmem_ram_1420), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n6730) );
NOR2_X1 MEM_stage_inst_dmem_U6857 ( .A1(MEM_stage_inst_dmem_n6728), .A2(MEM_stage_inst_dmem_n6727), .ZN(MEM_stage_inst_dmem_n6736) );
NAND2_X1 MEM_stage_inst_dmem_U6856 ( .A1(MEM_stage_inst_dmem_n6726), .A2(MEM_stage_inst_dmem_n6725), .ZN(MEM_stage_inst_dmem_n6727) );
NAND2_X1 MEM_stage_inst_dmem_U6855 ( .A1(MEM_stage_inst_dmem_ram_1276), .A2(MEM_stage_inst_dmem_n7914), .ZN(MEM_stage_inst_dmem_n6725) );
NAND2_X1 MEM_stage_inst_dmem_U6854 ( .A1(MEM_stage_inst_dmem_ram_1244), .A2(MEM_stage_inst_dmem_n8206), .ZN(MEM_stage_inst_dmem_n6726) );
NAND2_X1 MEM_stage_inst_dmem_U6853 ( .A1(MEM_stage_inst_dmem_n6724), .A2(MEM_stage_inst_dmem_n6723), .ZN(MEM_stage_inst_dmem_n6728) );
NAND2_X1 MEM_stage_inst_dmem_U6852 ( .A1(MEM_stage_inst_dmem_ram_2028), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n6723) );
NAND2_X1 MEM_stage_inst_dmem_U6851 ( .A1(MEM_stage_inst_dmem_ram_1132), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n6724) );
NOR2_X1 MEM_stage_inst_dmem_U6850 ( .A1(MEM_stage_inst_dmem_n6722), .A2(MEM_stage_inst_dmem_n6721), .ZN(MEM_stage_inst_dmem_n6980) );
NOR2_X1 MEM_stage_inst_dmem_U6849 ( .A1(MEM_stage_inst_dmem_n6720), .A2(MEM_stage_inst_dmem_n8417), .ZN(MEM_stage_inst_dmem_n6721) );
NOR2_X1 MEM_stage_inst_dmem_U6848 ( .A1(MEM_stage_inst_dmem_n6719), .A2(MEM_stage_inst_dmem_n6718), .ZN(MEM_stage_inst_dmem_n6720) );
NAND2_X1 MEM_stage_inst_dmem_U6847 ( .A1(MEM_stage_inst_dmem_n6717), .A2(MEM_stage_inst_dmem_n6716), .ZN(MEM_stage_inst_dmem_n6718) );
NOR2_X1 MEM_stage_inst_dmem_U6846 ( .A1(MEM_stage_inst_dmem_n6715), .A2(MEM_stage_inst_dmem_n6714), .ZN(MEM_stage_inst_dmem_n6716) );
NAND2_X1 MEM_stage_inst_dmem_U6845 ( .A1(MEM_stage_inst_dmem_n6713), .A2(MEM_stage_inst_dmem_n6712), .ZN(MEM_stage_inst_dmem_n6714) );
NOR2_X1 MEM_stage_inst_dmem_U6844 ( .A1(MEM_stage_inst_dmem_n6711), .A2(MEM_stage_inst_dmem_n6710), .ZN(MEM_stage_inst_dmem_n6712) );
NAND2_X1 MEM_stage_inst_dmem_U6843 ( .A1(MEM_stage_inst_dmem_n6709), .A2(MEM_stage_inst_dmem_n6708), .ZN(MEM_stage_inst_dmem_n6710) );
NAND2_X1 MEM_stage_inst_dmem_U6842 ( .A1(MEM_stage_inst_dmem_ram_3372), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n6708) );
NAND2_X1 MEM_stage_inst_dmem_U6841 ( .A1(MEM_stage_inst_dmem_ram_3676), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n6709) );
NAND2_X1 MEM_stage_inst_dmem_U6840 ( .A1(MEM_stage_inst_dmem_n6707), .A2(MEM_stage_inst_dmem_n6706), .ZN(MEM_stage_inst_dmem_n6711) );
NAND2_X1 MEM_stage_inst_dmem_U6839 ( .A1(MEM_stage_inst_dmem_ram_3628), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n6706) );
NAND2_X1 MEM_stage_inst_dmem_U6838 ( .A1(MEM_stage_inst_dmem_ram_3612), .A2(MEM_stage_inst_dmem_n7884), .ZN(MEM_stage_inst_dmem_n6707) );
NOR2_X1 MEM_stage_inst_dmem_U6837 ( .A1(MEM_stage_inst_dmem_n6705), .A2(MEM_stage_inst_dmem_n6704), .ZN(MEM_stage_inst_dmem_n6713) );
NAND2_X1 MEM_stage_inst_dmem_U6836 ( .A1(MEM_stage_inst_dmem_n6703), .A2(MEM_stage_inst_dmem_n6702), .ZN(MEM_stage_inst_dmem_n6704) );
NAND2_X1 MEM_stage_inst_dmem_U6835 ( .A1(MEM_stage_inst_dmem_ram_3212), .A2(MEM_stage_inst_dmem_n8174), .ZN(MEM_stage_inst_dmem_n6702) );
NAND2_X1 MEM_stage_inst_dmem_U6834 ( .A1(MEM_stage_inst_dmem_ram_3756), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n6703) );
NAND2_X1 MEM_stage_inst_dmem_U6833 ( .A1(MEM_stage_inst_dmem_n6701), .A2(MEM_stage_inst_dmem_n6700), .ZN(MEM_stage_inst_dmem_n6705) );
NAND2_X1 MEM_stage_inst_dmem_U6832 ( .A1(MEM_stage_inst_dmem_ram_3292), .A2(MEM_stage_inst_dmem_n8206), .ZN(MEM_stage_inst_dmem_n6700) );
NAND2_X1 MEM_stage_inst_dmem_U6831 ( .A1(MEM_stage_inst_dmem_ram_3228), .A2(MEM_stage_inst_dmem_n7903), .ZN(MEM_stage_inst_dmem_n6701) );
NAND2_X1 MEM_stage_inst_dmem_U6830 ( .A1(MEM_stage_inst_dmem_n6699), .A2(MEM_stage_inst_dmem_n6698), .ZN(MEM_stage_inst_dmem_n6715) );
NOR2_X1 MEM_stage_inst_dmem_U6829 ( .A1(MEM_stage_inst_dmem_n6697), .A2(MEM_stage_inst_dmem_n6696), .ZN(MEM_stage_inst_dmem_n6698) );
NAND2_X1 MEM_stage_inst_dmem_U6828 ( .A1(MEM_stage_inst_dmem_n6695), .A2(MEM_stage_inst_dmem_n6694), .ZN(MEM_stage_inst_dmem_n6696) );
NAND2_X1 MEM_stage_inst_dmem_U6827 ( .A1(MEM_stage_inst_dmem_ram_3852), .A2(MEM_stage_inst_dmem_n7992), .ZN(MEM_stage_inst_dmem_n6694) );
NAND2_X1 MEM_stage_inst_dmem_U6826 ( .A1(MEM_stage_inst_dmem_ram_3884), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n6695) );
NAND2_X1 MEM_stage_inst_dmem_U6825 ( .A1(MEM_stage_inst_dmem_n6693), .A2(MEM_stage_inst_dmem_n6692), .ZN(MEM_stage_inst_dmem_n6697) );
NAND2_X1 MEM_stage_inst_dmem_U6824 ( .A1(MEM_stage_inst_dmem_ram_4076), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n6692) );
NAND2_X1 MEM_stage_inst_dmem_U6823 ( .A1(MEM_stage_inst_dmem_ram_3468), .A2(MEM_stage_inst_dmem_n7930), .ZN(MEM_stage_inst_dmem_n6693) );
NOR2_X1 MEM_stage_inst_dmem_U6822 ( .A1(MEM_stage_inst_dmem_n6691), .A2(MEM_stage_inst_dmem_n6690), .ZN(MEM_stage_inst_dmem_n6699) );
NAND2_X1 MEM_stage_inst_dmem_U6821 ( .A1(MEM_stage_inst_dmem_n6689), .A2(MEM_stage_inst_dmem_n6688), .ZN(MEM_stage_inst_dmem_n6690) );
NAND2_X1 MEM_stage_inst_dmem_U6820 ( .A1(MEM_stage_inst_dmem_ram_3532), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n6688) );
NAND2_X1 MEM_stage_inst_dmem_U6819 ( .A1(MEM_stage_inst_dmem_ram_3244), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n6689) );
NAND2_X1 MEM_stage_inst_dmem_U6818 ( .A1(MEM_stage_inst_dmem_n6687), .A2(MEM_stage_inst_dmem_n6686), .ZN(MEM_stage_inst_dmem_n6691) );
NAND2_X1 MEM_stage_inst_dmem_U6817 ( .A1(MEM_stage_inst_dmem_ram_4092), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n6686) );
NAND2_X1 MEM_stage_inst_dmem_U6816 ( .A1(MEM_stage_inst_dmem_ram_3340), .A2(MEM_stage_inst_dmem_n7898), .ZN(MEM_stage_inst_dmem_n6687) );
NOR2_X1 MEM_stage_inst_dmem_U6815 ( .A1(MEM_stage_inst_dmem_n6685), .A2(MEM_stage_inst_dmem_n6684), .ZN(MEM_stage_inst_dmem_n6717) );
NAND2_X1 MEM_stage_inst_dmem_U6814 ( .A1(MEM_stage_inst_dmem_n6683), .A2(MEM_stage_inst_dmem_n6682), .ZN(MEM_stage_inst_dmem_n6684) );
NOR2_X1 MEM_stage_inst_dmem_U6813 ( .A1(MEM_stage_inst_dmem_n6681), .A2(MEM_stage_inst_dmem_n6680), .ZN(MEM_stage_inst_dmem_n6682) );
NAND2_X1 MEM_stage_inst_dmem_U6812 ( .A1(MEM_stage_inst_dmem_n6679), .A2(MEM_stage_inst_dmem_n6678), .ZN(MEM_stage_inst_dmem_n6680) );
NAND2_X1 MEM_stage_inst_dmem_U6811 ( .A1(MEM_stage_inst_dmem_ram_3772), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n6678) );
NAND2_X1 MEM_stage_inst_dmem_U6810 ( .A1(MEM_stage_inst_dmem_ram_3548), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n6679) );
NAND2_X1 MEM_stage_inst_dmem_U6809 ( .A1(MEM_stage_inst_dmem_n6677), .A2(MEM_stage_inst_dmem_n6676), .ZN(MEM_stage_inst_dmem_n6681) );
NAND2_X1 MEM_stage_inst_dmem_U6808 ( .A1(MEM_stage_inst_dmem_ram_3564), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n6676) );
NAND2_X1 MEM_stage_inst_dmem_U6807 ( .A1(MEM_stage_inst_dmem_ram_3900), .A2(MEM_stage_inst_dmem_n8005), .ZN(MEM_stage_inst_dmem_n6677) );
NOR2_X1 MEM_stage_inst_dmem_U6806 ( .A1(MEM_stage_inst_dmem_n6675), .A2(MEM_stage_inst_dmem_n6674), .ZN(MEM_stage_inst_dmem_n6683) );
NAND2_X1 MEM_stage_inst_dmem_U6805 ( .A1(MEM_stage_inst_dmem_n6673), .A2(MEM_stage_inst_dmem_n6672), .ZN(MEM_stage_inst_dmem_n6674) );
NAND2_X1 MEM_stage_inst_dmem_U6804 ( .A1(MEM_stage_inst_dmem_ram_3916), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n6672) );
NAND2_X1 MEM_stage_inst_dmem_U6803 ( .A1(MEM_stage_inst_dmem_ram_3740), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n6673) );
NAND2_X1 MEM_stage_inst_dmem_U6802 ( .A1(MEM_stage_inst_dmem_n6671), .A2(MEM_stage_inst_dmem_n6670), .ZN(MEM_stage_inst_dmem_n6675) );
NAND2_X1 MEM_stage_inst_dmem_U6801 ( .A1(MEM_stage_inst_dmem_ram_3932), .A2(MEM_stage_inst_dmem_n3141), .ZN(MEM_stage_inst_dmem_n6670) );
NAND2_X1 MEM_stage_inst_dmem_U6800 ( .A1(MEM_stage_inst_dmem_ram_3436), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n6671) );
NAND2_X1 MEM_stage_inst_dmem_U6799 ( .A1(MEM_stage_inst_dmem_n6669), .A2(MEM_stage_inst_dmem_n6668), .ZN(MEM_stage_inst_dmem_n6685) );
NOR2_X1 MEM_stage_inst_dmem_U6798 ( .A1(MEM_stage_inst_dmem_n6667), .A2(MEM_stage_inst_dmem_n6666), .ZN(MEM_stage_inst_dmem_n6668) );
NAND2_X1 MEM_stage_inst_dmem_U6797 ( .A1(MEM_stage_inst_dmem_n6665), .A2(MEM_stage_inst_dmem_n6664), .ZN(MEM_stage_inst_dmem_n6666) );
NAND2_X1 MEM_stage_inst_dmem_U6796 ( .A1(MEM_stage_inst_dmem_ram_3148), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n6664) );
NAND2_X1 MEM_stage_inst_dmem_U6795 ( .A1(MEM_stage_inst_dmem_ram_3500), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n6665) );
NAND2_X1 MEM_stage_inst_dmem_U6794 ( .A1(MEM_stage_inst_dmem_n6663), .A2(MEM_stage_inst_dmem_n6662), .ZN(MEM_stage_inst_dmem_n6667) );
NAND2_X1 MEM_stage_inst_dmem_U6793 ( .A1(MEM_stage_inst_dmem_ram_3276), .A2(MEM_stage_inst_dmem_n8256), .ZN(MEM_stage_inst_dmem_n6662) );
NAND2_X1 MEM_stage_inst_dmem_U6792 ( .A1(MEM_stage_inst_dmem_ram_3196), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n6663) );
NOR2_X1 MEM_stage_inst_dmem_U6791 ( .A1(MEM_stage_inst_dmem_n6661), .A2(MEM_stage_inst_dmem_n6660), .ZN(MEM_stage_inst_dmem_n6669) );
NAND2_X1 MEM_stage_inst_dmem_U6790 ( .A1(MEM_stage_inst_dmem_n6659), .A2(MEM_stage_inst_dmem_n6658), .ZN(MEM_stage_inst_dmem_n6660) );
NAND2_X1 MEM_stage_inst_dmem_U6789 ( .A1(MEM_stage_inst_dmem_ram_3788), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n6658) );
NAND2_X1 MEM_stage_inst_dmem_U6788 ( .A1(MEM_stage_inst_dmem_ram_3660), .A2(MEM_stage_inst_dmem_n7973), .ZN(MEM_stage_inst_dmem_n6659) );
NAND2_X1 MEM_stage_inst_dmem_U6787 ( .A1(MEM_stage_inst_dmem_n6657), .A2(MEM_stage_inst_dmem_n6656), .ZN(MEM_stage_inst_dmem_n6661) );
NAND2_X1 MEM_stage_inst_dmem_U6786 ( .A1(MEM_stage_inst_dmem_ram_3404), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n6656) );
NAND2_X1 MEM_stage_inst_dmem_U6785 ( .A1(MEM_stage_inst_dmem_ram_3996), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n6657) );
NAND2_X1 MEM_stage_inst_dmem_U6784 ( .A1(MEM_stage_inst_dmem_n6655), .A2(MEM_stage_inst_dmem_n6654), .ZN(MEM_stage_inst_dmem_n6719) );
NOR2_X1 MEM_stage_inst_dmem_U6783 ( .A1(MEM_stage_inst_dmem_n6653), .A2(MEM_stage_inst_dmem_n6652), .ZN(MEM_stage_inst_dmem_n6654) );
NAND2_X1 MEM_stage_inst_dmem_U6782 ( .A1(MEM_stage_inst_dmem_n6651), .A2(MEM_stage_inst_dmem_n6650), .ZN(MEM_stage_inst_dmem_n6652) );
NOR2_X1 MEM_stage_inst_dmem_U6781 ( .A1(MEM_stage_inst_dmem_n6649), .A2(MEM_stage_inst_dmem_n6648), .ZN(MEM_stage_inst_dmem_n6650) );
NAND2_X1 MEM_stage_inst_dmem_U6780 ( .A1(MEM_stage_inst_dmem_n6647), .A2(MEM_stage_inst_dmem_n6646), .ZN(MEM_stage_inst_dmem_n6648) );
NAND2_X1 MEM_stage_inst_dmem_U6779 ( .A1(MEM_stage_inst_dmem_ram_3516), .A2(MEM_stage_inst_dmem_n7888), .ZN(MEM_stage_inst_dmem_n6646) );
NAND2_X1 MEM_stage_inst_dmem_U6778 ( .A1(MEM_stage_inst_dmem_ram_4028), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n6647) );
NAND2_X1 MEM_stage_inst_dmem_U6777 ( .A1(MEM_stage_inst_dmem_n6645), .A2(MEM_stage_inst_dmem_n6644), .ZN(MEM_stage_inst_dmem_n6649) );
NAND2_X1 MEM_stage_inst_dmem_U6776 ( .A1(MEM_stage_inst_dmem_ram_3132), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n6644) );
NAND2_X1 MEM_stage_inst_dmem_U6775 ( .A1(MEM_stage_inst_dmem_ram_3804), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n6645) );
NOR2_X1 MEM_stage_inst_dmem_U6774 ( .A1(MEM_stage_inst_dmem_n6643), .A2(MEM_stage_inst_dmem_n6642), .ZN(MEM_stage_inst_dmem_n6651) );
NAND2_X1 MEM_stage_inst_dmem_U6773 ( .A1(MEM_stage_inst_dmem_n6641), .A2(MEM_stage_inst_dmem_n6640), .ZN(MEM_stage_inst_dmem_n6642) );
NAND2_X1 MEM_stage_inst_dmem_U6772 ( .A1(MEM_stage_inst_dmem_ram_3100), .A2(MEM_stage_inst_dmem_n7887), .ZN(MEM_stage_inst_dmem_n6640) );
NAND2_X1 MEM_stage_inst_dmem_U6771 ( .A1(MEM_stage_inst_dmem_ram_3868), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n6641) );
NAND2_X1 MEM_stage_inst_dmem_U6770 ( .A1(MEM_stage_inst_dmem_n6639), .A2(MEM_stage_inst_dmem_n6638), .ZN(MEM_stage_inst_dmem_n6643) );
NAND2_X1 MEM_stage_inst_dmem_U6769 ( .A1(MEM_stage_inst_dmem_ram_3692), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n6638) );
NAND2_X1 MEM_stage_inst_dmem_U6768 ( .A1(MEM_stage_inst_dmem_ram_3084), .A2(MEM_stage_inst_dmem_n7953), .ZN(MEM_stage_inst_dmem_n6639) );
NAND2_X1 MEM_stage_inst_dmem_U6767 ( .A1(MEM_stage_inst_dmem_n6637), .A2(MEM_stage_inst_dmem_n6636), .ZN(MEM_stage_inst_dmem_n6653) );
NOR2_X1 MEM_stage_inst_dmem_U6766 ( .A1(MEM_stage_inst_dmem_n6635), .A2(MEM_stage_inst_dmem_n6634), .ZN(MEM_stage_inst_dmem_n6636) );
NAND2_X1 MEM_stage_inst_dmem_U6765 ( .A1(MEM_stage_inst_dmem_n6633), .A2(MEM_stage_inst_dmem_n6632), .ZN(MEM_stage_inst_dmem_n6634) );
NAND2_X1 MEM_stage_inst_dmem_U6764 ( .A1(MEM_stage_inst_dmem_ram_4060), .A2(MEM_stage_inst_dmem_n7895), .ZN(MEM_stage_inst_dmem_n6632) );
NAND2_X1 MEM_stage_inst_dmem_U6763 ( .A1(MEM_stage_inst_dmem_ram_3420), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n6633) );
NAND2_X1 MEM_stage_inst_dmem_U6762 ( .A1(MEM_stage_inst_dmem_n6631), .A2(MEM_stage_inst_dmem_n6630), .ZN(MEM_stage_inst_dmem_n6635) );
NAND2_X1 MEM_stage_inst_dmem_U6761 ( .A1(MEM_stage_inst_dmem_ram_3964), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n6630) );
NAND2_X1 MEM_stage_inst_dmem_U6760 ( .A1(MEM_stage_inst_dmem_ram_3836), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n6631) );
NOR2_X1 MEM_stage_inst_dmem_U6759 ( .A1(MEM_stage_inst_dmem_n6629), .A2(MEM_stage_inst_dmem_n6628), .ZN(MEM_stage_inst_dmem_n6637) );
NAND2_X1 MEM_stage_inst_dmem_U6758 ( .A1(MEM_stage_inst_dmem_n6627), .A2(MEM_stage_inst_dmem_n6626), .ZN(MEM_stage_inst_dmem_n6628) );
NAND2_X1 MEM_stage_inst_dmem_U6757 ( .A1(MEM_stage_inst_dmem_ram_3644), .A2(MEM_stage_inst_dmem_n8169), .ZN(MEM_stage_inst_dmem_n6626) );
NAND2_X1 MEM_stage_inst_dmem_U6756 ( .A1(MEM_stage_inst_dmem_ram_3708), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n6627) );
NAND2_X1 MEM_stage_inst_dmem_U6755 ( .A1(MEM_stage_inst_dmem_n6625), .A2(MEM_stage_inst_dmem_n6624), .ZN(MEM_stage_inst_dmem_n6629) );
NAND2_X1 MEM_stage_inst_dmem_U6754 ( .A1(MEM_stage_inst_dmem_ram_3948), .A2(MEM_stage_inst_dmem_n7923), .ZN(MEM_stage_inst_dmem_n6624) );
NAND2_X1 MEM_stage_inst_dmem_U6753 ( .A1(MEM_stage_inst_dmem_ram_3260), .A2(MEM_stage_inst_dmem_n7937), .ZN(MEM_stage_inst_dmem_n6625) );
NOR2_X1 MEM_stage_inst_dmem_U6752 ( .A1(MEM_stage_inst_dmem_n6623), .A2(MEM_stage_inst_dmem_n6622), .ZN(MEM_stage_inst_dmem_n6655) );
NAND2_X1 MEM_stage_inst_dmem_U6751 ( .A1(MEM_stage_inst_dmem_n6621), .A2(MEM_stage_inst_dmem_n6620), .ZN(MEM_stage_inst_dmem_n6622) );
NOR2_X1 MEM_stage_inst_dmem_U6750 ( .A1(MEM_stage_inst_dmem_n6619), .A2(MEM_stage_inst_dmem_n6618), .ZN(MEM_stage_inst_dmem_n6620) );
NAND2_X1 MEM_stage_inst_dmem_U6749 ( .A1(MEM_stage_inst_dmem_n6617), .A2(MEM_stage_inst_dmem_n6616), .ZN(MEM_stage_inst_dmem_n6618) );
NAND2_X1 MEM_stage_inst_dmem_U6748 ( .A1(MEM_stage_inst_dmem_ram_3388), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n6616) );
NAND2_X1 MEM_stage_inst_dmem_U6747 ( .A1(MEM_stage_inst_dmem_ram_3116), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n6617) );
NAND2_X1 MEM_stage_inst_dmem_U6746 ( .A1(MEM_stage_inst_dmem_n6615), .A2(MEM_stage_inst_dmem_n6614), .ZN(MEM_stage_inst_dmem_n6619) );
NAND2_X1 MEM_stage_inst_dmem_U6745 ( .A1(MEM_stage_inst_dmem_ram_3164), .A2(MEM_stage_inst_dmem_n7938), .ZN(MEM_stage_inst_dmem_n6614) );
NAND2_X1 MEM_stage_inst_dmem_U6744 ( .A1(MEM_stage_inst_dmem_ram_3820), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n6615) );
NOR2_X1 MEM_stage_inst_dmem_U6743 ( .A1(MEM_stage_inst_dmem_n6613), .A2(MEM_stage_inst_dmem_n6612), .ZN(MEM_stage_inst_dmem_n6621) );
NAND2_X1 MEM_stage_inst_dmem_U6742 ( .A1(MEM_stage_inst_dmem_n6611), .A2(MEM_stage_inst_dmem_n6610), .ZN(MEM_stage_inst_dmem_n6612) );
NAND2_X1 MEM_stage_inst_dmem_U6741 ( .A1(MEM_stage_inst_dmem_ram_3980), .A2(MEM_stage_inst_dmem_n8193), .ZN(MEM_stage_inst_dmem_n6610) );
NAND2_X1 MEM_stage_inst_dmem_U6740 ( .A1(MEM_stage_inst_dmem_ram_3324), .A2(MEM_stage_inst_dmem_n7914), .ZN(MEM_stage_inst_dmem_n6611) );
NAND2_X1 MEM_stage_inst_dmem_U6739 ( .A1(MEM_stage_inst_dmem_n6609), .A2(MEM_stage_inst_dmem_n6608), .ZN(MEM_stage_inst_dmem_n6613) );
NAND2_X1 MEM_stage_inst_dmem_U6738 ( .A1(MEM_stage_inst_dmem_ram_3724), .A2(MEM_stage_inst_dmem_n7960), .ZN(MEM_stage_inst_dmem_n6608) );
NAND2_X1 MEM_stage_inst_dmem_U6737 ( .A1(MEM_stage_inst_dmem_ram_4044), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n6609) );
NAND2_X1 MEM_stage_inst_dmem_U6736 ( .A1(MEM_stage_inst_dmem_n6607), .A2(MEM_stage_inst_dmem_n6606), .ZN(MEM_stage_inst_dmem_n6623) );
NOR2_X1 MEM_stage_inst_dmem_U6735 ( .A1(MEM_stage_inst_dmem_n6605), .A2(MEM_stage_inst_dmem_n6604), .ZN(MEM_stage_inst_dmem_n6606) );
NAND2_X1 MEM_stage_inst_dmem_U6734 ( .A1(MEM_stage_inst_dmem_n6603), .A2(MEM_stage_inst_dmem_n6602), .ZN(MEM_stage_inst_dmem_n6604) );
NAND2_X1 MEM_stage_inst_dmem_U6733 ( .A1(MEM_stage_inst_dmem_ram_4012), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n6602) );
NAND2_X1 MEM_stage_inst_dmem_U6732 ( .A1(MEM_stage_inst_dmem_ram_3180), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n6603) );
NAND2_X1 MEM_stage_inst_dmem_U6731 ( .A1(MEM_stage_inst_dmem_n6601), .A2(MEM_stage_inst_dmem_n6600), .ZN(MEM_stage_inst_dmem_n6605) );
NAND2_X1 MEM_stage_inst_dmem_U6730 ( .A1(MEM_stage_inst_dmem_ram_3484), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n6600) );
NAND2_X1 MEM_stage_inst_dmem_U6729 ( .A1(MEM_stage_inst_dmem_ram_3452), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n6601) );
NOR2_X1 MEM_stage_inst_dmem_U6728 ( .A1(MEM_stage_inst_dmem_n6599), .A2(MEM_stage_inst_dmem_n6598), .ZN(MEM_stage_inst_dmem_n6607) );
NAND2_X1 MEM_stage_inst_dmem_U6727 ( .A1(MEM_stage_inst_dmem_n6597), .A2(MEM_stage_inst_dmem_n6596), .ZN(MEM_stage_inst_dmem_n6598) );
NAND2_X1 MEM_stage_inst_dmem_U6726 ( .A1(MEM_stage_inst_dmem_ram_3308), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n6596) );
NAND2_X1 MEM_stage_inst_dmem_U6725 ( .A1(MEM_stage_inst_dmem_ram_3356), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n6597) );
NAND2_X1 MEM_stage_inst_dmem_U6724 ( .A1(MEM_stage_inst_dmem_n6595), .A2(MEM_stage_inst_dmem_n6594), .ZN(MEM_stage_inst_dmem_n6599) );
NAND2_X1 MEM_stage_inst_dmem_U6723 ( .A1(MEM_stage_inst_dmem_ram_3580), .A2(MEM_stage_inst_dmem_n64), .ZN(MEM_stage_inst_dmem_n6594) );
NAND2_X1 MEM_stage_inst_dmem_U6722 ( .A1(MEM_stage_inst_dmem_ram_3596), .A2(MEM_stage_inst_dmem_n8225), .ZN(MEM_stage_inst_dmem_n6595) );
NOR2_X1 MEM_stage_inst_dmem_U6721 ( .A1(MEM_stage_inst_dmem_n6593), .A2(MEM_stage_inst_dmem_n8551), .ZN(MEM_stage_inst_dmem_n6722) );
NOR2_X1 MEM_stage_inst_dmem_U6720 ( .A1(MEM_stage_inst_dmem_n6592), .A2(MEM_stage_inst_dmem_n6591), .ZN(MEM_stage_inst_dmem_n6593) );
NAND2_X1 MEM_stage_inst_dmem_U6719 ( .A1(MEM_stage_inst_dmem_n6590), .A2(MEM_stage_inst_dmem_n6589), .ZN(MEM_stage_inst_dmem_n6591) );
NOR2_X1 MEM_stage_inst_dmem_U6718 ( .A1(MEM_stage_inst_dmem_n6588), .A2(MEM_stage_inst_dmem_n6587), .ZN(MEM_stage_inst_dmem_n6589) );
NAND2_X1 MEM_stage_inst_dmem_U6717 ( .A1(MEM_stage_inst_dmem_n6586), .A2(MEM_stage_inst_dmem_n6585), .ZN(MEM_stage_inst_dmem_n6587) );
NOR2_X1 MEM_stage_inst_dmem_U6716 ( .A1(MEM_stage_inst_dmem_n6584), .A2(MEM_stage_inst_dmem_n6583), .ZN(MEM_stage_inst_dmem_n6585) );
NAND2_X1 MEM_stage_inst_dmem_U6715 ( .A1(MEM_stage_inst_dmem_n6582), .A2(MEM_stage_inst_dmem_n6581), .ZN(MEM_stage_inst_dmem_n6583) );
NAND2_X1 MEM_stage_inst_dmem_U6714 ( .A1(MEM_stage_inst_dmem_ram_412), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n6581) );
NAND2_X1 MEM_stage_inst_dmem_U6713 ( .A1(MEM_stage_inst_dmem_ram_172), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n6582) );
NAND2_X1 MEM_stage_inst_dmem_U6712 ( .A1(MEM_stage_inst_dmem_n6580), .A2(MEM_stage_inst_dmem_n6579), .ZN(MEM_stage_inst_dmem_n6584) );
NAND2_X1 MEM_stage_inst_dmem_U6711 ( .A1(MEM_stage_inst_dmem_ram_684), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n6579) );
NAND2_X1 MEM_stage_inst_dmem_U6710 ( .A1(MEM_stage_inst_dmem_ram_124), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n6580) );
NOR2_X1 MEM_stage_inst_dmem_U6709 ( .A1(MEM_stage_inst_dmem_n6578), .A2(MEM_stage_inst_dmem_n6577), .ZN(MEM_stage_inst_dmem_n6586) );
NAND2_X1 MEM_stage_inst_dmem_U6708 ( .A1(MEM_stage_inst_dmem_n6576), .A2(MEM_stage_inst_dmem_n6575), .ZN(MEM_stage_inst_dmem_n6577) );
NAND2_X1 MEM_stage_inst_dmem_U6707 ( .A1(MEM_stage_inst_dmem_ram_892), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n6575) );
NAND2_X1 MEM_stage_inst_dmem_U6706 ( .A1(MEM_stage_inst_dmem_ram_140), .A2(MEM_stage_inst_dmem_n8174), .ZN(MEM_stage_inst_dmem_n6576) );
NAND2_X1 MEM_stage_inst_dmem_U6705 ( .A1(MEM_stage_inst_dmem_n6574), .A2(MEM_stage_inst_dmem_n6573), .ZN(MEM_stage_inst_dmem_n6578) );
NAND2_X1 MEM_stage_inst_dmem_U6704 ( .A1(MEM_stage_inst_dmem_ram_780), .A2(MEM_stage_inst_dmem_n8472), .ZN(MEM_stage_inst_dmem_n6573) );
NAND2_X1 MEM_stage_inst_dmem_U6703 ( .A1(MEM_stage_inst_dmem_ram_156), .A2(MEM_stage_inst_dmem_n44), .ZN(MEM_stage_inst_dmem_n6574) );
NAND2_X1 MEM_stage_inst_dmem_U6702 ( .A1(MEM_stage_inst_dmem_n6572), .A2(MEM_stage_inst_dmem_n6571), .ZN(MEM_stage_inst_dmem_n6588) );
NOR2_X1 MEM_stage_inst_dmem_U6701 ( .A1(MEM_stage_inst_dmem_n6570), .A2(MEM_stage_inst_dmem_n6569), .ZN(MEM_stage_inst_dmem_n6571) );
NAND2_X1 MEM_stage_inst_dmem_U6700 ( .A1(MEM_stage_inst_dmem_n6568), .A2(MEM_stage_inst_dmem_n6567), .ZN(MEM_stage_inst_dmem_n6569) );
NAND2_X1 MEM_stage_inst_dmem_U6699 ( .A1(MEM_stage_inst_dmem_ram_812), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n6567) );
NAND2_X1 MEM_stage_inst_dmem_U6698 ( .A1(MEM_stage_inst_dmem_ram_268), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n6568) );
NAND2_X1 MEM_stage_inst_dmem_U6697 ( .A1(MEM_stage_inst_dmem_n6566), .A2(MEM_stage_inst_dmem_n6565), .ZN(MEM_stage_inst_dmem_n6570) );
NAND2_X1 MEM_stage_inst_dmem_U6696 ( .A1(MEM_stage_inst_dmem_ram_396), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n6565) );
NAND2_X1 MEM_stage_inst_dmem_U6695 ( .A1(MEM_stage_inst_dmem_ram_668), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n6566) );
NOR2_X1 MEM_stage_inst_dmem_U6694 ( .A1(MEM_stage_inst_dmem_n6564), .A2(MEM_stage_inst_dmem_n6563), .ZN(MEM_stage_inst_dmem_n6572) );
NAND2_X1 MEM_stage_inst_dmem_U6693 ( .A1(MEM_stage_inst_dmem_n6562), .A2(MEM_stage_inst_dmem_n6561), .ZN(MEM_stage_inst_dmem_n6563) );
NAND2_X1 MEM_stage_inst_dmem_U6692 ( .A1(MEM_stage_inst_dmem_ram_444), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n6561) );
NAND2_X1 MEM_stage_inst_dmem_U6691 ( .A1(MEM_stage_inst_dmem_ram_492), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n6562) );
NAND2_X1 MEM_stage_inst_dmem_U6690 ( .A1(MEM_stage_inst_dmem_n6560), .A2(MEM_stage_inst_dmem_n6559), .ZN(MEM_stage_inst_dmem_n6564) );
NAND2_X1 MEM_stage_inst_dmem_U6689 ( .A1(MEM_stage_inst_dmem_ram_764), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n6559) );
NAND2_X1 MEM_stage_inst_dmem_U6688 ( .A1(MEM_stage_inst_dmem_ram_700), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n6560) );
NOR2_X1 MEM_stage_inst_dmem_U6687 ( .A1(MEM_stage_inst_dmem_n6558), .A2(MEM_stage_inst_dmem_n6557), .ZN(MEM_stage_inst_dmem_n6590) );
NAND2_X1 MEM_stage_inst_dmem_U6686 ( .A1(MEM_stage_inst_dmem_n6556), .A2(MEM_stage_inst_dmem_n6555), .ZN(MEM_stage_inst_dmem_n6557) );
NOR2_X1 MEM_stage_inst_dmem_U6685 ( .A1(MEM_stage_inst_dmem_n6554), .A2(MEM_stage_inst_dmem_n6553), .ZN(MEM_stage_inst_dmem_n6555) );
NAND2_X1 MEM_stage_inst_dmem_U6684 ( .A1(MEM_stage_inst_dmem_n6552), .A2(MEM_stage_inst_dmem_n6551), .ZN(MEM_stage_inst_dmem_n6553) );
NAND2_X1 MEM_stage_inst_dmem_U6683 ( .A1(MEM_stage_inst_dmem_ram_204), .A2(MEM_stage_inst_dmem_n8256), .ZN(MEM_stage_inst_dmem_n6551) );
NAND2_X1 MEM_stage_inst_dmem_U6682 ( .A1(MEM_stage_inst_dmem_ram_28), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n6552) );
NAND2_X1 MEM_stage_inst_dmem_U6681 ( .A1(MEM_stage_inst_dmem_n6550), .A2(MEM_stage_inst_dmem_n6549), .ZN(MEM_stage_inst_dmem_n6554) );
NAND2_X1 MEM_stage_inst_dmem_U6680 ( .A1(MEM_stage_inst_dmem_ram_716), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n6549) );
NAND2_X1 MEM_stage_inst_dmem_U6679 ( .A1(MEM_stage_inst_dmem_ram_732), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n6550) );
NOR2_X1 MEM_stage_inst_dmem_U6678 ( .A1(MEM_stage_inst_dmem_n6548), .A2(MEM_stage_inst_dmem_n6547), .ZN(MEM_stage_inst_dmem_n6556) );
NAND2_X1 MEM_stage_inst_dmem_U6677 ( .A1(MEM_stage_inst_dmem_n6546), .A2(MEM_stage_inst_dmem_n6545), .ZN(MEM_stage_inst_dmem_n6547) );
NAND2_X1 MEM_stage_inst_dmem_U6676 ( .A1(MEM_stage_inst_dmem_ram_972), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n6545) );
NAND2_X1 MEM_stage_inst_dmem_U6675 ( .A1(MEM_stage_inst_dmem_ram_620), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n6546) );
NAND2_X1 MEM_stage_inst_dmem_U6674 ( .A1(MEM_stage_inst_dmem_n6544), .A2(MEM_stage_inst_dmem_n6543), .ZN(MEM_stage_inst_dmem_n6548) );
NAND2_X1 MEM_stage_inst_dmem_U6673 ( .A1(MEM_stage_inst_dmem_ram_988), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n6543) );
NAND2_X1 MEM_stage_inst_dmem_U6672 ( .A1(MEM_stage_inst_dmem_ram_524), .A2(MEM_stage_inst_dmem_n8225), .ZN(MEM_stage_inst_dmem_n6544) );
NAND2_X1 MEM_stage_inst_dmem_U6671 ( .A1(MEM_stage_inst_dmem_n6542), .A2(MEM_stage_inst_dmem_n6541), .ZN(MEM_stage_inst_dmem_n6558) );
NOR2_X1 MEM_stage_inst_dmem_U6670 ( .A1(MEM_stage_inst_dmem_n6540), .A2(MEM_stage_inst_dmem_n6539), .ZN(MEM_stage_inst_dmem_n6541) );
NAND2_X1 MEM_stage_inst_dmem_U6669 ( .A1(MEM_stage_inst_dmem_n6538), .A2(MEM_stage_inst_dmem_n6537), .ZN(MEM_stage_inst_dmem_n6539) );
NAND2_X1 MEM_stage_inst_dmem_U6668 ( .A1(MEM_stage_inst_dmem_ram_300), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n6537) );
NAND2_X1 MEM_stage_inst_dmem_U6667 ( .A1(MEM_stage_inst_dmem_ram_12), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n6538) );
NAND2_X1 MEM_stage_inst_dmem_U6666 ( .A1(MEM_stage_inst_dmem_n6536), .A2(MEM_stage_inst_dmem_n6535), .ZN(MEM_stage_inst_dmem_n6540) );
NAND2_X1 MEM_stage_inst_dmem_U6665 ( .A1(MEM_stage_inst_dmem_ram_76), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n6535) );
NAND2_X1 MEM_stage_inst_dmem_U6664 ( .A1(MEM_stage_inst_dmem_ram_476), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n6536) );
NOR2_X1 MEM_stage_inst_dmem_U6663 ( .A1(MEM_stage_inst_dmem_n6534), .A2(MEM_stage_inst_dmem_n6533), .ZN(MEM_stage_inst_dmem_n6542) );
NAND2_X1 MEM_stage_inst_dmem_U6662 ( .A1(MEM_stage_inst_dmem_n6532), .A2(MEM_stage_inst_dmem_n6531), .ZN(MEM_stage_inst_dmem_n6533) );
NAND2_X1 MEM_stage_inst_dmem_U6661 ( .A1(MEM_stage_inst_dmem_ram_364), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n6531) );
NAND2_X1 MEM_stage_inst_dmem_U6660 ( .A1(MEM_stage_inst_dmem_ram_636), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n6532) );
NAND2_X1 MEM_stage_inst_dmem_U6659 ( .A1(MEM_stage_inst_dmem_n6530), .A2(MEM_stage_inst_dmem_n6529), .ZN(MEM_stage_inst_dmem_n6534) );
NAND2_X1 MEM_stage_inst_dmem_U6658 ( .A1(MEM_stage_inst_dmem_ram_860), .A2(MEM_stage_inst_dmem_n3141), .ZN(MEM_stage_inst_dmem_n6529) );
NAND2_X1 MEM_stage_inst_dmem_U6657 ( .A1(MEM_stage_inst_dmem_ram_460), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n6530) );
NAND2_X1 MEM_stage_inst_dmem_U6656 ( .A1(MEM_stage_inst_dmem_n6528), .A2(MEM_stage_inst_dmem_n6527), .ZN(MEM_stage_inst_dmem_n6592) );
NOR2_X1 MEM_stage_inst_dmem_U6655 ( .A1(MEM_stage_inst_dmem_n6526), .A2(MEM_stage_inst_dmem_n6525), .ZN(MEM_stage_inst_dmem_n6527) );
NAND2_X1 MEM_stage_inst_dmem_U6654 ( .A1(MEM_stage_inst_dmem_n6524), .A2(MEM_stage_inst_dmem_n6523), .ZN(MEM_stage_inst_dmem_n6525) );
NOR2_X1 MEM_stage_inst_dmem_U6653 ( .A1(MEM_stage_inst_dmem_n6522), .A2(MEM_stage_inst_dmem_n6521), .ZN(MEM_stage_inst_dmem_n6523) );
NAND2_X1 MEM_stage_inst_dmem_U6652 ( .A1(MEM_stage_inst_dmem_n6520), .A2(MEM_stage_inst_dmem_n6519), .ZN(MEM_stage_inst_dmem_n6521) );
NAND2_X1 MEM_stage_inst_dmem_U6651 ( .A1(MEM_stage_inst_dmem_ram_540), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n6519) );
NAND2_X1 MEM_stage_inst_dmem_U6650 ( .A1(MEM_stage_inst_dmem_ram_748), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n6520) );
NAND2_X1 MEM_stage_inst_dmem_U6649 ( .A1(MEM_stage_inst_dmem_n6518), .A2(MEM_stage_inst_dmem_n6517), .ZN(MEM_stage_inst_dmem_n6522) );
NAND2_X1 MEM_stage_inst_dmem_U6648 ( .A1(MEM_stage_inst_dmem_ram_316), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n6517) );
NAND2_X1 MEM_stage_inst_dmem_U6647 ( .A1(MEM_stage_inst_dmem_ram_604), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n6518) );
NOR2_X1 MEM_stage_inst_dmem_U6646 ( .A1(MEM_stage_inst_dmem_n6516), .A2(MEM_stage_inst_dmem_n6515), .ZN(MEM_stage_inst_dmem_n6524) );
NAND2_X1 MEM_stage_inst_dmem_U6645 ( .A1(MEM_stage_inst_dmem_n6514), .A2(MEM_stage_inst_dmem_n6513), .ZN(MEM_stage_inst_dmem_n6515) );
NAND2_X1 MEM_stage_inst_dmem_U6644 ( .A1(MEM_stage_inst_dmem_ram_572), .A2(MEM_stage_inst_dmem_n8169), .ZN(MEM_stage_inst_dmem_n6513) );
NAND2_X1 MEM_stage_inst_dmem_U6643 ( .A1(MEM_stage_inst_dmem_ram_284), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n6514) );
NAND2_X1 MEM_stage_inst_dmem_U6642 ( .A1(MEM_stage_inst_dmem_n6512), .A2(MEM_stage_inst_dmem_n6511), .ZN(MEM_stage_inst_dmem_n6516) );
NAND2_X1 MEM_stage_inst_dmem_U6641 ( .A1(MEM_stage_inst_dmem_ram_908), .A2(MEM_stage_inst_dmem_n8193), .ZN(MEM_stage_inst_dmem_n6511) );
NAND2_X1 MEM_stage_inst_dmem_U6640 ( .A1(MEM_stage_inst_dmem_ram_92), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n6512) );
NAND2_X1 MEM_stage_inst_dmem_U6639 ( .A1(MEM_stage_inst_dmem_n6510), .A2(MEM_stage_inst_dmem_n6509), .ZN(MEM_stage_inst_dmem_n6526) );
NOR2_X1 MEM_stage_inst_dmem_U6638 ( .A1(MEM_stage_inst_dmem_n6508), .A2(MEM_stage_inst_dmem_n6507), .ZN(MEM_stage_inst_dmem_n6509) );
NAND2_X1 MEM_stage_inst_dmem_U6637 ( .A1(MEM_stage_inst_dmem_n6506), .A2(MEM_stage_inst_dmem_n6505), .ZN(MEM_stage_inst_dmem_n6507) );
NAND2_X1 MEM_stage_inst_dmem_U6636 ( .A1(MEM_stage_inst_dmem_ram_1020), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n6505) );
NAND2_X1 MEM_stage_inst_dmem_U6635 ( .A1(MEM_stage_inst_dmem_ram_940), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n6506) );
NAND2_X1 MEM_stage_inst_dmem_U6634 ( .A1(MEM_stage_inst_dmem_n6504), .A2(MEM_stage_inst_dmem_n6503), .ZN(MEM_stage_inst_dmem_n6508) );
NAND2_X1 MEM_stage_inst_dmem_U6633 ( .A1(MEM_stage_inst_dmem_ram_956), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n6503) );
NAND2_X1 MEM_stage_inst_dmem_U6632 ( .A1(MEM_stage_inst_dmem_ram_924), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n6504) );
NOR2_X1 MEM_stage_inst_dmem_U6631 ( .A1(MEM_stage_inst_dmem_n6502), .A2(MEM_stage_inst_dmem_n6501), .ZN(MEM_stage_inst_dmem_n6510) );
NAND2_X1 MEM_stage_inst_dmem_U6630 ( .A1(MEM_stage_inst_dmem_n6500), .A2(MEM_stage_inst_dmem_n6499), .ZN(MEM_stage_inst_dmem_n6501) );
NAND2_X1 MEM_stage_inst_dmem_U6629 ( .A1(MEM_stage_inst_dmem_ram_332), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n6499) );
NAND2_X1 MEM_stage_inst_dmem_U6628 ( .A1(MEM_stage_inst_dmem_ram_844), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n6500) );
NAND2_X1 MEM_stage_inst_dmem_U6627 ( .A1(MEM_stage_inst_dmem_n6498), .A2(MEM_stage_inst_dmem_n6497), .ZN(MEM_stage_inst_dmem_n6502) );
NAND2_X1 MEM_stage_inst_dmem_U6626 ( .A1(MEM_stage_inst_dmem_ram_108), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n6497) );
NAND2_X1 MEM_stage_inst_dmem_U6625 ( .A1(MEM_stage_inst_dmem_ram_588), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n6498) );
NOR2_X1 MEM_stage_inst_dmem_U6624 ( .A1(MEM_stage_inst_dmem_n6496), .A2(MEM_stage_inst_dmem_n6495), .ZN(MEM_stage_inst_dmem_n6528) );
NAND2_X1 MEM_stage_inst_dmem_U6623 ( .A1(MEM_stage_inst_dmem_n6494), .A2(MEM_stage_inst_dmem_n6493), .ZN(MEM_stage_inst_dmem_n6495) );
NOR2_X1 MEM_stage_inst_dmem_U6622 ( .A1(MEM_stage_inst_dmem_n6492), .A2(MEM_stage_inst_dmem_n6491), .ZN(MEM_stage_inst_dmem_n6493) );
NAND2_X1 MEM_stage_inst_dmem_U6621 ( .A1(MEM_stage_inst_dmem_n6490), .A2(MEM_stage_inst_dmem_n6489), .ZN(MEM_stage_inst_dmem_n6491) );
NAND2_X1 MEM_stage_inst_dmem_U6620 ( .A1(MEM_stage_inst_dmem_ram_508), .A2(MEM_stage_inst_dmem_n64), .ZN(MEM_stage_inst_dmem_n6489) );
NAND2_X1 MEM_stage_inst_dmem_U6619 ( .A1(MEM_stage_inst_dmem_ram_556), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n6490) );
NAND2_X1 MEM_stage_inst_dmem_U6618 ( .A1(MEM_stage_inst_dmem_n6488), .A2(MEM_stage_inst_dmem_n6487), .ZN(MEM_stage_inst_dmem_n6492) );
NAND2_X1 MEM_stage_inst_dmem_U6617 ( .A1(MEM_stage_inst_dmem_ram_428), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n6487) );
NAND2_X1 MEM_stage_inst_dmem_U6616 ( .A1(MEM_stage_inst_dmem_ram_44), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n6488) );
NOR2_X1 MEM_stage_inst_dmem_U6615 ( .A1(MEM_stage_inst_dmem_n6486), .A2(MEM_stage_inst_dmem_n6485), .ZN(MEM_stage_inst_dmem_n6494) );
NAND2_X1 MEM_stage_inst_dmem_U6614 ( .A1(MEM_stage_inst_dmem_n6484), .A2(MEM_stage_inst_dmem_n6483), .ZN(MEM_stage_inst_dmem_n6485) );
NAND2_X1 MEM_stage_inst_dmem_U6613 ( .A1(MEM_stage_inst_dmem_ram_60), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n6483) );
NAND2_X1 MEM_stage_inst_dmem_U6612 ( .A1(MEM_stage_inst_dmem_ram_828), .A2(MEM_stage_inst_dmem_n8005), .ZN(MEM_stage_inst_dmem_n6484) );
NAND2_X1 MEM_stage_inst_dmem_U6611 ( .A1(MEM_stage_inst_dmem_n6482), .A2(MEM_stage_inst_dmem_n6481), .ZN(MEM_stage_inst_dmem_n6486) );
NAND2_X1 MEM_stage_inst_dmem_U6610 ( .A1(MEM_stage_inst_dmem_ram_188), .A2(MEM_stage_inst_dmem_n8434), .ZN(MEM_stage_inst_dmem_n6481) );
NAND2_X1 MEM_stage_inst_dmem_U6609 ( .A1(MEM_stage_inst_dmem_ram_380), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n6482) );
NAND2_X1 MEM_stage_inst_dmem_U6608 ( .A1(MEM_stage_inst_dmem_n6480), .A2(MEM_stage_inst_dmem_n6479), .ZN(MEM_stage_inst_dmem_n6496) );
NOR2_X1 MEM_stage_inst_dmem_U6607 ( .A1(MEM_stage_inst_dmem_n6478), .A2(MEM_stage_inst_dmem_n6477), .ZN(MEM_stage_inst_dmem_n6479) );
NAND2_X1 MEM_stage_inst_dmem_U6606 ( .A1(MEM_stage_inst_dmem_n6476), .A2(MEM_stage_inst_dmem_n6475), .ZN(MEM_stage_inst_dmem_n6477) );
NAND2_X1 MEM_stage_inst_dmem_U6605 ( .A1(MEM_stage_inst_dmem_ram_876), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n6475) );
NAND2_X1 MEM_stage_inst_dmem_U6604 ( .A1(MEM_stage_inst_dmem_ram_252), .A2(MEM_stage_inst_dmem_n7914), .ZN(MEM_stage_inst_dmem_n6476) );
NAND2_X1 MEM_stage_inst_dmem_U6603 ( .A1(MEM_stage_inst_dmem_n6474), .A2(MEM_stage_inst_dmem_n6473), .ZN(MEM_stage_inst_dmem_n6478) );
NAND2_X1 MEM_stage_inst_dmem_U6602 ( .A1(MEM_stage_inst_dmem_ram_1004), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n6473) );
NAND2_X1 MEM_stage_inst_dmem_U6601 ( .A1(MEM_stage_inst_dmem_ram_348), .A2(MEM_stage_inst_dmem_n3216), .ZN(MEM_stage_inst_dmem_n6474) );
NOR2_X1 MEM_stage_inst_dmem_U6600 ( .A1(MEM_stage_inst_dmem_n6472), .A2(MEM_stage_inst_dmem_n6471), .ZN(MEM_stage_inst_dmem_n6480) );
NAND2_X1 MEM_stage_inst_dmem_U6599 ( .A1(MEM_stage_inst_dmem_n6470), .A2(MEM_stage_inst_dmem_n6469), .ZN(MEM_stage_inst_dmem_n6471) );
NAND2_X1 MEM_stage_inst_dmem_U6598 ( .A1(MEM_stage_inst_dmem_ram_652), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n6469) );
NAND2_X1 MEM_stage_inst_dmem_U6597 ( .A1(MEM_stage_inst_dmem_ram_220), .A2(MEM_stage_inst_dmem_n8206), .ZN(MEM_stage_inst_dmem_n6470) );
NAND2_X1 MEM_stage_inst_dmem_U6596 ( .A1(MEM_stage_inst_dmem_n6468), .A2(MEM_stage_inst_dmem_n6467), .ZN(MEM_stage_inst_dmem_n6472) );
NAND2_X1 MEM_stage_inst_dmem_U6595 ( .A1(MEM_stage_inst_dmem_ram_236), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n6467) );
NAND2_X1 MEM_stage_inst_dmem_U6594 ( .A1(MEM_stage_inst_dmem_ram_796), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n6468) );
NAND2_X1 MEM_stage_inst_dmem_U6593 ( .A1(MEM_stage_inst_dmem_n6466), .A2(MEM_stage_inst_dmem_n6465), .ZN(MEM_stage_inst_mem_read_data_11) );
NOR2_X1 MEM_stage_inst_dmem_U6592 ( .A1(MEM_stage_inst_dmem_n6464), .A2(MEM_stage_inst_dmem_n6463), .ZN(MEM_stage_inst_dmem_n6465) );
NOR2_X1 MEM_stage_inst_dmem_U6591 ( .A1(MEM_stage_inst_dmem_n6462), .A2(MEM_stage_inst_dmem_n8286), .ZN(MEM_stage_inst_dmem_n6463) );
NOR2_X1 MEM_stage_inst_dmem_U6590 ( .A1(MEM_stage_inst_dmem_n6461), .A2(MEM_stage_inst_dmem_n6460), .ZN(MEM_stage_inst_dmem_n6462) );
NAND2_X1 MEM_stage_inst_dmem_U6589 ( .A1(MEM_stage_inst_dmem_n6459), .A2(MEM_stage_inst_dmem_n6458), .ZN(MEM_stage_inst_dmem_n6460) );
NOR2_X1 MEM_stage_inst_dmem_U6588 ( .A1(MEM_stage_inst_dmem_n6457), .A2(MEM_stage_inst_dmem_n6456), .ZN(MEM_stage_inst_dmem_n6458) );
NAND2_X1 MEM_stage_inst_dmem_U6587 ( .A1(MEM_stage_inst_dmem_n6455), .A2(MEM_stage_inst_dmem_n6454), .ZN(MEM_stage_inst_dmem_n6456) );
NOR2_X1 MEM_stage_inst_dmem_U6586 ( .A1(MEM_stage_inst_dmem_n6453), .A2(MEM_stage_inst_dmem_n6452), .ZN(MEM_stage_inst_dmem_n6454) );
NAND2_X1 MEM_stage_inst_dmem_U6585 ( .A1(MEM_stage_inst_dmem_n6451), .A2(MEM_stage_inst_dmem_n6450), .ZN(MEM_stage_inst_dmem_n6452) );
NAND2_X1 MEM_stage_inst_dmem_U6584 ( .A1(MEM_stage_inst_dmem_ram_2907), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n6450) );
NAND2_X1 MEM_stage_inst_dmem_U6583 ( .A1(MEM_stage_inst_dmem_ram_2315), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n6451) );
NAND2_X1 MEM_stage_inst_dmem_U6582 ( .A1(MEM_stage_inst_dmem_n6449), .A2(MEM_stage_inst_dmem_n6448), .ZN(MEM_stage_inst_dmem_n6453) );
NAND2_X1 MEM_stage_inst_dmem_U6581 ( .A1(MEM_stage_inst_dmem_ram_2203), .A2(MEM_stage_inst_dmem_n44), .ZN(MEM_stage_inst_dmem_n6448) );
NAND2_X1 MEM_stage_inst_dmem_U6580 ( .A1(MEM_stage_inst_dmem_ram_2779), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n6449) );
NOR2_X1 MEM_stage_inst_dmem_U6579 ( .A1(MEM_stage_inst_dmem_n6447), .A2(MEM_stage_inst_dmem_n6446), .ZN(MEM_stage_inst_dmem_n6455) );
NAND2_X1 MEM_stage_inst_dmem_U6578 ( .A1(MEM_stage_inst_dmem_n6445), .A2(MEM_stage_inst_dmem_n6444), .ZN(MEM_stage_inst_dmem_n6446) );
NAND2_X1 MEM_stage_inst_dmem_U6577 ( .A1(MEM_stage_inst_dmem_ram_2603), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n6444) );
NAND2_X1 MEM_stage_inst_dmem_U6576 ( .A1(MEM_stage_inst_dmem_ram_2571), .A2(MEM_stage_inst_dmem_n8225), .ZN(MEM_stage_inst_dmem_n6445) );
NAND2_X1 MEM_stage_inst_dmem_U6575 ( .A1(MEM_stage_inst_dmem_n6443), .A2(MEM_stage_inst_dmem_n6442), .ZN(MEM_stage_inst_dmem_n6447) );
NAND2_X1 MEM_stage_inst_dmem_U6574 ( .A1(MEM_stage_inst_dmem_ram_2939), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n6442) );
NAND2_X1 MEM_stage_inst_dmem_U6573 ( .A1(MEM_stage_inst_dmem_ram_2267), .A2(MEM_stage_inst_dmem_n8206), .ZN(MEM_stage_inst_dmem_n6443) );
NAND2_X1 MEM_stage_inst_dmem_U6572 ( .A1(MEM_stage_inst_dmem_n6441), .A2(MEM_stage_inst_dmem_n6440), .ZN(MEM_stage_inst_dmem_n6457) );
NOR2_X1 MEM_stage_inst_dmem_U6571 ( .A1(MEM_stage_inst_dmem_n6439), .A2(MEM_stage_inst_dmem_n6438), .ZN(MEM_stage_inst_dmem_n6440) );
NAND2_X1 MEM_stage_inst_dmem_U6570 ( .A1(MEM_stage_inst_dmem_n6437), .A2(MEM_stage_inst_dmem_n6436), .ZN(MEM_stage_inst_dmem_n6438) );
NAND2_X1 MEM_stage_inst_dmem_U6569 ( .A1(MEM_stage_inst_dmem_ram_3019), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n6436) );
NAND2_X1 MEM_stage_inst_dmem_U6568 ( .A1(MEM_stage_inst_dmem_ram_2075), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n6437) );
NAND2_X1 MEM_stage_inst_dmem_U6567 ( .A1(MEM_stage_inst_dmem_n6435), .A2(MEM_stage_inst_dmem_n6434), .ZN(MEM_stage_inst_dmem_n6439) );
NAND2_X1 MEM_stage_inst_dmem_U6566 ( .A1(MEM_stage_inst_dmem_ram_2971), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n6434) );
NAND2_X1 MEM_stage_inst_dmem_U6565 ( .A1(MEM_stage_inst_dmem_ram_2635), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n6435) );
NOR2_X1 MEM_stage_inst_dmem_U6564 ( .A1(MEM_stage_inst_dmem_n6433), .A2(MEM_stage_inst_dmem_n6432), .ZN(MEM_stage_inst_dmem_n6441) );
NAND2_X1 MEM_stage_inst_dmem_U6563 ( .A1(MEM_stage_inst_dmem_n6431), .A2(MEM_stage_inst_dmem_n6430), .ZN(MEM_stage_inst_dmem_n6432) );
NAND2_X1 MEM_stage_inst_dmem_U6562 ( .A1(MEM_stage_inst_dmem_ram_2587), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n6430) );
NAND2_X1 MEM_stage_inst_dmem_U6561 ( .A1(MEM_stage_inst_dmem_ram_2651), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n6431) );
NAND2_X1 MEM_stage_inst_dmem_U6560 ( .A1(MEM_stage_inst_dmem_n6429), .A2(MEM_stage_inst_dmem_n6428), .ZN(MEM_stage_inst_dmem_n6433) );
NAND2_X1 MEM_stage_inst_dmem_U6559 ( .A1(MEM_stage_inst_dmem_ram_2923), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n6428) );
NAND2_X1 MEM_stage_inst_dmem_U6558 ( .A1(MEM_stage_inst_dmem_ram_2283), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n6429) );
NOR2_X1 MEM_stage_inst_dmem_U6557 ( .A1(MEM_stage_inst_dmem_n6427), .A2(MEM_stage_inst_dmem_n6426), .ZN(MEM_stage_inst_dmem_n6459) );
NAND2_X1 MEM_stage_inst_dmem_U6556 ( .A1(MEM_stage_inst_dmem_n6425), .A2(MEM_stage_inst_dmem_n6424), .ZN(MEM_stage_inst_dmem_n6426) );
NOR2_X1 MEM_stage_inst_dmem_U6555 ( .A1(MEM_stage_inst_dmem_n6423), .A2(MEM_stage_inst_dmem_n6422), .ZN(MEM_stage_inst_dmem_n6424) );
NAND2_X1 MEM_stage_inst_dmem_U6554 ( .A1(MEM_stage_inst_dmem_n6421), .A2(MEM_stage_inst_dmem_n6420), .ZN(MEM_stage_inst_dmem_n6422) );
NAND2_X1 MEM_stage_inst_dmem_U6553 ( .A1(MEM_stage_inst_dmem_ram_2891), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n6420) );
NAND2_X1 MEM_stage_inst_dmem_U6552 ( .A1(MEM_stage_inst_dmem_ram_2059), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n6421) );
NAND2_X1 MEM_stage_inst_dmem_U6551 ( .A1(MEM_stage_inst_dmem_n6419), .A2(MEM_stage_inst_dmem_n6418), .ZN(MEM_stage_inst_dmem_n6423) );
NAND2_X1 MEM_stage_inst_dmem_U6550 ( .A1(MEM_stage_inst_dmem_ram_2459), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n6418) );
NAND2_X1 MEM_stage_inst_dmem_U6549 ( .A1(MEM_stage_inst_dmem_ram_2859), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n6419) );
NOR2_X1 MEM_stage_inst_dmem_U6548 ( .A1(MEM_stage_inst_dmem_n6417), .A2(MEM_stage_inst_dmem_n6416), .ZN(MEM_stage_inst_dmem_n6425) );
NAND2_X1 MEM_stage_inst_dmem_U6547 ( .A1(MEM_stage_inst_dmem_n6415), .A2(MEM_stage_inst_dmem_n6414), .ZN(MEM_stage_inst_dmem_n6416) );
NAND2_X1 MEM_stage_inst_dmem_U6546 ( .A1(MEM_stage_inst_dmem_ram_2187), .A2(MEM_stage_inst_dmem_n8174), .ZN(MEM_stage_inst_dmem_n6414) );
NAND2_X1 MEM_stage_inst_dmem_U6545 ( .A1(MEM_stage_inst_dmem_ram_2875), .A2(MEM_stage_inst_dmem_n46), .ZN(MEM_stage_inst_dmem_n6415) );
NAND2_X1 MEM_stage_inst_dmem_U6544 ( .A1(MEM_stage_inst_dmem_n6413), .A2(MEM_stage_inst_dmem_n6412), .ZN(MEM_stage_inst_dmem_n6417) );
NAND2_X1 MEM_stage_inst_dmem_U6543 ( .A1(MEM_stage_inst_dmem_ram_2251), .A2(MEM_stage_inst_dmem_n8256), .ZN(MEM_stage_inst_dmem_n6412) );
NAND2_X1 MEM_stage_inst_dmem_U6542 ( .A1(MEM_stage_inst_dmem_ram_2987), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n6413) );
NAND2_X1 MEM_stage_inst_dmem_U6541 ( .A1(MEM_stage_inst_dmem_n6411), .A2(MEM_stage_inst_dmem_n6410), .ZN(MEM_stage_inst_dmem_n6427) );
NOR2_X1 MEM_stage_inst_dmem_U6540 ( .A1(MEM_stage_inst_dmem_n6409), .A2(MEM_stage_inst_dmem_n6408), .ZN(MEM_stage_inst_dmem_n6410) );
NAND2_X1 MEM_stage_inst_dmem_U6539 ( .A1(MEM_stage_inst_dmem_n6407), .A2(MEM_stage_inst_dmem_n6406), .ZN(MEM_stage_inst_dmem_n6408) );
NAND2_X1 MEM_stage_inst_dmem_U6538 ( .A1(MEM_stage_inst_dmem_ram_2475), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n6406) );
NAND2_X1 MEM_stage_inst_dmem_U6537 ( .A1(MEM_stage_inst_dmem_ram_2683), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n6407) );
NAND2_X1 MEM_stage_inst_dmem_U6536 ( .A1(MEM_stage_inst_dmem_n6405), .A2(MEM_stage_inst_dmem_n6404), .ZN(MEM_stage_inst_dmem_n6409) );
NAND2_X1 MEM_stage_inst_dmem_U6535 ( .A1(MEM_stage_inst_dmem_ram_2219), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n6404) );
NAND2_X1 MEM_stage_inst_dmem_U6534 ( .A1(MEM_stage_inst_dmem_ram_2427), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n6405) );
NOR2_X1 MEM_stage_inst_dmem_U6533 ( .A1(MEM_stage_inst_dmem_n6403), .A2(MEM_stage_inst_dmem_n6402), .ZN(MEM_stage_inst_dmem_n6411) );
NAND2_X1 MEM_stage_inst_dmem_U6532 ( .A1(MEM_stage_inst_dmem_n6401), .A2(MEM_stage_inst_dmem_n6400), .ZN(MEM_stage_inst_dmem_n6402) );
NAND2_X1 MEM_stage_inst_dmem_U6531 ( .A1(MEM_stage_inst_dmem_ram_2763), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n6400) );
NAND2_X1 MEM_stage_inst_dmem_U6530 ( .A1(MEM_stage_inst_dmem_ram_2667), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n6401) );
NAND2_X1 MEM_stage_inst_dmem_U6529 ( .A1(MEM_stage_inst_dmem_n6399), .A2(MEM_stage_inst_dmem_n6398), .ZN(MEM_stage_inst_dmem_n6403) );
NAND2_X1 MEM_stage_inst_dmem_U6528 ( .A1(MEM_stage_inst_dmem_ram_2827), .A2(MEM_stage_inst_dmem_n8472), .ZN(MEM_stage_inst_dmem_n6398) );
NAND2_X1 MEM_stage_inst_dmem_U6527 ( .A1(MEM_stage_inst_dmem_ram_2491), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n6399) );
NAND2_X1 MEM_stage_inst_dmem_U6526 ( .A1(MEM_stage_inst_dmem_n6397), .A2(MEM_stage_inst_dmem_n6396), .ZN(MEM_stage_inst_dmem_n6461) );
NOR2_X1 MEM_stage_inst_dmem_U6525 ( .A1(MEM_stage_inst_dmem_n6395), .A2(MEM_stage_inst_dmem_n6394), .ZN(MEM_stage_inst_dmem_n6396) );
NAND2_X1 MEM_stage_inst_dmem_U6524 ( .A1(MEM_stage_inst_dmem_n6393), .A2(MEM_stage_inst_dmem_n6392), .ZN(MEM_stage_inst_dmem_n6394) );
NOR2_X1 MEM_stage_inst_dmem_U6523 ( .A1(MEM_stage_inst_dmem_n6391), .A2(MEM_stage_inst_dmem_n6390), .ZN(MEM_stage_inst_dmem_n6392) );
NAND2_X1 MEM_stage_inst_dmem_U6522 ( .A1(MEM_stage_inst_dmem_n6389), .A2(MEM_stage_inst_dmem_n6388), .ZN(MEM_stage_inst_dmem_n6390) );
NAND2_X1 MEM_stage_inst_dmem_U6521 ( .A1(MEM_stage_inst_dmem_ram_2619), .A2(MEM_stage_inst_dmem_n8169), .ZN(MEM_stage_inst_dmem_n6388) );
NAND2_X1 MEM_stage_inst_dmem_U6520 ( .A1(MEM_stage_inst_dmem_ram_2811), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n6389) );
NAND2_X1 MEM_stage_inst_dmem_U6519 ( .A1(MEM_stage_inst_dmem_n6387), .A2(MEM_stage_inst_dmem_n6386), .ZN(MEM_stage_inst_dmem_n6391) );
NAND2_X1 MEM_stage_inst_dmem_U6518 ( .A1(MEM_stage_inst_dmem_ram_2699), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n6386) );
NAND2_X1 MEM_stage_inst_dmem_U6517 ( .A1(MEM_stage_inst_dmem_ram_2507), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n6387) );
NOR2_X1 MEM_stage_inst_dmem_U6516 ( .A1(MEM_stage_inst_dmem_n6385), .A2(MEM_stage_inst_dmem_n6384), .ZN(MEM_stage_inst_dmem_n6393) );
NAND2_X1 MEM_stage_inst_dmem_U6515 ( .A1(MEM_stage_inst_dmem_n6383), .A2(MEM_stage_inst_dmem_n6382), .ZN(MEM_stage_inst_dmem_n6384) );
NAND2_X1 MEM_stage_inst_dmem_U6514 ( .A1(MEM_stage_inst_dmem_ram_2363), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n6382) );
NAND2_X1 MEM_stage_inst_dmem_U6513 ( .A1(MEM_stage_inst_dmem_ram_2123), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n6383) );
NAND2_X1 MEM_stage_inst_dmem_U6512 ( .A1(MEM_stage_inst_dmem_n6381), .A2(MEM_stage_inst_dmem_n6380), .ZN(MEM_stage_inst_dmem_n6385) );
NAND2_X1 MEM_stage_inst_dmem_U6511 ( .A1(MEM_stage_inst_dmem_ram_2331), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n6380) );
NAND2_X1 MEM_stage_inst_dmem_U6510 ( .A1(MEM_stage_inst_dmem_ram_2171), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n6381) );
NAND2_X1 MEM_stage_inst_dmem_U6509 ( .A1(MEM_stage_inst_dmem_n6379), .A2(MEM_stage_inst_dmem_n6378), .ZN(MEM_stage_inst_dmem_n6395) );
NOR2_X1 MEM_stage_inst_dmem_U6508 ( .A1(MEM_stage_inst_dmem_n6377), .A2(MEM_stage_inst_dmem_n6376), .ZN(MEM_stage_inst_dmem_n6378) );
NAND2_X1 MEM_stage_inst_dmem_U6507 ( .A1(MEM_stage_inst_dmem_n6375), .A2(MEM_stage_inst_dmem_n6374), .ZN(MEM_stage_inst_dmem_n6376) );
NAND2_X1 MEM_stage_inst_dmem_U6506 ( .A1(MEM_stage_inst_dmem_ram_2411), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n6374) );
NAND2_X1 MEM_stage_inst_dmem_U6505 ( .A1(MEM_stage_inst_dmem_ram_3067), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n6375) );
NAND2_X1 MEM_stage_inst_dmem_U6504 ( .A1(MEM_stage_inst_dmem_n6373), .A2(MEM_stage_inst_dmem_n6372), .ZN(MEM_stage_inst_dmem_n6377) );
NAND2_X1 MEM_stage_inst_dmem_U6503 ( .A1(MEM_stage_inst_dmem_ram_2555), .A2(MEM_stage_inst_dmem_n64), .ZN(MEM_stage_inst_dmem_n6372) );
NAND2_X1 MEM_stage_inst_dmem_U6502 ( .A1(MEM_stage_inst_dmem_ram_2523), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n6373) );
NOR2_X1 MEM_stage_inst_dmem_U6501 ( .A1(MEM_stage_inst_dmem_n6371), .A2(MEM_stage_inst_dmem_n6370), .ZN(MEM_stage_inst_dmem_n6379) );
NAND2_X1 MEM_stage_inst_dmem_U6500 ( .A1(MEM_stage_inst_dmem_n6369), .A2(MEM_stage_inst_dmem_n6368), .ZN(MEM_stage_inst_dmem_n6370) );
NAND2_X1 MEM_stage_inst_dmem_U6499 ( .A1(MEM_stage_inst_dmem_ram_2091), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n6368) );
NAND2_X1 MEM_stage_inst_dmem_U6498 ( .A1(MEM_stage_inst_dmem_ram_2715), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n6369) );
NAND2_X1 MEM_stage_inst_dmem_U6497 ( .A1(MEM_stage_inst_dmem_n6367), .A2(MEM_stage_inst_dmem_n6366), .ZN(MEM_stage_inst_dmem_n6371) );
NAND2_X1 MEM_stage_inst_dmem_U6496 ( .A1(MEM_stage_inst_dmem_ram_2107), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n6366) );
NAND2_X1 MEM_stage_inst_dmem_U6495 ( .A1(MEM_stage_inst_dmem_ram_2235), .A2(MEM_stage_inst_dmem_n8434), .ZN(MEM_stage_inst_dmem_n6367) );
NOR2_X1 MEM_stage_inst_dmem_U6494 ( .A1(MEM_stage_inst_dmem_n6365), .A2(MEM_stage_inst_dmem_n6364), .ZN(MEM_stage_inst_dmem_n6397) );
NAND2_X1 MEM_stage_inst_dmem_U6493 ( .A1(MEM_stage_inst_dmem_n6363), .A2(MEM_stage_inst_dmem_n6362), .ZN(MEM_stage_inst_dmem_n6364) );
NOR2_X1 MEM_stage_inst_dmem_U6492 ( .A1(MEM_stage_inst_dmem_n6361), .A2(MEM_stage_inst_dmem_n6360), .ZN(MEM_stage_inst_dmem_n6362) );
NAND2_X1 MEM_stage_inst_dmem_U6491 ( .A1(MEM_stage_inst_dmem_n6359), .A2(MEM_stage_inst_dmem_n6358), .ZN(MEM_stage_inst_dmem_n6360) );
NAND2_X1 MEM_stage_inst_dmem_U6490 ( .A1(MEM_stage_inst_dmem_ram_2139), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n6358) );
NAND2_X1 MEM_stage_inst_dmem_U6489 ( .A1(MEM_stage_inst_dmem_ram_2347), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n6359) );
NAND2_X1 MEM_stage_inst_dmem_U6488 ( .A1(MEM_stage_inst_dmem_n6357), .A2(MEM_stage_inst_dmem_n6356), .ZN(MEM_stage_inst_dmem_n6361) );
NAND2_X1 MEM_stage_inst_dmem_U6487 ( .A1(MEM_stage_inst_dmem_ram_2443), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n6356) );
NAND2_X1 MEM_stage_inst_dmem_U6486 ( .A1(MEM_stage_inst_dmem_ram_2843), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n6357) );
NOR2_X1 MEM_stage_inst_dmem_U6485 ( .A1(MEM_stage_inst_dmem_n6355), .A2(MEM_stage_inst_dmem_n6354), .ZN(MEM_stage_inst_dmem_n6363) );
NAND2_X1 MEM_stage_inst_dmem_U6484 ( .A1(MEM_stage_inst_dmem_n6353), .A2(MEM_stage_inst_dmem_n6352), .ZN(MEM_stage_inst_dmem_n6354) );
NAND2_X1 MEM_stage_inst_dmem_U6483 ( .A1(MEM_stage_inst_dmem_ram_3003), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n6352) );
NAND2_X1 MEM_stage_inst_dmem_U6482 ( .A1(MEM_stage_inst_dmem_ram_3051), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n6353) );
NAND2_X1 MEM_stage_inst_dmem_U6481 ( .A1(MEM_stage_inst_dmem_n6351), .A2(MEM_stage_inst_dmem_n6350), .ZN(MEM_stage_inst_dmem_n6355) );
NAND2_X1 MEM_stage_inst_dmem_U6480 ( .A1(MEM_stage_inst_dmem_ram_2299), .A2(MEM_stage_inst_dmem_n39), .ZN(MEM_stage_inst_dmem_n6350) );
NAND2_X1 MEM_stage_inst_dmem_U6479 ( .A1(MEM_stage_inst_dmem_ram_2731), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n6351) );
NAND2_X1 MEM_stage_inst_dmem_U6478 ( .A1(MEM_stage_inst_dmem_n6349), .A2(MEM_stage_inst_dmem_n6348), .ZN(MEM_stage_inst_dmem_n6365) );
NOR2_X1 MEM_stage_inst_dmem_U6477 ( .A1(MEM_stage_inst_dmem_n6347), .A2(MEM_stage_inst_dmem_n6346), .ZN(MEM_stage_inst_dmem_n6348) );
NAND2_X1 MEM_stage_inst_dmem_U6476 ( .A1(MEM_stage_inst_dmem_n6345), .A2(MEM_stage_inst_dmem_n6344), .ZN(MEM_stage_inst_dmem_n6346) );
NAND2_X1 MEM_stage_inst_dmem_U6475 ( .A1(MEM_stage_inst_dmem_ram_2747), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n6344) );
NAND2_X1 MEM_stage_inst_dmem_U6474 ( .A1(MEM_stage_inst_dmem_ram_2155), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n6345) );
NAND2_X1 MEM_stage_inst_dmem_U6473 ( .A1(MEM_stage_inst_dmem_n6343), .A2(MEM_stage_inst_dmem_n6342), .ZN(MEM_stage_inst_dmem_n6347) );
NAND2_X1 MEM_stage_inst_dmem_U6472 ( .A1(MEM_stage_inst_dmem_ram_2379), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n6342) );
NAND2_X1 MEM_stage_inst_dmem_U6471 ( .A1(MEM_stage_inst_dmem_ram_2539), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n6343) );
NOR2_X1 MEM_stage_inst_dmem_U6470 ( .A1(MEM_stage_inst_dmem_n6341), .A2(MEM_stage_inst_dmem_n6340), .ZN(MEM_stage_inst_dmem_n6349) );
NAND2_X1 MEM_stage_inst_dmem_U6469 ( .A1(MEM_stage_inst_dmem_n6339), .A2(MEM_stage_inst_dmem_n6338), .ZN(MEM_stage_inst_dmem_n6340) );
NAND2_X1 MEM_stage_inst_dmem_U6468 ( .A1(MEM_stage_inst_dmem_ram_3035), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n6338) );
NAND2_X1 MEM_stage_inst_dmem_U6467 ( .A1(MEM_stage_inst_dmem_ram_2395), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n6339) );
NAND2_X1 MEM_stage_inst_dmem_U6466 ( .A1(MEM_stage_inst_dmem_n6337), .A2(MEM_stage_inst_dmem_n6336), .ZN(MEM_stage_inst_dmem_n6341) );
NAND2_X1 MEM_stage_inst_dmem_U6465 ( .A1(MEM_stage_inst_dmem_ram_2955), .A2(MEM_stage_inst_dmem_n8193), .ZN(MEM_stage_inst_dmem_n6336) );
NAND2_X1 MEM_stage_inst_dmem_U6464 ( .A1(MEM_stage_inst_dmem_ram_2795), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n6337) );
NOR2_X1 MEM_stage_inst_dmem_U6463 ( .A1(MEM_stage_inst_dmem_n6335), .A2(MEM_stage_inst_dmem_n8152), .ZN(MEM_stage_inst_dmem_n6464) );
NOR2_X1 MEM_stage_inst_dmem_U6462 ( .A1(MEM_stage_inst_dmem_n6334), .A2(MEM_stage_inst_dmem_n6333), .ZN(MEM_stage_inst_dmem_n6335) );
NAND2_X1 MEM_stage_inst_dmem_U6461 ( .A1(MEM_stage_inst_dmem_n6332), .A2(MEM_stage_inst_dmem_n6331), .ZN(MEM_stage_inst_dmem_n6333) );
NOR2_X1 MEM_stage_inst_dmem_U6460 ( .A1(MEM_stage_inst_dmem_n6330), .A2(MEM_stage_inst_dmem_n6329), .ZN(MEM_stage_inst_dmem_n6331) );
NAND2_X1 MEM_stage_inst_dmem_U6459 ( .A1(MEM_stage_inst_dmem_n6328), .A2(MEM_stage_inst_dmem_n6327), .ZN(MEM_stage_inst_dmem_n6329) );
NOR2_X1 MEM_stage_inst_dmem_U6458 ( .A1(MEM_stage_inst_dmem_n6326), .A2(MEM_stage_inst_dmem_n6325), .ZN(MEM_stage_inst_dmem_n6327) );
NAND2_X1 MEM_stage_inst_dmem_U6457 ( .A1(MEM_stage_inst_dmem_n6324), .A2(MEM_stage_inst_dmem_n6323), .ZN(MEM_stage_inst_dmem_n6325) );
NAND2_X1 MEM_stage_inst_dmem_U6456 ( .A1(MEM_stage_inst_dmem_ram_1243), .A2(MEM_stage_inst_dmem_n8206), .ZN(MEM_stage_inst_dmem_n6323) );
NAND2_X1 MEM_stage_inst_dmem_U6455 ( .A1(MEM_stage_inst_dmem_ram_1627), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n6324) );
NAND2_X1 MEM_stage_inst_dmem_U6454 ( .A1(MEM_stage_inst_dmem_n6322), .A2(MEM_stage_inst_dmem_n6321), .ZN(MEM_stage_inst_dmem_n6326) );
NAND2_X1 MEM_stage_inst_dmem_U6453 ( .A1(MEM_stage_inst_dmem_ram_1259), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n6321) );
NAND2_X1 MEM_stage_inst_dmem_U6452 ( .A1(MEM_stage_inst_dmem_ram_1499), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n6322) );
NOR2_X1 MEM_stage_inst_dmem_U6451 ( .A1(MEM_stage_inst_dmem_n6320), .A2(MEM_stage_inst_dmem_n6319), .ZN(MEM_stage_inst_dmem_n6328) );
NAND2_X1 MEM_stage_inst_dmem_U6450 ( .A1(MEM_stage_inst_dmem_n6318), .A2(MEM_stage_inst_dmem_n6317), .ZN(MEM_stage_inst_dmem_n6319) );
NAND2_X1 MEM_stage_inst_dmem_U6449 ( .A1(MEM_stage_inst_dmem_ram_1899), .A2(MEM_stage_inst_dmem_n7923), .ZN(MEM_stage_inst_dmem_n6317) );
NAND2_X1 MEM_stage_inst_dmem_U6448 ( .A1(MEM_stage_inst_dmem_ram_1131), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n6318) );
NAND2_X1 MEM_stage_inst_dmem_U6447 ( .A1(MEM_stage_inst_dmem_n6316), .A2(MEM_stage_inst_dmem_n6315), .ZN(MEM_stage_inst_dmem_n6320) );
NAND2_X1 MEM_stage_inst_dmem_U6446 ( .A1(MEM_stage_inst_dmem_ram_1883), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n6315) );
NAND2_X1 MEM_stage_inst_dmem_U6445 ( .A1(MEM_stage_inst_dmem_ram_1947), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n6316) );
NAND2_X1 MEM_stage_inst_dmem_U6444 ( .A1(MEM_stage_inst_dmem_n6314), .A2(MEM_stage_inst_dmem_n6313), .ZN(MEM_stage_inst_dmem_n6330) );
NOR2_X1 MEM_stage_inst_dmem_U6443 ( .A1(MEM_stage_inst_dmem_n6312), .A2(MEM_stage_inst_dmem_n6311), .ZN(MEM_stage_inst_dmem_n6313) );
NAND2_X1 MEM_stage_inst_dmem_U6442 ( .A1(MEM_stage_inst_dmem_n6310), .A2(MEM_stage_inst_dmem_n6309), .ZN(MEM_stage_inst_dmem_n6311) );
NAND2_X1 MEM_stage_inst_dmem_U6441 ( .A1(MEM_stage_inst_dmem_ram_1515), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n6309) );
NAND2_X1 MEM_stage_inst_dmem_U6440 ( .A1(MEM_stage_inst_dmem_ram_1371), .A2(MEM_stage_inst_dmem_n3216), .ZN(MEM_stage_inst_dmem_n6310) );
NAND2_X1 MEM_stage_inst_dmem_U6439 ( .A1(MEM_stage_inst_dmem_n6308), .A2(MEM_stage_inst_dmem_n6307), .ZN(MEM_stage_inst_dmem_n6312) );
NAND2_X1 MEM_stage_inst_dmem_U6438 ( .A1(MEM_stage_inst_dmem_ram_1755), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n6307) );
NAND2_X1 MEM_stage_inst_dmem_U6437 ( .A1(MEM_stage_inst_dmem_ram_1611), .A2(MEM_stage_inst_dmem_n7973), .ZN(MEM_stage_inst_dmem_n6308) );
NOR2_X1 MEM_stage_inst_dmem_U6436 ( .A1(MEM_stage_inst_dmem_n6306), .A2(MEM_stage_inst_dmem_n6305), .ZN(MEM_stage_inst_dmem_n6314) );
NAND2_X1 MEM_stage_inst_dmem_U6435 ( .A1(MEM_stage_inst_dmem_n6304), .A2(MEM_stage_inst_dmem_n6303), .ZN(MEM_stage_inst_dmem_n6305) );
NAND2_X1 MEM_stage_inst_dmem_U6434 ( .A1(MEM_stage_inst_dmem_ram_1163), .A2(MEM_stage_inst_dmem_n8174), .ZN(MEM_stage_inst_dmem_n6303) );
NAND2_X1 MEM_stage_inst_dmem_U6433 ( .A1(MEM_stage_inst_dmem_ram_1835), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n6304) );
NAND2_X1 MEM_stage_inst_dmem_U6432 ( .A1(MEM_stage_inst_dmem_n6302), .A2(MEM_stage_inst_dmem_n6301), .ZN(MEM_stage_inst_dmem_n6306) );
NAND2_X1 MEM_stage_inst_dmem_U6431 ( .A1(MEM_stage_inst_dmem_ram_1355), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n6301) );
NAND2_X1 MEM_stage_inst_dmem_U6430 ( .A1(MEM_stage_inst_dmem_ram_1179), .A2(MEM_stage_inst_dmem_n7903), .ZN(MEM_stage_inst_dmem_n6302) );
NOR2_X1 MEM_stage_inst_dmem_U6429 ( .A1(MEM_stage_inst_dmem_n6300), .A2(MEM_stage_inst_dmem_n6299), .ZN(MEM_stage_inst_dmem_n6332) );
NAND2_X1 MEM_stage_inst_dmem_U6428 ( .A1(MEM_stage_inst_dmem_n6298), .A2(MEM_stage_inst_dmem_n6297), .ZN(MEM_stage_inst_dmem_n6299) );
NOR2_X1 MEM_stage_inst_dmem_U6427 ( .A1(MEM_stage_inst_dmem_n6296), .A2(MEM_stage_inst_dmem_n6295), .ZN(MEM_stage_inst_dmem_n6297) );
NAND2_X1 MEM_stage_inst_dmem_U6426 ( .A1(MEM_stage_inst_dmem_n6294), .A2(MEM_stage_inst_dmem_n6293), .ZN(MEM_stage_inst_dmem_n6295) );
NAND2_X1 MEM_stage_inst_dmem_U6425 ( .A1(MEM_stage_inst_dmem_ram_1915), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n6293) );
NAND2_X1 MEM_stage_inst_dmem_U6424 ( .A1(MEM_stage_inst_dmem_ram_1291), .A2(MEM_stage_inst_dmem_n7898), .ZN(MEM_stage_inst_dmem_n6294) );
NAND2_X1 MEM_stage_inst_dmem_U6423 ( .A1(MEM_stage_inst_dmem_n6292), .A2(MEM_stage_inst_dmem_n6291), .ZN(MEM_stage_inst_dmem_n6296) );
NAND2_X1 MEM_stage_inst_dmem_U6422 ( .A1(MEM_stage_inst_dmem_ram_1803), .A2(MEM_stage_inst_dmem_n7992), .ZN(MEM_stage_inst_dmem_n6291) );
NAND2_X1 MEM_stage_inst_dmem_U6421 ( .A1(MEM_stage_inst_dmem_ram_1787), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n6292) );
NOR2_X1 MEM_stage_inst_dmem_U6420 ( .A1(MEM_stage_inst_dmem_n6290), .A2(MEM_stage_inst_dmem_n6289), .ZN(MEM_stage_inst_dmem_n6298) );
NAND2_X1 MEM_stage_inst_dmem_U6419 ( .A1(MEM_stage_inst_dmem_n6288), .A2(MEM_stage_inst_dmem_n6287), .ZN(MEM_stage_inst_dmem_n6289) );
NAND2_X1 MEM_stage_inst_dmem_U6418 ( .A1(MEM_stage_inst_dmem_ram_1931), .A2(MEM_stage_inst_dmem_n8193), .ZN(MEM_stage_inst_dmem_n6287) );
NAND2_X1 MEM_stage_inst_dmem_U6417 ( .A1(MEM_stage_inst_dmem_ram_1035), .A2(MEM_stage_inst_dmem_n7953), .ZN(MEM_stage_inst_dmem_n6288) );
NAND2_X1 MEM_stage_inst_dmem_U6416 ( .A1(MEM_stage_inst_dmem_n6286), .A2(MEM_stage_inst_dmem_n6285), .ZN(MEM_stage_inst_dmem_n6290) );
NAND2_X1 MEM_stage_inst_dmem_U6415 ( .A1(MEM_stage_inst_dmem_ram_1867), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n6285) );
NAND2_X1 MEM_stage_inst_dmem_U6414 ( .A1(MEM_stage_inst_dmem_ram_1739), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n6286) );
NAND2_X1 MEM_stage_inst_dmem_U6413 ( .A1(MEM_stage_inst_dmem_n6284), .A2(MEM_stage_inst_dmem_n6283), .ZN(MEM_stage_inst_dmem_n6300) );
NOR2_X1 MEM_stage_inst_dmem_U6412 ( .A1(MEM_stage_inst_dmem_n6282), .A2(MEM_stage_inst_dmem_n6281), .ZN(MEM_stage_inst_dmem_n6283) );
NAND2_X1 MEM_stage_inst_dmem_U6411 ( .A1(MEM_stage_inst_dmem_n6280), .A2(MEM_stage_inst_dmem_n6279), .ZN(MEM_stage_inst_dmem_n6281) );
NAND2_X1 MEM_stage_inst_dmem_U6410 ( .A1(MEM_stage_inst_dmem_ram_1451), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n6279) );
NAND2_X1 MEM_stage_inst_dmem_U6409 ( .A1(MEM_stage_inst_dmem_ram_1963), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n6280) );
NAND2_X1 MEM_stage_inst_dmem_U6408 ( .A1(MEM_stage_inst_dmem_n6278), .A2(MEM_stage_inst_dmem_n6277), .ZN(MEM_stage_inst_dmem_n6282) );
NAND2_X1 MEM_stage_inst_dmem_U6407 ( .A1(MEM_stage_inst_dmem_ram_1227), .A2(MEM_stage_inst_dmem_n8256), .ZN(MEM_stage_inst_dmem_n6277) );
NAND2_X1 MEM_stage_inst_dmem_U6406 ( .A1(MEM_stage_inst_dmem_ram_1595), .A2(MEM_stage_inst_dmem_n8169), .ZN(MEM_stage_inst_dmem_n6278) );
NOR2_X1 MEM_stage_inst_dmem_U6405 ( .A1(MEM_stage_inst_dmem_n6276), .A2(MEM_stage_inst_dmem_n6275), .ZN(MEM_stage_inst_dmem_n6284) );
NAND2_X1 MEM_stage_inst_dmem_U6404 ( .A1(MEM_stage_inst_dmem_n6274), .A2(MEM_stage_inst_dmem_n6273), .ZN(MEM_stage_inst_dmem_n6275) );
NAND2_X1 MEM_stage_inst_dmem_U6403 ( .A1(MEM_stage_inst_dmem_ram_1339), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n6273) );
NAND2_X1 MEM_stage_inst_dmem_U6402 ( .A1(MEM_stage_inst_dmem_ram_1979), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n6274) );
NAND2_X1 MEM_stage_inst_dmem_U6401 ( .A1(MEM_stage_inst_dmem_n6272), .A2(MEM_stage_inst_dmem_n6271), .ZN(MEM_stage_inst_dmem_n6276) );
NAND2_X1 MEM_stage_inst_dmem_U6400 ( .A1(MEM_stage_inst_dmem_ram_1467), .A2(MEM_stage_inst_dmem_n7888), .ZN(MEM_stage_inst_dmem_n6271) );
NAND2_X1 MEM_stage_inst_dmem_U6399 ( .A1(MEM_stage_inst_dmem_ram_1851), .A2(MEM_stage_inst_dmem_n46), .ZN(MEM_stage_inst_dmem_n6272) );
NAND2_X1 MEM_stage_inst_dmem_U6398 ( .A1(MEM_stage_inst_dmem_n6270), .A2(MEM_stage_inst_dmem_n6269), .ZN(MEM_stage_inst_dmem_n6334) );
NOR2_X1 MEM_stage_inst_dmem_U6397 ( .A1(MEM_stage_inst_dmem_n6268), .A2(MEM_stage_inst_dmem_n6267), .ZN(MEM_stage_inst_dmem_n6269) );
NAND2_X1 MEM_stage_inst_dmem_U6396 ( .A1(MEM_stage_inst_dmem_n6266), .A2(MEM_stage_inst_dmem_n6265), .ZN(MEM_stage_inst_dmem_n6267) );
NOR2_X1 MEM_stage_inst_dmem_U6395 ( .A1(MEM_stage_inst_dmem_n6264), .A2(MEM_stage_inst_dmem_n6263), .ZN(MEM_stage_inst_dmem_n6265) );
NAND2_X1 MEM_stage_inst_dmem_U6394 ( .A1(MEM_stage_inst_dmem_n6262), .A2(MEM_stage_inst_dmem_n6261), .ZN(MEM_stage_inst_dmem_n6263) );
NAND2_X1 MEM_stage_inst_dmem_U6393 ( .A1(MEM_stage_inst_dmem_ram_1707), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n6261) );
NAND2_X1 MEM_stage_inst_dmem_U6392 ( .A1(MEM_stage_inst_dmem_ram_1723), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n6262) );
NAND2_X1 MEM_stage_inst_dmem_U6391 ( .A1(MEM_stage_inst_dmem_n6260), .A2(MEM_stage_inst_dmem_n6259), .ZN(MEM_stage_inst_dmem_n6264) );
NAND2_X1 MEM_stage_inst_dmem_U6390 ( .A1(MEM_stage_inst_dmem_ram_1435), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n6259) );
NAND2_X1 MEM_stage_inst_dmem_U6389 ( .A1(MEM_stage_inst_dmem_ram_2043), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n6260) );
NOR2_X1 MEM_stage_inst_dmem_U6388 ( .A1(MEM_stage_inst_dmem_n6258), .A2(MEM_stage_inst_dmem_n6257), .ZN(MEM_stage_inst_dmem_n6266) );
NAND2_X1 MEM_stage_inst_dmem_U6387 ( .A1(MEM_stage_inst_dmem_n6256), .A2(MEM_stage_inst_dmem_n6255), .ZN(MEM_stage_inst_dmem_n6257) );
NAND2_X1 MEM_stage_inst_dmem_U6386 ( .A1(MEM_stage_inst_dmem_ram_2011), .A2(MEM_stage_inst_dmem_n7895), .ZN(MEM_stage_inst_dmem_n6255) );
NAND2_X1 MEM_stage_inst_dmem_U6385 ( .A1(MEM_stage_inst_dmem_ram_1771), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n6256) );
NAND2_X1 MEM_stage_inst_dmem_U6384 ( .A1(MEM_stage_inst_dmem_n6254), .A2(MEM_stage_inst_dmem_n6253), .ZN(MEM_stage_inst_dmem_n6258) );
NAND2_X1 MEM_stage_inst_dmem_U6383 ( .A1(MEM_stage_inst_dmem_ram_1099), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n6253) );
NAND2_X1 MEM_stage_inst_dmem_U6382 ( .A1(MEM_stage_inst_dmem_ram_1995), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n6254) );
NAND2_X1 MEM_stage_inst_dmem_U6381 ( .A1(MEM_stage_inst_dmem_n6252), .A2(MEM_stage_inst_dmem_n6251), .ZN(MEM_stage_inst_dmem_n6268) );
NOR2_X1 MEM_stage_inst_dmem_U6380 ( .A1(MEM_stage_inst_dmem_n6250), .A2(MEM_stage_inst_dmem_n6249), .ZN(MEM_stage_inst_dmem_n6251) );
NAND2_X1 MEM_stage_inst_dmem_U6379 ( .A1(MEM_stage_inst_dmem_n6248), .A2(MEM_stage_inst_dmem_n6247), .ZN(MEM_stage_inst_dmem_n6249) );
NAND2_X1 MEM_stage_inst_dmem_U6378 ( .A1(MEM_stage_inst_dmem_ram_1531), .A2(MEM_stage_inst_dmem_n64), .ZN(MEM_stage_inst_dmem_n6247) );
NAND2_X1 MEM_stage_inst_dmem_U6377 ( .A1(MEM_stage_inst_dmem_ram_1691), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n6248) );
NAND2_X1 MEM_stage_inst_dmem_U6376 ( .A1(MEM_stage_inst_dmem_n6246), .A2(MEM_stage_inst_dmem_n6245), .ZN(MEM_stage_inst_dmem_n6250) );
NAND2_X1 MEM_stage_inst_dmem_U6375 ( .A1(MEM_stage_inst_dmem_ram_1051), .A2(MEM_stage_inst_dmem_n7887), .ZN(MEM_stage_inst_dmem_n6245) );
NAND2_X1 MEM_stage_inst_dmem_U6374 ( .A1(MEM_stage_inst_dmem_ram_1643), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n6246) );
NOR2_X1 MEM_stage_inst_dmem_U6373 ( .A1(MEM_stage_inst_dmem_n6244), .A2(MEM_stage_inst_dmem_n6243), .ZN(MEM_stage_inst_dmem_n6252) );
NAND2_X1 MEM_stage_inst_dmem_U6372 ( .A1(MEM_stage_inst_dmem_n6242), .A2(MEM_stage_inst_dmem_n6241), .ZN(MEM_stage_inst_dmem_n6243) );
NAND2_X1 MEM_stage_inst_dmem_U6371 ( .A1(MEM_stage_inst_dmem_ram_1387), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n6241) );
NAND2_X1 MEM_stage_inst_dmem_U6370 ( .A1(MEM_stage_inst_dmem_ram_1275), .A2(MEM_stage_inst_dmem_n39), .ZN(MEM_stage_inst_dmem_n6242) );
NAND2_X1 MEM_stage_inst_dmem_U6369 ( .A1(MEM_stage_inst_dmem_n6240), .A2(MEM_stage_inst_dmem_n6239), .ZN(MEM_stage_inst_dmem_n6244) );
NAND2_X1 MEM_stage_inst_dmem_U6368 ( .A1(MEM_stage_inst_dmem_ram_1579), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n6239) );
NAND2_X1 MEM_stage_inst_dmem_U6367 ( .A1(MEM_stage_inst_dmem_ram_1419), .A2(MEM_stage_inst_dmem_n7930), .ZN(MEM_stage_inst_dmem_n6240) );
NOR2_X1 MEM_stage_inst_dmem_U6366 ( .A1(MEM_stage_inst_dmem_n6238), .A2(MEM_stage_inst_dmem_n6237), .ZN(MEM_stage_inst_dmem_n6270) );
NAND2_X1 MEM_stage_inst_dmem_U6365 ( .A1(MEM_stage_inst_dmem_n6236), .A2(MEM_stage_inst_dmem_n6235), .ZN(MEM_stage_inst_dmem_n6237) );
NOR2_X1 MEM_stage_inst_dmem_U6364 ( .A1(MEM_stage_inst_dmem_n6234), .A2(MEM_stage_inst_dmem_n6233), .ZN(MEM_stage_inst_dmem_n6235) );
NAND2_X1 MEM_stage_inst_dmem_U6363 ( .A1(MEM_stage_inst_dmem_n6232), .A2(MEM_stage_inst_dmem_n6231), .ZN(MEM_stage_inst_dmem_n6233) );
NAND2_X1 MEM_stage_inst_dmem_U6362 ( .A1(MEM_stage_inst_dmem_ram_1675), .A2(MEM_stage_inst_dmem_n7960), .ZN(MEM_stage_inst_dmem_n6231) );
NAND2_X1 MEM_stage_inst_dmem_U6361 ( .A1(MEM_stage_inst_dmem_ram_1323), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n6232) );
NAND2_X1 MEM_stage_inst_dmem_U6360 ( .A1(MEM_stage_inst_dmem_n6230), .A2(MEM_stage_inst_dmem_n6229), .ZN(MEM_stage_inst_dmem_n6234) );
NAND2_X1 MEM_stage_inst_dmem_U6359 ( .A1(MEM_stage_inst_dmem_ram_1083), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n6229) );
NAND2_X1 MEM_stage_inst_dmem_U6358 ( .A1(MEM_stage_inst_dmem_ram_1547), .A2(MEM_stage_inst_dmem_n8225), .ZN(MEM_stage_inst_dmem_n6230) );
NOR2_X1 MEM_stage_inst_dmem_U6357 ( .A1(MEM_stage_inst_dmem_n6228), .A2(MEM_stage_inst_dmem_n6227), .ZN(MEM_stage_inst_dmem_n6236) );
NAND2_X1 MEM_stage_inst_dmem_U6356 ( .A1(MEM_stage_inst_dmem_n6226), .A2(MEM_stage_inst_dmem_n6225), .ZN(MEM_stage_inst_dmem_n6227) );
NAND2_X1 MEM_stage_inst_dmem_U6355 ( .A1(MEM_stage_inst_dmem_ram_1147), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n6225) );
NAND2_X1 MEM_stage_inst_dmem_U6354 ( .A1(MEM_stage_inst_dmem_ram_1403), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n6226) );
NAND2_X1 MEM_stage_inst_dmem_U6353 ( .A1(MEM_stage_inst_dmem_n6224), .A2(MEM_stage_inst_dmem_n6223), .ZN(MEM_stage_inst_dmem_n6228) );
NAND2_X1 MEM_stage_inst_dmem_U6352 ( .A1(MEM_stage_inst_dmem_ram_1211), .A2(MEM_stage_inst_dmem_n7937), .ZN(MEM_stage_inst_dmem_n6223) );
NAND2_X1 MEM_stage_inst_dmem_U6351 ( .A1(MEM_stage_inst_dmem_ram_1819), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n6224) );
NAND2_X1 MEM_stage_inst_dmem_U6350 ( .A1(MEM_stage_inst_dmem_n6222), .A2(MEM_stage_inst_dmem_n6221), .ZN(MEM_stage_inst_dmem_n6238) );
NOR2_X1 MEM_stage_inst_dmem_U6349 ( .A1(MEM_stage_inst_dmem_n6220), .A2(MEM_stage_inst_dmem_n6219), .ZN(MEM_stage_inst_dmem_n6221) );
NAND2_X1 MEM_stage_inst_dmem_U6348 ( .A1(MEM_stage_inst_dmem_n6218), .A2(MEM_stage_inst_dmem_n6217), .ZN(MEM_stage_inst_dmem_n6219) );
NAND2_X1 MEM_stage_inst_dmem_U6347 ( .A1(MEM_stage_inst_dmem_ram_1483), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n6217) );
NAND2_X1 MEM_stage_inst_dmem_U6346 ( .A1(MEM_stage_inst_dmem_ram_1195), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n6218) );
NAND2_X1 MEM_stage_inst_dmem_U6345 ( .A1(MEM_stage_inst_dmem_n6216), .A2(MEM_stage_inst_dmem_n6215), .ZN(MEM_stage_inst_dmem_n6220) );
NAND2_X1 MEM_stage_inst_dmem_U6344 ( .A1(MEM_stage_inst_dmem_ram_2027), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n6215) );
NAND2_X1 MEM_stage_inst_dmem_U6343 ( .A1(MEM_stage_inst_dmem_ram_1115), .A2(MEM_stage_inst_dmem_n7938), .ZN(MEM_stage_inst_dmem_n6216) );
NOR2_X1 MEM_stage_inst_dmem_U6342 ( .A1(MEM_stage_inst_dmem_n6214), .A2(MEM_stage_inst_dmem_n6213), .ZN(MEM_stage_inst_dmem_n6222) );
NAND2_X1 MEM_stage_inst_dmem_U6341 ( .A1(MEM_stage_inst_dmem_n6212), .A2(MEM_stage_inst_dmem_n6211), .ZN(MEM_stage_inst_dmem_n6213) );
NAND2_X1 MEM_stage_inst_dmem_U6340 ( .A1(MEM_stage_inst_dmem_ram_1067), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n6211) );
NAND2_X1 MEM_stage_inst_dmem_U6339 ( .A1(MEM_stage_inst_dmem_ram_1563), .A2(MEM_stage_inst_dmem_n7884), .ZN(MEM_stage_inst_dmem_n6212) );
NAND2_X1 MEM_stage_inst_dmem_U6338 ( .A1(MEM_stage_inst_dmem_n6210), .A2(MEM_stage_inst_dmem_n6209), .ZN(MEM_stage_inst_dmem_n6214) );
NAND2_X1 MEM_stage_inst_dmem_U6337 ( .A1(MEM_stage_inst_dmem_ram_1307), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n6209) );
NAND2_X1 MEM_stage_inst_dmem_U6336 ( .A1(MEM_stage_inst_dmem_ram_1659), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n6210) );
NOR2_X1 MEM_stage_inst_dmem_U6335 ( .A1(MEM_stage_inst_dmem_n6208), .A2(MEM_stage_inst_dmem_n6207), .ZN(MEM_stage_inst_dmem_n6466) );
NOR2_X1 MEM_stage_inst_dmem_U6334 ( .A1(MEM_stage_inst_dmem_n6206), .A2(MEM_stage_inst_dmem_n8551), .ZN(MEM_stage_inst_dmem_n6207) );
NOR2_X1 MEM_stage_inst_dmem_U6333 ( .A1(MEM_stage_inst_dmem_n6205), .A2(MEM_stage_inst_dmem_n6204), .ZN(MEM_stage_inst_dmem_n6206) );
NAND2_X1 MEM_stage_inst_dmem_U6332 ( .A1(MEM_stage_inst_dmem_n6203), .A2(MEM_stage_inst_dmem_n6202), .ZN(MEM_stage_inst_dmem_n6204) );
NOR2_X1 MEM_stage_inst_dmem_U6331 ( .A1(MEM_stage_inst_dmem_n6201), .A2(MEM_stage_inst_dmem_n6200), .ZN(MEM_stage_inst_dmem_n6202) );
NAND2_X1 MEM_stage_inst_dmem_U6330 ( .A1(MEM_stage_inst_dmem_n6199), .A2(MEM_stage_inst_dmem_n6198), .ZN(MEM_stage_inst_dmem_n6200) );
NOR2_X1 MEM_stage_inst_dmem_U6329 ( .A1(MEM_stage_inst_dmem_n6197), .A2(MEM_stage_inst_dmem_n6196), .ZN(MEM_stage_inst_dmem_n6198) );
NAND2_X1 MEM_stage_inst_dmem_U6328 ( .A1(MEM_stage_inst_dmem_n6195), .A2(MEM_stage_inst_dmem_n6194), .ZN(MEM_stage_inst_dmem_n6196) );
NAND2_X1 MEM_stage_inst_dmem_U6327 ( .A1(MEM_stage_inst_dmem_ram_139), .A2(MEM_stage_inst_dmem_n8174), .ZN(MEM_stage_inst_dmem_n6194) );
NAND2_X1 MEM_stage_inst_dmem_U6326 ( .A1(MEM_stage_inst_dmem_ram_283), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n6195) );
NAND2_X1 MEM_stage_inst_dmem_U6325 ( .A1(MEM_stage_inst_dmem_n6193), .A2(MEM_stage_inst_dmem_n6192), .ZN(MEM_stage_inst_dmem_n6197) );
NAND2_X1 MEM_stage_inst_dmem_U6324 ( .A1(MEM_stage_inst_dmem_ram_1003), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n6192) );
NAND2_X1 MEM_stage_inst_dmem_U6323 ( .A1(MEM_stage_inst_dmem_ram_299), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n6193) );
NOR2_X1 MEM_stage_inst_dmem_U6322 ( .A1(MEM_stage_inst_dmem_n6191), .A2(MEM_stage_inst_dmem_n6190), .ZN(MEM_stage_inst_dmem_n6199) );
NAND2_X1 MEM_stage_inst_dmem_U6321 ( .A1(MEM_stage_inst_dmem_n6189), .A2(MEM_stage_inst_dmem_n6188), .ZN(MEM_stage_inst_dmem_n6190) );
NAND2_X1 MEM_stage_inst_dmem_U6320 ( .A1(MEM_stage_inst_dmem_ram_187), .A2(MEM_stage_inst_dmem_n7937), .ZN(MEM_stage_inst_dmem_n6188) );
NAND2_X1 MEM_stage_inst_dmem_U6319 ( .A1(MEM_stage_inst_dmem_ram_379), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n6189) );
NAND2_X1 MEM_stage_inst_dmem_U6318 ( .A1(MEM_stage_inst_dmem_n6187), .A2(MEM_stage_inst_dmem_n6186), .ZN(MEM_stage_inst_dmem_n6191) );
NAND2_X1 MEM_stage_inst_dmem_U6317 ( .A1(MEM_stage_inst_dmem_ram_955), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n6186) );
NAND2_X1 MEM_stage_inst_dmem_U6316 ( .A1(MEM_stage_inst_dmem_ram_587), .A2(MEM_stage_inst_dmem_n7973), .ZN(MEM_stage_inst_dmem_n6187) );
NAND2_X1 MEM_stage_inst_dmem_U6315 ( .A1(MEM_stage_inst_dmem_n6185), .A2(MEM_stage_inst_dmem_n6184), .ZN(MEM_stage_inst_dmem_n6201) );
NOR2_X1 MEM_stage_inst_dmem_U6314 ( .A1(MEM_stage_inst_dmem_n6183), .A2(MEM_stage_inst_dmem_n6182), .ZN(MEM_stage_inst_dmem_n6184) );
NAND2_X1 MEM_stage_inst_dmem_U6313 ( .A1(MEM_stage_inst_dmem_n6181), .A2(MEM_stage_inst_dmem_n6180), .ZN(MEM_stage_inst_dmem_n6182) );
NAND2_X1 MEM_stage_inst_dmem_U6312 ( .A1(MEM_stage_inst_dmem_ram_27), .A2(MEM_stage_inst_dmem_n7887), .ZN(MEM_stage_inst_dmem_n6180) );
NAND2_X1 MEM_stage_inst_dmem_U6311 ( .A1(MEM_stage_inst_dmem_ram_347), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n6181) );
NAND2_X1 MEM_stage_inst_dmem_U6310 ( .A1(MEM_stage_inst_dmem_n6179), .A2(MEM_stage_inst_dmem_n6178), .ZN(MEM_stage_inst_dmem_n6183) );
NAND2_X1 MEM_stage_inst_dmem_U6309 ( .A1(MEM_stage_inst_dmem_ram_363), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n6178) );
NAND2_X1 MEM_stage_inst_dmem_U6308 ( .A1(MEM_stage_inst_dmem_ram_59), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n6179) );
NOR2_X1 MEM_stage_inst_dmem_U6307 ( .A1(MEM_stage_inst_dmem_n6177), .A2(MEM_stage_inst_dmem_n6176), .ZN(MEM_stage_inst_dmem_n6185) );
NAND2_X1 MEM_stage_inst_dmem_U6306 ( .A1(MEM_stage_inst_dmem_n6175), .A2(MEM_stage_inst_dmem_n6174), .ZN(MEM_stage_inst_dmem_n6176) );
NAND2_X1 MEM_stage_inst_dmem_U6305 ( .A1(MEM_stage_inst_dmem_ram_251), .A2(MEM_stage_inst_dmem_n39), .ZN(MEM_stage_inst_dmem_n6174) );
NAND2_X1 MEM_stage_inst_dmem_U6304 ( .A1(MEM_stage_inst_dmem_ram_603), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n6175) );
NAND2_X1 MEM_stage_inst_dmem_U6303 ( .A1(MEM_stage_inst_dmem_n6173), .A2(MEM_stage_inst_dmem_n6172), .ZN(MEM_stage_inst_dmem_n6177) );
NAND2_X1 MEM_stage_inst_dmem_U6302 ( .A1(MEM_stage_inst_dmem_ram_43), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n6172) );
NAND2_X1 MEM_stage_inst_dmem_U6301 ( .A1(MEM_stage_inst_dmem_ram_11), .A2(MEM_stage_inst_dmem_n7953), .ZN(MEM_stage_inst_dmem_n6173) );
NOR2_X1 MEM_stage_inst_dmem_U6300 ( .A1(MEM_stage_inst_dmem_n6171), .A2(MEM_stage_inst_dmem_n6170), .ZN(MEM_stage_inst_dmem_n6203) );
NAND2_X1 MEM_stage_inst_dmem_U6299 ( .A1(MEM_stage_inst_dmem_n6169), .A2(MEM_stage_inst_dmem_n6168), .ZN(MEM_stage_inst_dmem_n6170) );
NOR2_X1 MEM_stage_inst_dmem_U6298 ( .A1(MEM_stage_inst_dmem_n6167), .A2(MEM_stage_inst_dmem_n6166), .ZN(MEM_stage_inst_dmem_n6168) );
NAND2_X1 MEM_stage_inst_dmem_U6297 ( .A1(MEM_stage_inst_dmem_n6165), .A2(MEM_stage_inst_dmem_n6164), .ZN(MEM_stage_inst_dmem_n6166) );
NAND2_X1 MEM_stage_inst_dmem_U6296 ( .A1(MEM_stage_inst_dmem_ram_555), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n6164) );
NAND2_X1 MEM_stage_inst_dmem_U6295 ( .A1(MEM_stage_inst_dmem_ram_219), .A2(MEM_stage_inst_dmem_n8206), .ZN(MEM_stage_inst_dmem_n6165) );
NAND2_X1 MEM_stage_inst_dmem_U6294 ( .A1(MEM_stage_inst_dmem_n6163), .A2(MEM_stage_inst_dmem_n6162), .ZN(MEM_stage_inst_dmem_n6167) );
NAND2_X1 MEM_stage_inst_dmem_U6293 ( .A1(MEM_stage_inst_dmem_ram_75), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n6162) );
NAND2_X1 MEM_stage_inst_dmem_U6292 ( .A1(MEM_stage_inst_dmem_ram_827), .A2(MEM_stage_inst_dmem_n46), .ZN(MEM_stage_inst_dmem_n6163) );
NOR2_X1 MEM_stage_inst_dmem_U6291 ( .A1(MEM_stage_inst_dmem_n6161), .A2(MEM_stage_inst_dmem_n6160), .ZN(MEM_stage_inst_dmem_n6169) );
NAND2_X1 MEM_stage_inst_dmem_U6290 ( .A1(MEM_stage_inst_dmem_n6159), .A2(MEM_stage_inst_dmem_n6158), .ZN(MEM_stage_inst_dmem_n6160) );
NAND2_X1 MEM_stage_inst_dmem_U6289 ( .A1(MEM_stage_inst_dmem_ram_859), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n6158) );
NAND2_X1 MEM_stage_inst_dmem_U6288 ( .A1(MEM_stage_inst_dmem_ram_635), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n6159) );
NAND2_X1 MEM_stage_inst_dmem_U6287 ( .A1(MEM_stage_inst_dmem_n6157), .A2(MEM_stage_inst_dmem_n6156), .ZN(MEM_stage_inst_dmem_n6161) );
NAND2_X1 MEM_stage_inst_dmem_U6286 ( .A1(MEM_stage_inst_dmem_ram_891), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n6156) );
NAND2_X1 MEM_stage_inst_dmem_U6285 ( .A1(MEM_stage_inst_dmem_ram_795), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n6157) );
NAND2_X1 MEM_stage_inst_dmem_U6284 ( .A1(MEM_stage_inst_dmem_n6155), .A2(MEM_stage_inst_dmem_n6154), .ZN(MEM_stage_inst_dmem_n6171) );
NOR2_X1 MEM_stage_inst_dmem_U6283 ( .A1(MEM_stage_inst_dmem_n6153), .A2(MEM_stage_inst_dmem_n6152), .ZN(MEM_stage_inst_dmem_n6154) );
NAND2_X1 MEM_stage_inst_dmem_U6282 ( .A1(MEM_stage_inst_dmem_n6151), .A2(MEM_stage_inst_dmem_n6150), .ZN(MEM_stage_inst_dmem_n6152) );
NAND2_X1 MEM_stage_inst_dmem_U6281 ( .A1(MEM_stage_inst_dmem_ram_123), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n6150) );
NAND2_X1 MEM_stage_inst_dmem_U6280 ( .A1(MEM_stage_inst_dmem_ram_459), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n6151) );
NAND2_X1 MEM_stage_inst_dmem_U6279 ( .A1(MEM_stage_inst_dmem_n6149), .A2(MEM_stage_inst_dmem_n6148), .ZN(MEM_stage_inst_dmem_n6153) );
NAND2_X1 MEM_stage_inst_dmem_U6278 ( .A1(MEM_stage_inst_dmem_ram_507), .A2(MEM_stage_inst_dmem_n64), .ZN(MEM_stage_inst_dmem_n6148) );
NAND2_X1 MEM_stage_inst_dmem_U6277 ( .A1(MEM_stage_inst_dmem_ram_267), .A2(MEM_stage_inst_dmem_n7898), .ZN(MEM_stage_inst_dmem_n6149) );
NOR2_X1 MEM_stage_inst_dmem_U6276 ( .A1(MEM_stage_inst_dmem_n6147), .A2(MEM_stage_inst_dmem_n6146), .ZN(MEM_stage_inst_dmem_n6155) );
NAND2_X1 MEM_stage_inst_dmem_U6275 ( .A1(MEM_stage_inst_dmem_n6145), .A2(MEM_stage_inst_dmem_n6144), .ZN(MEM_stage_inst_dmem_n6146) );
NAND2_X1 MEM_stage_inst_dmem_U6274 ( .A1(MEM_stage_inst_dmem_ram_875), .A2(MEM_stage_inst_dmem_n7923), .ZN(MEM_stage_inst_dmem_n6144) );
NAND2_X1 MEM_stage_inst_dmem_U6273 ( .A1(MEM_stage_inst_dmem_ram_699), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n6145) );
NAND2_X1 MEM_stage_inst_dmem_U6272 ( .A1(MEM_stage_inst_dmem_n6143), .A2(MEM_stage_inst_dmem_n6142), .ZN(MEM_stage_inst_dmem_n6147) );
NAND2_X1 MEM_stage_inst_dmem_U6271 ( .A1(MEM_stage_inst_dmem_ram_971), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n6142) );
NAND2_X1 MEM_stage_inst_dmem_U6270 ( .A1(MEM_stage_inst_dmem_ram_763), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n6143) );
NAND2_X1 MEM_stage_inst_dmem_U6269 ( .A1(MEM_stage_inst_dmem_n6141), .A2(MEM_stage_inst_dmem_n6140), .ZN(MEM_stage_inst_dmem_n6205) );
NOR2_X1 MEM_stage_inst_dmem_U6268 ( .A1(MEM_stage_inst_dmem_n6139), .A2(MEM_stage_inst_dmem_n6138), .ZN(MEM_stage_inst_dmem_n6140) );
NAND2_X1 MEM_stage_inst_dmem_U6267 ( .A1(MEM_stage_inst_dmem_n6137), .A2(MEM_stage_inst_dmem_n6136), .ZN(MEM_stage_inst_dmem_n6138) );
NOR2_X1 MEM_stage_inst_dmem_U6266 ( .A1(MEM_stage_inst_dmem_n6135), .A2(MEM_stage_inst_dmem_n6134), .ZN(MEM_stage_inst_dmem_n6136) );
NAND2_X1 MEM_stage_inst_dmem_U6265 ( .A1(MEM_stage_inst_dmem_n6133), .A2(MEM_stage_inst_dmem_n6132), .ZN(MEM_stage_inst_dmem_n6134) );
NAND2_X1 MEM_stage_inst_dmem_U6264 ( .A1(MEM_stage_inst_dmem_ram_571), .A2(MEM_stage_inst_dmem_n8169), .ZN(MEM_stage_inst_dmem_n6132) );
NAND2_X1 MEM_stage_inst_dmem_U6263 ( .A1(MEM_stage_inst_dmem_ram_939), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n6133) );
NAND2_X1 MEM_stage_inst_dmem_U6262 ( .A1(MEM_stage_inst_dmem_n6131), .A2(MEM_stage_inst_dmem_n6130), .ZN(MEM_stage_inst_dmem_n6135) );
NAND2_X1 MEM_stage_inst_dmem_U6261 ( .A1(MEM_stage_inst_dmem_ram_1019), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n6130) );
NAND2_X1 MEM_stage_inst_dmem_U6260 ( .A1(MEM_stage_inst_dmem_ram_667), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n6131) );
NOR2_X1 MEM_stage_inst_dmem_U6259 ( .A1(MEM_stage_inst_dmem_n6129), .A2(MEM_stage_inst_dmem_n6128), .ZN(MEM_stage_inst_dmem_n6137) );
NAND2_X1 MEM_stage_inst_dmem_U6258 ( .A1(MEM_stage_inst_dmem_n6127), .A2(MEM_stage_inst_dmem_n6126), .ZN(MEM_stage_inst_dmem_n6128) );
NAND2_X1 MEM_stage_inst_dmem_U6257 ( .A1(MEM_stage_inst_dmem_ram_203), .A2(MEM_stage_inst_dmem_n8256), .ZN(MEM_stage_inst_dmem_n6126) );
NAND2_X1 MEM_stage_inst_dmem_U6256 ( .A1(MEM_stage_inst_dmem_ram_683), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n6127) );
NAND2_X1 MEM_stage_inst_dmem_U6255 ( .A1(MEM_stage_inst_dmem_n6125), .A2(MEM_stage_inst_dmem_n6124), .ZN(MEM_stage_inst_dmem_n6129) );
NAND2_X1 MEM_stage_inst_dmem_U6254 ( .A1(MEM_stage_inst_dmem_ram_523), .A2(MEM_stage_inst_dmem_n8225), .ZN(MEM_stage_inst_dmem_n6124) );
NAND2_X1 MEM_stage_inst_dmem_U6253 ( .A1(MEM_stage_inst_dmem_ram_107), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n6125) );
NAND2_X1 MEM_stage_inst_dmem_U6252 ( .A1(MEM_stage_inst_dmem_n6123), .A2(MEM_stage_inst_dmem_n6122), .ZN(MEM_stage_inst_dmem_n6139) );
NOR2_X1 MEM_stage_inst_dmem_U6251 ( .A1(MEM_stage_inst_dmem_n6121), .A2(MEM_stage_inst_dmem_n6120), .ZN(MEM_stage_inst_dmem_n6122) );
NAND2_X1 MEM_stage_inst_dmem_U6250 ( .A1(MEM_stage_inst_dmem_n6119), .A2(MEM_stage_inst_dmem_n6118), .ZN(MEM_stage_inst_dmem_n6120) );
NAND2_X1 MEM_stage_inst_dmem_U6249 ( .A1(MEM_stage_inst_dmem_ram_811), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n6118) );
NAND2_X1 MEM_stage_inst_dmem_U6248 ( .A1(MEM_stage_inst_dmem_ram_155), .A2(MEM_stage_inst_dmem_n7903), .ZN(MEM_stage_inst_dmem_n6119) );
NAND2_X1 MEM_stage_inst_dmem_U6247 ( .A1(MEM_stage_inst_dmem_n6117), .A2(MEM_stage_inst_dmem_n6116), .ZN(MEM_stage_inst_dmem_n6121) );
NAND2_X1 MEM_stage_inst_dmem_U6246 ( .A1(MEM_stage_inst_dmem_ram_331), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n6116) );
NAND2_X1 MEM_stage_inst_dmem_U6245 ( .A1(MEM_stage_inst_dmem_ram_427), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n6117) );
NOR2_X1 MEM_stage_inst_dmem_U6244 ( .A1(MEM_stage_inst_dmem_n6115), .A2(MEM_stage_inst_dmem_n6114), .ZN(MEM_stage_inst_dmem_n6123) );
NAND2_X1 MEM_stage_inst_dmem_U6243 ( .A1(MEM_stage_inst_dmem_n6113), .A2(MEM_stage_inst_dmem_n6112), .ZN(MEM_stage_inst_dmem_n6114) );
NAND2_X1 MEM_stage_inst_dmem_U6242 ( .A1(MEM_stage_inst_dmem_ram_779), .A2(MEM_stage_inst_dmem_n7992), .ZN(MEM_stage_inst_dmem_n6112) );
NAND2_X1 MEM_stage_inst_dmem_U6241 ( .A1(MEM_stage_inst_dmem_ram_171), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n6113) );
NAND2_X1 MEM_stage_inst_dmem_U6240 ( .A1(MEM_stage_inst_dmem_n6111), .A2(MEM_stage_inst_dmem_n6110), .ZN(MEM_stage_inst_dmem_n6115) );
NAND2_X1 MEM_stage_inst_dmem_U6239 ( .A1(MEM_stage_inst_dmem_ram_843), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n6110) );
NAND2_X1 MEM_stage_inst_dmem_U6238 ( .A1(MEM_stage_inst_dmem_ram_987), .A2(MEM_stage_inst_dmem_n7895), .ZN(MEM_stage_inst_dmem_n6111) );
NOR2_X1 MEM_stage_inst_dmem_U6237 ( .A1(MEM_stage_inst_dmem_n6109), .A2(MEM_stage_inst_dmem_n6108), .ZN(MEM_stage_inst_dmem_n6141) );
NAND2_X1 MEM_stage_inst_dmem_U6236 ( .A1(MEM_stage_inst_dmem_n6107), .A2(MEM_stage_inst_dmem_n6106), .ZN(MEM_stage_inst_dmem_n6108) );
NOR2_X1 MEM_stage_inst_dmem_U6235 ( .A1(MEM_stage_inst_dmem_n6105), .A2(MEM_stage_inst_dmem_n6104), .ZN(MEM_stage_inst_dmem_n6106) );
NAND2_X1 MEM_stage_inst_dmem_U6234 ( .A1(MEM_stage_inst_dmem_n6103), .A2(MEM_stage_inst_dmem_n6102), .ZN(MEM_stage_inst_dmem_n6104) );
NAND2_X1 MEM_stage_inst_dmem_U6233 ( .A1(MEM_stage_inst_dmem_ram_235), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n6102) );
NAND2_X1 MEM_stage_inst_dmem_U6232 ( .A1(MEM_stage_inst_dmem_ram_715), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n6103) );
NAND2_X1 MEM_stage_inst_dmem_U6231 ( .A1(MEM_stage_inst_dmem_n6101), .A2(MEM_stage_inst_dmem_n6100), .ZN(MEM_stage_inst_dmem_n6105) );
NAND2_X1 MEM_stage_inst_dmem_U6230 ( .A1(MEM_stage_inst_dmem_ram_315), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n6100) );
NAND2_X1 MEM_stage_inst_dmem_U6229 ( .A1(MEM_stage_inst_dmem_ram_91), .A2(MEM_stage_inst_dmem_n7938), .ZN(MEM_stage_inst_dmem_n6101) );
NOR2_X1 MEM_stage_inst_dmem_U6228 ( .A1(MEM_stage_inst_dmem_n6099), .A2(MEM_stage_inst_dmem_n6098), .ZN(MEM_stage_inst_dmem_n6107) );
NAND2_X1 MEM_stage_inst_dmem_U6227 ( .A1(MEM_stage_inst_dmem_n6097), .A2(MEM_stage_inst_dmem_n6096), .ZN(MEM_stage_inst_dmem_n6098) );
NAND2_X1 MEM_stage_inst_dmem_U6226 ( .A1(MEM_stage_inst_dmem_ram_475), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n6096) );
NAND2_X1 MEM_stage_inst_dmem_U6225 ( .A1(MEM_stage_inst_dmem_ram_395), .A2(MEM_stage_inst_dmem_n7930), .ZN(MEM_stage_inst_dmem_n6097) );
NAND2_X1 MEM_stage_inst_dmem_U6224 ( .A1(MEM_stage_inst_dmem_n6095), .A2(MEM_stage_inst_dmem_n6094), .ZN(MEM_stage_inst_dmem_n6099) );
NAND2_X1 MEM_stage_inst_dmem_U6223 ( .A1(MEM_stage_inst_dmem_ram_443), .A2(MEM_stage_inst_dmem_n7888), .ZN(MEM_stage_inst_dmem_n6094) );
NAND2_X1 MEM_stage_inst_dmem_U6222 ( .A1(MEM_stage_inst_dmem_ram_731), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n6095) );
NAND2_X1 MEM_stage_inst_dmem_U6221 ( .A1(MEM_stage_inst_dmem_n6093), .A2(MEM_stage_inst_dmem_n6092), .ZN(MEM_stage_inst_dmem_n6109) );
NOR2_X1 MEM_stage_inst_dmem_U6220 ( .A1(MEM_stage_inst_dmem_n6091), .A2(MEM_stage_inst_dmem_n6090), .ZN(MEM_stage_inst_dmem_n6092) );
NAND2_X1 MEM_stage_inst_dmem_U6219 ( .A1(MEM_stage_inst_dmem_n6089), .A2(MEM_stage_inst_dmem_n6088), .ZN(MEM_stage_inst_dmem_n6090) );
NAND2_X1 MEM_stage_inst_dmem_U6218 ( .A1(MEM_stage_inst_dmem_ram_619), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n6088) );
NAND2_X1 MEM_stage_inst_dmem_U6217 ( .A1(MEM_stage_inst_dmem_ram_539), .A2(MEM_stage_inst_dmem_n7884), .ZN(MEM_stage_inst_dmem_n6089) );
NAND2_X1 MEM_stage_inst_dmem_U6216 ( .A1(MEM_stage_inst_dmem_n6087), .A2(MEM_stage_inst_dmem_n6086), .ZN(MEM_stage_inst_dmem_n6091) );
NAND2_X1 MEM_stage_inst_dmem_U6215 ( .A1(MEM_stage_inst_dmem_ram_651), .A2(MEM_stage_inst_dmem_n7960), .ZN(MEM_stage_inst_dmem_n6086) );
NAND2_X1 MEM_stage_inst_dmem_U6214 ( .A1(MEM_stage_inst_dmem_ram_923), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n6087) );
NOR2_X1 MEM_stage_inst_dmem_U6213 ( .A1(MEM_stage_inst_dmem_n6085), .A2(MEM_stage_inst_dmem_n6084), .ZN(MEM_stage_inst_dmem_n6093) );
NAND2_X1 MEM_stage_inst_dmem_U6212 ( .A1(MEM_stage_inst_dmem_n6083), .A2(MEM_stage_inst_dmem_n6082), .ZN(MEM_stage_inst_dmem_n6084) );
NAND2_X1 MEM_stage_inst_dmem_U6211 ( .A1(MEM_stage_inst_dmem_ram_491), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n6082) );
NAND2_X1 MEM_stage_inst_dmem_U6210 ( .A1(MEM_stage_inst_dmem_ram_411), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n6083) );
NAND2_X1 MEM_stage_inst_dmem_U6209 ( .A1(MEM_stage_inst_dmem_n6081), .A2(MEM_stage_inst_dmem_n6080), .ZN(MEM_stage_inst_dmem_n6085) );
NAND2_X1 MEM_stage_inst_dmem_U6208 ( .A1(MEM_stage_inst_dmem_ram_907), .A2(MEM_stage_inst_dmem_n8193), .ZN(MEM_stage_inst_dmem_n6080) );
NAND2_X1 MEM_stage_inst_dmem_U6207 ( .A1(MEM_stage_inst_dmem_ram_747), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n6081) );
NOR2_X1 MEM_stage_inst_dmem_U6206 ( .A1(MEM_stage_inst_dmem_n6079), .A2(MEM_stage_inst_dmem_n8417), .ZN(MEM_stage_inst_dmem_n6208) );
NOR2_X1 MEM_stage_inst_dmem_U6205 ( .A1(MEM_stage_inst_dmem_n6078), .A2(MEM_stage_inst_dmem_n6077), .ZN(MEM_stage_inst_dmem_n6079) );
NAND2_X1 MEM_stage_inst_dmem_U6204 ( .A1(MEM_stage_inst_dmem_n6076), .A2(MEM_stage_inst_dmem_n6075), .ZN(MEM_stage_inst_dmem_n6077) );
NOR2_X1 MEM_stage_inst_dmem_U6203 ( .A1(MEM_stage_inst_dmem_n6074), .A2(MEM_stage_inst_dmem_n6073), .ZN(MEM_stage_inst_dmem_n6075) );
NAND2_X1 MEM_stage_inst_dmem_U6202 ( .A1(MEM_stage_inst_dmem_n6072), .A2(MEM_stage_inst_dmem_n6071), .ZN(MEM_stage_inst_dmem_n6073) );
NOR2_X1 MEM_stage_inst_dmem_U6201 ( .A1(MEM_stage_inst_dmem_n6070), .A2(MEM_stage_inst_dmem_n6069), .ZN(MEM_stage_inst_dmem_n6071) );
NAND2_X1 MEM_stage_inst_dmem_U6200 ( .A1(MEM_stage_inst_dmem_n6068), .A2(MEM_stage_inst_dmem_n6067), .ZN(MEM_stage_inst_dmem_n6069) );
NAND2_X1 MEM_stage_inst_dmem_U6199 ( .A1(MEM_stage_inst_dmem_ram_3563), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n6067) );
NAND2_X1 MEM_stage_inst_dmem_U6198 ( .A1(MEM_stage_inst_dmem_ram_3771), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n6068) );
NAND2_X1 MEM_stage_inst_dmem_U6197 ( .A1(MEM_stage_inst_dmem_n6066), .A2(MEM_stage_inst_dmem_n6065), .ZN(MEM_stage_inst_dmem_n6070) );
NAND2_X1 MEM_stage_inst_dmem_U6196 ( .A1(MEM_stage_inst_dmem_ram_3291), .A2(MEM_stage_inst_dmem_n8206), .ZN(MEM_stage_inst_dmem_n6065) );
NAND2_X1 MEM_stage_inst_dmem_U6195 ( .A1(MEM_stage_inst_dmem_ram_3179), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n6066) );
NOR2_X1 MEM_stage_inst_dmem_U6194 ( .A1(MEM_stage_inst_dmem_n6064), .A2(MEM_stage_inst_dmem_n6063), .ZN(MEM_stage_inst_dmem_n6072) );
NAND2_X1 MEM_stage_inst_dmem_U6193 ( .A1(MEM_stage_inst_dmem_n6062), .A2(MEM_stage_inst_dmem_n6061), .ZN(MEM_stage_inst_dmem_n6063) );
NAND2_X1 MEM_stage_inst_dmem_U6192 ( .A1(MEM_stage_inst_dmem_ram_3979), .A2(MEM_stage_inst_dmem_n8193), .ZN(MEM_stage_inst_dmem_n6061) );
NAND2_X1 MEM_stage_inst_dmem_U6191 ( .A1(MEM_stage_inst_dmem_ram_3547), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n6062) );
NAND2_X1 MEM_stage_inst_dmem_U6190 ( .A1(MEM_stage_inst_dmem_n6060), .A2(MEM_stage_inst_dmem_n6059), .ZN(MEM_stage_inst_dmem_n6064) );
NAND2_X1 MEM_stage_inst_dmem_U6189 ( .A1(MEM_stage_inst_dmem_ram_3755), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n6059) );
NAND2_X1 MEM_stage_inst_dmem_U6188 ( .A1(MEM_stage_inst_dmem_ram_4091), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n6060) );
NAND2_X1 MEM_stage_inst_dmem_U6187 ( .A1(MEM_stage_inst_dmem_n6058), .A2(MEM_stage_inst_dmem_n6057), .ZN(MEM_stage_inst_dmem_n6074) );
NOR2_X1 MEM_stage_inst_dmem_U6186 ( .A1(MEM_stage_inst_dmem_n6056), .A2(MEM_stage_inst_dmem_n6055), .ZN(MEM_stage_inst_dmem_n6057) );
NAND2_X1 MEM_stage_inst_dmem_U6185 ( .A1(MEM_stage_inst_dmem_n6054), .A2(MEM_stage_inst_dmem_n6053), .ZN(MEM_stage_inst_dmem_n6055) );
NAND2_X1 MEM_stage_inst_dmem_U6184 ( .A1(MEM_stage_inst_dmem_ram_3275), .A2(MEM_stage_inst_dmem_n8256), .ZN(MEM_stage_inst_dmem_n6053) );
NAND2_X1 MEM_stage_inst_dmem_U6183 ( .A1(MEM_stage_inst_dmem_ram_3915), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n6054) );
NAND2_X1 MEM_stage_inst_dmem_U6182 ( .A1(MEM_stage_inst_dmem_n6052), .A2(MEM_stage_inst_dmem_n6051), .ZN(MEM_stage_inst_dmem_n6056) );
NAND2_X1 MEM_stage_inst_dmem_U6181 ( .A1(MEM_stage_inst_dmem_ram_3403), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n6051) );
NAND2_X1 MEM_stage_inst_dmem_U6180 ( .A1(MEM_stage_inst_dmem_ram_4043), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n6052) );
NOR2_X1 MEM_stage_inst_dmem_U6179 ( .A1(MEM_stage_inst_dmem_n6050), .A2(MEM_stage_inst_dmem_n6049), .ZN(MEM_stage_inst_dmem_n6058) );
NAND2_X1 MEM_stage_inst_dmem_U6178 ( .A1(MEM_stage_inst_dmem_n6048), .A2(MEM_stage_inst_dmem_n6047), .ZN(MEM_stage_inst_dmem_n6049) );
NAND2_X1 MEM_stage_inst_dmem_U6177 ( .A1(MEM_stage_inst_dmem_ram_3883), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n6047) );
NAND2_X1 MEM_stage_inst_dmem_U6176 ( .A1(MEM_stage_inst_dmem_ram_3083), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n6048) );
NAND2_X1 MEM_stage_inst_dmem_U6175 ( .A1(MEM_stage_inst_dmem_n6046), .A2(MEM_stage_inst_dmem_n6045), .ZN(MEM_stage_inst_dmem_n6050) );
NAND2_X1 MEM_stage_inst_dmem_U6174 ( .A1(MEM_stage_inst_dmem_ram_4011), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n6045) );
NAND2_X1 MEM_stage_inst_dmem_U6173 ( .A1(MEM_stage_inst_dmem_ram_3707), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n6046) );
NOR2_X1 MEM_stage_inst_dmem_U6172 ( .A1(MEM_stage_inst_dmem_n6044), .A2(MEM_stage_inst_dmem_n6043), .ZN(MEM_stage_inst_dmem_n6076) );
NAND2_X1 MEM_stage_inst_dmem_U6171 ( .A1(MEM_stage_inst_dmem_n6042), .A2(MEM_stage_inst_dmem_n6041), .ZN(MEM_stage_inst_dmem_n6043) );
NOR2_X1 MEM_stage_inst_dmem_U6170 ( .A1(MEM_stage_inst_dmem_n6040), .A2(MEM_stage_inst_dmem_n6039), .ZN(MEM_stage_inst_dmem_n6041) );
NAND2_X1 MEM_stage_inst_dmem_U6169 ( .A1(MEM_stage_inst_dmem_n6038), .A2(MEM_stage_inst_dmem_n6037), .ZN(MEM_stage_inst_dmem_n6039) );
NAND2_X1 MEM_stage_inst_dmem_U6168 ( .A1(MEM_stage_inst_dmem_ram_3579), .A2(MEM_stage_inst_dmem_n64), .ZN(MEM_stage_inst_dmem_n6037) );
NAND2_X1 MEM_stage_inst_dmem_U6167 ( .A1(MEM_stage_inst_dmem_ram_3499), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n6038) );
NAND2_X1 MEM_stage_inst_dmem_U6166 ( .A1(MEM_stage_inst_dmem_n6036), .A2(MEM_stage_inst_dmem_n6035), .ZN(MEM_stage_inst_dmem_n6040) );
NAND2_X1 MEM_stage_inst_dmem_U6165 ( .A1(MEM_stage_inst_dmem_ram_3147), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n6035) );
NAND2_X1 MEM_stage_inst_dmem_U6164 ( .A1(MEM_stage_inst_dmem_ram_3163), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n6036) );
NOR2_X1 MEM_stage_inst_dmem_U6163 ( .A1(MEM_stage_inst_dmem_n6034), .A2(MEM_stage_inst_dmem_n6033), .ZN(MEM_stage_inst_dmem_n6042) );
NAND2_X1 MEM_stage_inst_dmem_U6162 ( .A1(MEM_stage_inst_dmem_n6032), .A2(MEM_stage_inst_dmem_n6031), .ZN(MEM_stage_inst_dmem_n6033) );
NAND2_X1 MEM_stage_inst_dmem_U6161 ( .A1(MEM_stage_inst_dmem_ram_3851), .A2(MEM_stage_inst_dmem_n8472), .ZN(MEM_stage_inst_dmem_n6031) );
NAND2_X1 MEM_stage_inst_dmem_U6160 ( .A1(MEM_stage_inst_dmem_ram_3131), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n6032) );
NAND2_X1 MEM_stage_inst_dmem_U6159 ( .A1(MEM_stage_inst_dmem_n6030), .A2(MEM_stage_inst_dmem_n6029), .ZN(MEM_stage_inst_dmem_n6034) );
NAND2_X1 MEM_stage_inst_dmem_U6158 ( .A1(MEM_stage_inst_dmem_ram_3947), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n6029) );
NAND2_X1 MEM_stage_inst_dmem_U6157 ( .A1(MEM_stage_inst_dmem_ram_3259), .A2(MEM_stage_inst_dmem_n8434), .ZN(MEM_stage_inst_dmem_n6030) );
NAND2_X1 MEM_stage_inst_dmem_U6156 ( .A1(MEM_stage_inst_dmem_n6028), .A2(MEM_stage_inst_dmem_n6027), .ZN(MEM_stage_inst_dmem_n6044) );
NOR2_X1 MEM_stage_inst_dmem_U6155 ( .A1(MEM_stage_inst_dmem_n6026), .A2(MEM_stage_inst_dmem_n6025), .ZN(MEM_stage_inst_dmem_n6027) );
NAND2_X1 MEM_stage_inst_dmem_U6154 ( .A1(MEM_stage_inst_dmem_n6024), .A2(MEM_stage_inst_dmem_n6023), .ZN(MEM_stage_inst_dmem_n6025) );
NAND2_X1 MEM_stage_inst_dmem_U6153 ( .A1(MEM_stage_inst_dmem_ram_3243), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n6023) );
NAND2_X1 MEM_stage_inst_dmem_U6152 ( .A1(MEM_stage_inst_dmem_ram_3659), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n6024) );
NAND2_X1 MEM_stage_inst_dmem_U6151 ( .A1(MEM_stage_inst_dmem_n6022), .A2(MEM_stage_inst_dmem_n6021), .ZN(MEM_stage_inst_dmem_n6026) );
NAND2_X1 MEM_stage_inst_dmem_U6150 ( .A1(MEM_stage_inst_dmem_ram_3115), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n6021) );
NAND2_X1 MEM_stage_inst_dmem_U6149 ( .A1(MEM_stage_inst_dmem_ram_3339), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n6022) );
NOR2_X1 MEM_stage_inst_dmem_U6148 ( .A1(MEM_stage_inst_dmem_n6020), .A2(MEM_stage_inst_dmem_n6019), .ZN(MEM_stage_inst_dmem_n6028) );
NAND2_X1 MEM_stage_inst_dmem_U6147 ( .A1(MEM_stage_inst_dmem_n6018), .A2(MEM_stage_inst_dmem_n6017), .ZN(MEM_stage_inst_dmem_n6019) );
NAND2_X1 MEM_stage_inst_dmem_U6146 ( .A1(MEM_stage_inst_dmem_ram_3963), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n6017) );
NAND2_X1 MEM_stage_inst_dmem_U6145 ( .A1(MEM_stage_inst_dmem_ram_3819), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n6018) );
NAND2_X1 MEM_stage_inst_dmem_U6144 ( .A1(MEM_stage_inst_dmem_n6016), .A2(MEM_stage_inst_dmem_n6015), .ZN(MEM_stage_inst_dmem_n6020) );
NAND2_X1 MEM_stage_inst_dmem_U6143 ( .A1(MEM_stage_inst_dmem_ram_3467), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n6015) );
NAND2_X1 MEM_stage_inst_dmem_U6142 ( .A1(MEM_stage_inst_dmem_ram_3611), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n6016) );
NAND2_X1 MEM_stage_inst_dmem_U6141 ( .A1(MEM_stage_inst_dmem_n6014), .A2(MEM_stage_inst_dmem_n6013), .ZN(MEM_stage_inst_dmem_n6078) );
NOR2_X1 MEM_stage_inst_dmem_U6140 ( .A1(MEM_stage_inst_dmem_n6012), .A2(MEM_stage_inst_dmem_n6011), .ZN(MEM_stage_inst_dmem_n6013) );
NAND2_X1 MEM_stage_inst_dmem_U6139 ( .A1(MEM_stage_inst_dmem_n6010), .A2(MEM_stage_inst_dmem_n6009), .ZN(MEM_stage_inst_dmem_n6011) );
NOR2_X1 MEM_stage_inst_dmem_U6138 ( .A1(MEM_stage_inst_dmem_n6008), .A2(MEM_stage_inst_dmem_n6007), .ZN(MEM_stage_inst_dmem_n6009) );
NAND2_X1 MEM_stage_inst_dmem_U6137 ( .A1(MEM_stage_inst_dmem_n6006), .A2(MEM_stage_inst_dmem_n6005), .ZN(MEM_stage_inst_dmem_n6007) );
NAND2_X1 MEM_stage_inst_dmem_U6136 ( .A1(MEM_stage_inst_dmem_ram_3435), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n6005) );
NAND2_X1 MEM_stage_inst_dmem_U6135 ( .A1(MEM_stage_inst_dmem_ram_3451), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n6006) );
NAND2_X1 MEM_stage_inst_dmem_U6134 ( .A1(MEM_stage_inst_dmem_n6004), .A2(MEM_stage_inst_dmem_n6003), .ZN(MEM_stage_inst_dmem_n6008) );
NAND2_X1 MEM_stage_inst_dmem_U6133 ( .A1(MEM_stage_inst_dmem_ram_3531), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n6003) );
NAND2_X1 MEM_stage_inst_dmem_U6132 ( .A1(MEM_stage_inst_dmem_ram_3803), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n6004) );
NOR2_X1 MEM_stage_inst_dmem_U6131 ( .A1(MEM_stage_inst_dmem_n6002), .A2(MEM_stage_inst_dmem_n6001), .ZN(MEM_stage_inst_dmem_n6010) );
NAND2_X1 MEM_stage_inst_dmem_U6130 ( .A1(MEM_stage_inst_dmem_n6000), .A2(MEM_stage_inst_dmem_n5999), .ZN(MEM_stage_inst_dmem_n6001) );
NAND2_X1 MEM_stage_inst_dmem_U6129 ( .A1(MEM_stage_inst_dmem_ram_3355), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n5999) );
NAND2_X1 MEM_stage_inst_dmem_U6128 ( .A1(MEM_stage_inst_dmem_ram_3675), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n6000) );
NAND2_X1 MEM_stage_inst_dmem_U6127 ( .A1(MEM_stage_inst_dmem_n5998), .A2(MEM_stage_inst_dmem_n5997), .ZN(MEM_stage_inst_dmem_n6002) );
NAND2_X1 MEM_stage_inst_dmem_U6126 ( .A1(MEM_stage_inst_dmem_ram_3899), .A2(MEM_stage_inst_dmem_n46), .ZN(MEM_stage_inst_dmem_n5997) );
NAND2_X1 MEM_stage_inst_dmem_U6125 ( .A1(MEM_stage_inst_dmem_ram_3195), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n5998) );
NAND2_X1 MEM_stage_inst_dmem_U6124 ( .A1(MEM_stage_inst_dmem_n5996), .A2(MEM_stage_inst_dmem_n5995), .ZN(MEM_stage_inst_dmem_n6012) );
NOR2_X1 MEM_stage_inst_dmem_U6123 ( .A1(MEM_stage_inst_dmem_n5994), .A2(MEM_stage_inst_dmem_n5993), .ZN(MEM_stage_inst_dmem_n5995) );
NAND2_X1 MEM_stage_inst_dmem_U6122 ( .A1(MEM_stage_inst_dmem_n5992), .A2(MEM_stage_inst_dmem_n5991), .ZN(MEM_stage_inst_dmem_n5993) );
NAND2_X1 MEM_stage_inst_dmem_U6121 ( .A1(MEM_stage_inst_dmem_ram_4027), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n5991) );
NAND2_X1 MEM_stage_inst_dmem_U6120 ( .A1(MEM_stage_inst_dmem_ram_3627), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n5992) );
NAND2_X1 MEM_stage_inst_dmem_U6119 ( .A1(MEM_stage_inst_dmem_n5990), .A2(MEM_stage_inst_dmem_n5989), .ZN(MEM_stage_inst_dmem_n5994) );
NAND2_X1 MEM_stage_inst_dmem_U6118 ( .A1(MEM_stage_inst_dmem_ram_3099), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n5989) );
NAND2_X1 MEM_stage_inst_dmem_U6117 ( .A1(MEM_stage_inst_dmem_ram_3739), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n5990) );
NOR2_X1 MEM_stage_inst_dmem_U6116 ( .A1(MEM_stage_inst_dmem_n5988), .A2(MEM_stage_inst_dmem_n5987), .ZN(MEM_stage_inst_dmem_n5996) );
NAND2_X1 MEM_stage_inst_dmem_U6115 ( .A1(MEM_stage_inst_dmem_n5986), .A2(MEM_stage_inst_dmem_n5985), .ZN(MEM_stage_inst_dmem_n5987) );
NAND2_X1 MEM_stage_inst_dmem_U6114 ( .A1(MEM_stage_inst_dmem_ram_3371), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n5985) );
NAND2_X1 MEM_stage_inst_dmem_U6113 ( .A1(MEM_stage_inst_dmem_ram_3595), .A2(MEM_stage_inst_dmem_n8225), .ZN(MEM_stage_inst_dmem_n5986) );
NAND2_X1 MEM_stage_inst_dmem_U6112 ( .A1(MEM_stage_inst_dmem_n5984), .A2(MEM_stage_inst_dmem_n5983), .ZN(MEM_stage_inst_dmem_n5988) );
NAND2_X1 MEM_stage_inst_dmem_U6111 ( .A1(MEM_stage_inst_dmem_ram_3643), .A2(MEM_stage_inst_dmem_n8169), .ZN(MEM_stage_inst_dmem_n5983) );
NAND2_X1 MEM_stage_inst_dmem_U6110 ( .A1(MEM_stage_inst_dmem_ram_4075), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n5984) );
NOR2_X1 MEM_stage_inst_dmem_U6109 ( .A1(MEM_stage_inst_dmem_n5982), .A2(MEM_stage_inst_dmem_n5981), .ZN(MEM_stage_inst_dmem_n6014) );
NAND2_X1 MEM_stage_inst_dmem_U6108 ( .A1(MEM_stage_inst_dmem_n5980), .A2(MEM_stage_inst_dmem_n5979), .ZN(MEM_stage_inst_dmem_n5981) );
NOR2_X1 MEM_stage_inst_dmem_U6107 ( .A1(MEM_stage_inst_dmem_n5978), .A2(MEM_stage_inst_dmem_n5977), .ZN(MEM_stage_inst_dmem_n5979) );
NAND2_X1 MEM_stage_inst_dmem_U6106 ( .A1(MEM_stage_inst_dmem_n5976), .A2(MEM_stage_inst_dmem_n5975), .ZN(MEM_stage_inst_dmem_n5977) );
NAND2_X1 MEM_stage_inst_dmem_U6105 ( .A1(MEM_stage_inst_dmem_ram_3995), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n5975) );
NAND2_X1 MEM_stage_inst_dmem_U6104 ( .A1(MEM_stage_inst_dmem_ram_3323), .A2(MEM_stage_inst_dmem_n39), .ZN(MEM_stage_inst_dmem_n5976) );
NAND2_X1 MEM_stage_inst_dmem_U6103 ( .A1(MEM_stage_inst_dmem_n5974), .A2(MEM_stage_inst_dmem_n5973), .ZN(MEM_stage_inst_dmem_n5978) );
NAND2_X1 MEM_stage_inst_dmem_U6102 ( .A1(MEM_stage_inst_dmem_ram_3387), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n5973) );
NAND2_X1 MEM_stage_inst_dmem_U6101 ( .A1(MEM_stage_inst_dmem_ram_3691), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n5974) );
NOR2_X1 MEM_stage_inst_dmem_U6100 ( .A1(MEM_stage_inst_dmem_n5972), .A2(MEM_stage_inst_dmem_n5971), .ZN(MEM_stage_inst_dmem_n5980) );
NAND2_X1 MEM_stage_inst_dmem_U6099 ( .A1(MEM_stage_inst_dmem_n5970), .A2(MEM_stage_inst_dmem_n5969), .ZN(MEM_stage_inst_dmem_n5971) );
NAND2_X1 MEM_stage_inst_dmem_U6098 ( .A1(MEM_stage_inst_dmem_ram_3723), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n5969) );
NAND2_X1 MEM_stage_inst_dmem_U6097 ( .A1(MEM_stage_inst_dmem_ram_3867), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n5970) );
NAND2_X1 MEM_stage_inst_dmem_U6096 ( .A1(MEM_stage_inst_dmem_n5968), .A2(MEM_stage_inst_dmem_n5967), .ZN(MEM_stage_inst_dmem_n5972) );
NAND2_X1 MEM_stage_inst_dmem_U6095 ( .A1(MEM_stage_inst_dmem_ram_3483), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n5967) );
NAND2_X1 MEM_stage_inst_dmem_U6094 ( .A1(MEM_stage_inst_dmem_ram_3419), .A2(MEM_stage_inst_dmem_n3216), .ZN(MEM_stage_inst_dmem_n5968) );
NAND2_X1 MEM_stage_inst_dmem_U6093 ( .A1(MEM_stage_inst_dmem_n5966), .A2(MEM_stage_inst_dmem_n5965), .ZN(MEM_stage_inst_dmem_n5982) );
NOR2_X1 MEM_stage_inst_dmem_U6092 ( .A1(MEM_stage_inst_dmem_n5964), .A2(MEM_stage_inst_dmem_n5963), .ZN(MEM_stage_inst_dmem_n5965) );
NAND2_X1 MEM_stage_inst_dmem_U6091 ( .A1(MEM_stage_inst_dmem_n5962), .A2(MEM_stage_inst_dmem_n5961), .ZN(MEM_stage_inst_dmem_n5963) );
NAND2_X1 MEM_stage_inst_dmem_U6090 ( .A1(MEM_stage_inst_dmem_ram_3307), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n5961) );
NAND2_X1 MEM_stage_inst_dmem_U6089 ( .A1(MEM_stage_inst_dmem_ram_3787), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n5962) );
NAND2_X1 MEM_stage_inst_dmem_U6088 ( .A1(MEM_stage_inst_dmem_n5960), .A2(MEM_stage_inst_dmem_n5959), .ZN(MEM_stage_inst_dmem_n5964) );
NAND2_X1 MEM_stage_inst_dmem_U6087 ( .A1(MEM_stage_inst_dmem_ram_3211), .A2(MEM_stage_inst_dmem_n8174), .ZN(MEM_stage_inst_dmem_n5959) );
NAND2_X1 MEM_stage_inst_dmem_U6086 ( .A1(MEM_stage_inst_dmem_ram_3227), .A2(MEM_stage_inst_dmem_n44), .ZN(MEM_stage_inst_dmem_n5960) );
NOR2_X1 MEM_stage_inst_dmem_U6085 ( .A1(MEM_stage_inst_dmem_n5958), .A2(MEM_stage_inst_dmem_n5957), .ZN(MEM_stage_inst_dmem_n5966) );
NAND2_X1 MEM_stage_inst_dmem_U6084 ( .A1(MEM_stage_inst_dmem_n5956), .A2(MEM_stage_inst_dmem_n5955), .ZN(MEM_stage_inst_dmem_n5957) );
NAND2_X1 MEM_stage_inst_dmem_U6083 ( .A1(MEM_stage_inst_dmem_ram_3931), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n5955) );
NAND2_X1 MEM_stage_inst_dmem_U6082 ( .A1(MEM_stage_inst_dmem_ram_3515), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n5956) );
NAND2_X1 MEM_stage_inst_dmem_U6081 ( .A1(MEM_stage_inst_dmem_n5954), .A2(MEM_stage_inst_dmem_n5953), .ZN(MEM_stage_inst_dmem_n5958) );
NAND2_X1 MEM_stage_inst_dmem_U6080 ( .A1(MEM_stage_inst_dmem_ram_3835), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n5953) );
NAND2_X1 MEM_stage_inst_dmem_U6079 ( .A1(MEM_stage_inst_dmem_ram_4059), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n5954) );
NAND2_X1 MEM_stage_inst_dmem_U6078 ( .A1(MEM_stage_inst_dmem_n5952), .A2(MEM_stage_inst_dmem_n5951), .ZN(MEM_stage_inst_mem_read_data_10) );
NOR2_X1 MEM_stage_inst_dmem_U6077 ( .A1(MEM_stage_inst_dmem_n5950), .A2(MEM_stage_inst_dmem_n5949), .ZN(MEM_stage_inst_dmem_n5951) );
NOR2_X1 MEM_stage_inst_dmem_U6076 ( .A1(MEM_stage_inst_dmem_n5948), .A2(MEM_stage_inst_dmem_n8152), .ZN(MEM_stage_inst_dmem_n5949) );
NOR2_X1 MEM_stage_inst_dmem_U6075 ( .A1(MEM_stage_inst_dmem_n5947), .A2(MEM_stage_inst_dmem_n5946), .ZN(MEM_stage_inst_dmem_n5948) );
NAND2_X1 MEM_stage_inst_dmem_U6074 ( .A1(MEM_stage_inst_dmem_n5945), .A2(MEM_stage_inst_dmem_n5944), .ZN(MEM_stage_inst_dmem_n5946) );
NOR2_X1 MEM_stage_inst_dmem_U6073 ( .A1(MEM_stage_inst_dmem_n5943), .A2(MEM_stage_inst_dmem_n5942), .ZN(MEM_stage_inst_dmem_n5944) );
NAND2_X1 MEM_stage_inst_dmem_U6072 ( .A1(MEM_stage_inst_dmem_n5941), .A2(MEM_stage_inst_dmem_n5940), .ZN(MEM_stage_inst_dmem_n5942) );
NOR2_X1 MEM_stage_inst_dmem_U6071 ( .A1(MEM_stage_inst_dmem_n5939), .A2(MEM_stage_inst_dmem_n5938), .ZN(MEM_stage_inst_dmem_n5940) );
NAND2_X1 MEM_stage_inst_dmem_U6070 ( .A1(MEM_stage_inst_dmem_n5937), .A2(MEM_stage_inst_dmem_n5936), .ZN(MEM_stage_inst_dmem_n5938) );
NAND2_X1 MEM_stage_inst_dmem_U6069 ( .A1(MEM_stage_inst_dmem_ram_1402), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n5936) );
NAND2_X1 MEM_stage_inst_dmem_U6068 ( .A1(MEM_stage_inst_dmem_ram_1690), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n5937) );
NAND2_X1 MEM_stage_inst_dmem_U6067 ( .A1(MEM_stage_inst_dmem_n5935), .A2(MEM_stage_inst_dmem_n5934), .ZN(MEM_stage_inst_dmem_n5939) );
NAND2_X1 MEM_stage_inst_dmem_U6066 ( .A1(MEM_stage_inst_dmem_ram_1338), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n5934) );
NAND2_X1 MEM_stage_inst_dmem_U6065 ( .A1(MEM_stage_inst_dmem_ram_1994), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n5935) );
NOR2_X1 MEM_stage_inst_dmem_U6064 ( .A1(MEM_stage_inst_dmem_n5933), .A2(MEM_stage_inst_dmem_n5932), .ZN(MEM_stage_inst_dmem_n5941) );
NAND2_X1 MEM_stage_inst_dmem_U6063 ( .A1(MEM_stage_inst_dmem_n5931), .A2(MEM_stage_inst_dmem_n5930), .ZN(MEM_stage_inst_dmem_n5932) );
NAND2_X1 MEM_stage_inst_dmem_U6062 ( .A1(MEM_stage_inst_dmem_ram_1306), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n5930) );
NAND2_X1 MEM_stage_inst_dmem_U6061 ( .A1(MEM_stage_inst_dmem_ram_1658), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n5931) );
NAND2_X1 MEM_stage_inst_dmem_U6060 ( .A1(MEM_stage_inst_dmem_n5929), .A2(MEM_stage_inst_dmem_n5928), .ZN(MEM_stage_inst_dmem_n5933) );
NAND2_X1 MEM_stage_inst_dmem_U6059 ( .A1(MEM_stage_inst_dmem_ram_1098), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n5928) );
NAND2_X1 MEM_stage_inst_dmem_U6058 ( .A1(MEM_stage_inst_dmem_ram_1162), .A2(MEM_stage_inst_dmem_n8174), .ZN(MEM_stage_inst_dmem_n5929) );
NAND2_X1 MEM_stage_inst_dmem_U6057 ( .A1(MEM_stage_inst_dmem_n5927), .A2(MEM_stage_inst_dmem_n5926), .ZN(MEM_stage_inst_dmem_n5943) );
NOR2_X1 MEM_stage_inst_dmem_U6056 ( .A1(MEM_stage_inst_dmem_n5925), .A2(MEM_stage_inst_dmem_n5924), .ZN(MEM_stage_inst_dmem_n5926) );
NAND2_X1 MEM_stage_inst_dmem_U6055 ( .A1(MEM_stage_inst_dmem_n5923), .A2(MEM_stage_inst_dmem_n5922), .ZN(MEM_stage_inst_dmem_n5924) );
NAND2_X1 MEM_stage_inst_dmem_U6054 ( .A1(MEM_stage_inst_dmem_ram_1738), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n5922) );
NAND2_X1 MEM_stage_inst_dmem_U6053 ( .A1(MEM_stage_inst_dmem_ram_1242), .A2(MEM_stage_inst_dmem_n8206), .ZN(MEM_stage_inst_dmem_n5923) );
NAND2_X1 MEM_stage_inst_dmem_U6052 ( .A1(MEM_stage_inst_dmem_n5921), .A2(MEM_stage_inst_dmem_n5920), .ZN(MEM_stage_inst_dmem_n5925) );
NAND2_X1 MEM_stage_inst_dmem_U6051 ( .A1(MEM_stage_inst_dmem_ram_1258), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n5920) );
NAND2_X1 MEM_stage_inst_dmem_U6050 ( .A1(MEM_stage_inst_dmem_ram_2042), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n5921) );
NOR2_X1 MEM_stage_inst_dmem_U6049 ( .A1(MEM_stage_inst_dmem_n5919), .A2(MEM_stage_inst_dmem_n5918), .ZN(MEM_stage_inst_dmem_n5927) );
NAND2_X1 MEM_stage_inst_dmem_U6048 ( .A1(MEM_stage_inst_dmem_n5917), .A2(MEM_stage_inst_dmem_n5916), .ZN(MEM_stage_inst_dmem_n5918) );
NAND2_X1 MEM_stage_inst_dmem_U6047 ( .A1(MEM_stage_inst_dmem_ram_1194), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n5916) );
NAND2_X1 MEM_stage_inst_dmem_U6046 ( .A1(MEM_stage_inst_dmem_ram_1034), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n5917) );
NAND2_X1 MEM_stage_inst_dmem_U6045 ( .A1(MEM_stage_inst_dmem_n5915), .A2(MEM_stage_inst_dmem_n5914), .ZN(MEM_stage_inst_dmem_n5919) );
NAND2_X1 MEM_stage_inst_dmem_U6044 ( .A1(MEM_stage_inst_dmem_ram_1898), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n5914) );
NAND2_X1 MEM_stage_inst_dmem_U6043 ( .A1(MEM_stage_inst_dmem_ram_1802), .A2(MEM_stage_inst_dmem_n37), .ZN(MEM_stage_inst_dmem_n5915) );
NOR2_X1 MEM_stage_inst_dmem_U6042 ( .A1(MEM_stage_inst_dmem_n5913), .A2(MEM_stage_inst_dmem_n5912), .ZN(MEM_stage_inst_dmem_n5945) );
NAND2_X1 MEM_stage_inst_dmem_U6041 ( .A1(MEM_stage_inst_dmem_n5911), .A2(MEM_stage_inst_dmem_n5910), .ZN(MEM_stage_inst_dmem_n5912) );
NOR2_X1 MEM_stage_inst_dmem_U6040 ( .A1(MEM_stage_inst_dmem_n5909), .A2(MEM_stage_inst_dmem_n5908), .ZN(MEM_stage_inst_dmem_n5910) );
NAND2_X1 MEM_stage_inst_dmem_U6039 ( .A1(MEM_stage_inst_dmem_n5907), .A2(MEM_stage_inst_dmem_n5906), .ZN(MEM_stage_inst_dmem_n5908) );
NAND2_X1 MEM_stage_inst_dmem_U6038 ( .A1(MEM_stage_inst_dmem_ram_1946), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n5906) );
NAND2_X1 MEM_stage_inst_dmem_U6037 ( .A1(MEM_stage_inst_dmem_ram_1770), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n5907) );
NAND2_X1 MEM_stage_inst_dmem_U6036 ( .A1(MEM_stage_inst_dmem_n5905), .A2(MEM_stage_inst_dmem_n5904), .ZN(MEM_stage_inst_dmem_n5909) );
NAND2_X1 MEM_stage_inst_dmem_U6035 ( .A1(MEM_stage_inst_dmem_ram_1674), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n5904) );
NAND2_X1 MEM_stage_inst_dmem_U6034 ( .A1(MEM_stage_inst_dmem_ram_1146), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n5905) );
NOR2_X1 MEM_stage_inst_dmem_U6033 ( .A1(MEM_stage_inst_dmem_n5903), .A2(MEM_stage_inst_dmem_n5902), .ZN(MEM_stage_inst_dmem_n5911) );
NAND2_X1 MEM_stage_inst_dmem_U6032 ( .A1(MEM_stage_inst_dmem_n5901), .A2(MEM_stage_inst_dmem_n5900), .ZN(MEM_stage_inst_dmem_n5902) );
NAND2_X1 MEM_stage_inst_dmem_U6031 ( .A1(MEM_stage_inst_dmem_ram_1882), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n5900) );
NAND2_X1 MEM_stage_inst_dmem_U6030 ( .A1(MEM_stage_inst_dmem_ram_1130), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n5901) );
NAND2_X1 MEM_stage_inst_dmem_U6029 ( .A1(MEM_stage_inst_dmem_n5899), .A2(MEM_stage_inst_dmem_n5898), .ZN(MEM_stage_inst_dmem_n5903) );
NAND2_X1 MEM_stage_inst_dmem_U6028 ( .A1(MEM_stage_inst_dmem_ram_1434), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n5898) );
NAND2_X1 MEM_stage_inst_dmem_U6027 ( .A1(MEM_stage_inst_dmem_ram_1786), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n5899) );
NAND2_X1 MEM_stage_inst_dmem_U6026 ( .A1(MEM_stage_inst_dmem_n5897), .A2(MEM_stage_inst_dmem_n5896), .ZN(MEM_stage_inst_dmem_n5913) );
NOR2_X1 MEM_stage_inst_dmem_U6025 ( .A1(MEM_stage_inst_dmem_n5895), .A2(MEM_stage_inst_dmem_n5894), .ZN(MEM_stage_inst_dmem_n5896) );
NAND2_X1 MEM_stage_inst_dmem_U6024 ( .A1(MEM_stage_inst_dmem_n5893), .A2(MEM_stage_inst_dmem_n5892), .ZN(MEM_stage_inst_dmem_n5894) );
NAND2_X1 MEM_stage_inst_dmem_U6023 ( .A1(MEM_stage_inst_dmem_ram_1386), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n5892) );
NAND2_X1 MEM_stage_inst_dmem_U6022 ( .A1(MEM_stage_inst_dmem_ram_1706), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n5893) );
NAND2_X1 MEM_stage_inst_dmem_U6021 ( .A1(MEM_stage_inst_dmem_n5891), .A2(MEM_stage_inst_dmem_n5890), .ZN(MEM_stage_inst_dmem_n5895) );
NAND2_X1 MEM_stage_inst_dmem_U6020 ( .A1(MEM_stage_inst_dmem_ram_1834), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n5890) );
NAND2_X1 MEM_stage_inst_dmem_U6019 ( .A1(MEM_stage_inst_dmem_ram_1642), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n5891) );
NOR2_X1 MEM_stage_inst_dmem_U6018 ( .A1(MEM_stage_inst_dmem_n5889), .A2(MEM_stage_inst_dmem_n5888), .ZN(MEM_stage_inst_dmem_n5897) );
NAND2_X1 MEM_stage_inst_dmem_U6017 ( .A1(MEM_stage_inst_dmem_n5887), .A2(MEM_stage_inst_dmem_n5886), .ZN(MEM_stage_inst_dmem_n5888) );
NAND2_X1 MEM_stage_inst_dmem_U6016 ( .A1(MEM_stage_inst_dmem_ram_1418), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n5886) );
NAND2_X1 MEM_stage_inst_dmem_U6015 ( .A1(MEM_stage_inst_dmem_ram_1370), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n5887) );
NAND2_X1 MEM_stage_inst_dmem_U6014 ( .A1(MEM_stage_inst_dmem_n5885), .A2(MEM_stage_inst_dmem_n5884), .ZN(MEM_stage_inst_dmem_n5889) );
NAND2_X1 MEM_stage_inst_dmem_U6013 ( .A1(MEM_stage_inst_dmem_ram_1914), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n5884) );
NAND2_X1 MEM_stage_inst_dmem_U6012 ( .A1(MEM_stage_inst_dmem_ram_1114), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n5885) );
NAND2_X1 MEM_stage_inst_dmem_U6011 ( .A1(MEM_stage_inst_dmem_n5883), .A2(MEM_stage_inst_dmem_n5882), .ZN(MEM_stage_inst_dmem_n5947) );
NOR2_X1 MEM_stage_inst_dmem_U6010 ( .A1(MEM_stage_inst_dmem_n5881), .A2(MEM_stage_inst_dmem_n5880), .ZN(MEM_stage_inst_dmem_n5882) );
NAND2_X1 MEM_stage_inst_dmem_U6009 ( .A1(MEM_stage_inst_dmem_n5879), .A2(MEM_stage_inst_dmem_n5878), .ZN(MEM_stage_inst_dmem_n5880) );
NOR2_X1 MEM_stage_inst_dmem_U6008 ( .A1(MEM_stage_inst_dmem_n5877), .A2(MEM_stage_inst_dmem_n5876), .ZN(MEM_stage_inst_dmem_n5878) );
NAND2_X1 MEM_stage_inst_dmem_U6007 ( .A1(MEM_stage_inst_dmem_n5875), .A2(MEM_stage_inst_dmem_n5874), .ZN(MEM_stage_inst_dmem_n5876) );
NAND2_X1 MEM_stage_inst_dmem_U6006 ( .A1(MEM_stage_inst_dmem_ram_1450), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n5874) );
NAND2_X1 MEM_stage_inst_dmem_U6005 ( .A1(MEM_stage_inst_dmem_ram_1210), .A2(MEM_stage_inst_dmem_n55), .ZN(MEM_stage_inst_dmem_n5875) );
NAND2_X1 MEM_stage_inst_dmem_U6004 ( .A1(MEM_stage_inst_dmem_n5873), .A2(MEM_stage_inst_dmem_n5872), .ZN(MEM_stage_inst_dmem_n5877) );
NAND2_X1 MEM_stage_inst_dmem_U6003 ( .A1(MEM_stage_inst_dmem_ram_1082), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n5872) );
NAND2_X1 MEM_stage_inst_dmem_U6002 ( .A1(MEM_stage_inst_dmem_ram_1178), .A2(MEM_stage_inst_dmem_n44), .ZN(MEM_stage_inst_dmem_n5873) );
NOR2_X1 MEM_stage_inst_dmem_U6001 ( .A1(MEM_stage_inst_dmem_n5871), .A2(MEM_stage_inst_dmem_n5870), .ZN(MEM_stage_inst_dmem_n5879) );
NAND2_X1 MEM_stage_inst_dmem_U6000 ( .A1(MEM_stage_inst_dmem_n5869), .A2(MEM_stage_inst_dmem_n5868), .ZN(MEM_stage_inst_dmem_n5870) );
NAND2_X1 MEM_stage_inst_dmem_U5999 ( .A1(MEM_stage_inst_dmem_ram_1578), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n5868) );
NAND2_X1 MEM_stage_inst_dmem_U5998 ( .A1(MEM_stage_inst_dmem_ram_1962), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n5869) );
NAND2_X1 MEM_stage_inst_dmem_U5997 ( .A1(MEM_stage_inst_dmem_n5867), .A2(MEM_stage_inst_dmem_n5866), .ZN(MEM_stage_inst_dmem_n5871) );
NAND2_X1 MEM_stage_inst_dmem_U5996 ( .A1(MEM_stage_inst_dmem_ram_1466), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n5866) );
NAND2_X1 MEM_stage_inst_dmem_U5995 ( .A1(MEM_stage_inst_dmem_ram_1594), .A2(MEM_stage_inst_dmem_n8169), .ZN(MEM_stage_inst_dmem_n5867) );
NAND2_X1 MEM_stage_inst_dmem_U5994 ( .A1(MEM_stage_inst_dmem_n5865), .A2(MEM_stage_inst_dmem_n5864), .ZN(MEM_stage_inst_dmem_n5881) );
NOR2_X1 MEM_stage_inst_dmem_U5993 ( .A1(MEM_stage_inst_dmem_n5863), .A2(MEM_stage_inst_dmem_n5862), .ZN(MEM_stage_inst_dmem_n5864) );
NAND2_X1 MEM_stage_inst_dmem_U5992 ( .A1(MEM_stage_inst_dmem_n5861), .A2(MEM_stage_inst_dmem_n5860), .ZN(MEM_stage_inst_dmem_n5862) );
NAND2_X1 MEM_stage_inst_dmem_U5991 ( .A1(MEM_stage_inst_dmem_ram_2026), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n5860) );
NAND2_X1 MEM_stage_inst_dmem_U5990 ( .A1(MEM_stage_inst_dmem_ram_1818), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n5861) );
NAND2_X1 MEM_stage_inst_dmem_U5989 ( .A1(MEM_stage_inst_dmem_n5859), .A2(MEM_stage_inst_dmem_n5858), .ZN(MEM_stage_inst_dmem_n5863) );
NAND2_X1 MEM_stage_inst_dmem_U5988 ( .A1(MEM_stage_inst_dmem_ram_1354), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n5858) );
NAND2_X1 MEM_stage_inst_dmem_U5987 ( .A1(MEM_stage_inst_dmem_ram_1290), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n5859) );
NOR2_X1 MEM_stage_inst_dmem_U5986 ( .A1(MEM_stage_inst_dmem_n5856), .A2(MEM_stage_inst_dmem_n5855), .ZN(MEM_stage_inst_dmem_n5865) );
NAND2_X1 MEM_stage_inst_dmem_U5985 ( .A1(MEM_stage_inst_dmem_n5854), .A2(MEM_stage_inst_dmem_n5853), .ZN(MEM_stage_inst_dmem_n5855) );
NAND2_X1 MEM_stage_inst_dmem_U5984 ( .A1(MEM_stage_inst_dmem_ram_1274), .A2(MEM_stage_inst_dmem_n39), .ZN(MEM_stage_inst_dmem_n5853) );
NAND2_X1 MEM_stage_inst_dmem_U5983 ( .A1(MEM_stage_inst_dmem_ram_1850), .A2(MEM_stage_inst_dmem_n46), .ZN(MEM_stage_inst_dmem_n5854) );
NAND2_X1 MEM_stage_inst_dmem_U5982 ( .A1(MEM_stage_inst_dmem_n5852), .A2(MEM_stage_inst_dmem_n5851), .ZN(MEM_stage_inst_dmem_n5856) );
NAND2_X1 MEM_stage_inst_dmem_U5981 ( .A1(MEM_stage_inst_dmem_ram_1322), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n5851) );
NAND2_X1 MEM_stage_inst_dmem_U5980 ( .A1(MEM_stage_inst_dmem_ram_1626), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n5852) );
NOR2_X1 MEM_stage_inst_dmem_U5979 ( .A1(MEM_stage_inst_dmem_n5850), .A2(MEM_stage_inst_dmem_n5849), .ZN(MEM_stage_inst_dmem_n5883) );
NAND2_X1 MEM_stage_inst_dmem_U5978 ( .A1(MEM_stage_inst_dmem_n5848), .A2(MEM_stage_inst_dmem_n5847), .ZN(MEM_stage_inst_dmem_n5849) );
NOR2_X1 MEM_stage_inst_dmem_U5977 ( .A1(MEM_stage_inst_dmem_n5846), .A2(MEM_stage_inst_dmem_n5845), .ZN(MEM_stage_inst_dmem_n5847) );
NAND2_X1 MEM_stage_inst_dmem_U5976 ( .A1(MEM_stage_inst_dmem_n5844), .A2(MEM_stage_inst_dmem_n5843), .ZN(MEM_stage_inst_dmem_n5845) );
NAND2_X1 MEM_stage_inst_dmem_U5975 ( .A1(MEM_stage_inst_dmem_ram_1866), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n5843) );
NAND2_X1 MEM_stage_inst_dmem_U5974 ( .A1(MEM_stage_inst_dmem_ram_1978), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n5844) );
NAND2_X1 MEM_stage_inst_dmem_U5973 ( .A1(MEM_stage_inst_dmem_n5842), .A2(MEM_stage_inst_dmem_n5841), .ZN(MEM_stage_inst_dmem_n5846) );
NAND2_X1 MEM_stage_inst_dmem_U5972 ( .A1(MEM_stage_inst_dmem_ram_1226), .A2(MEM_stage_inst_dmem_n8256), .ZN(MEM_stage_inst_dmem_n5841) );
NAND2_X1 MEM_stage_inst_dmem_U5971 ( .A1(MEM_stage_inst_dmem_ram_1754), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n5842) );
NOR2_X1 MEM_stage_inst_dmem_U5970 ( .A1(MEM_stage_inst_dmem_n5840), .A2(MEM_stage_inst_dmem_n5839), .ZN(MEM_stage_inst_dmem_n5848) );
NAND2_X1 MEM_stage_inst_dmem_U5969 ( .A1(MEM_stage_inst_dmem_n5838), .A2(MEM_stage_inst_dmem_n5837), .ZN(MEM_stage_inst_dmem_n5839) );
NAND2_X1 MEM_stage_inst_dmem_U5968 ( .A1(MEM_stage_inst_dmem_ram_1498), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n5837) );
NAND2_X1 MEM_stage_inst_dmem_U5967 ( .A1(MEM_stage_inst_dmem_ram_1610), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n5838) );
NAND2_X1 MEM_stage_inst_dmem_U5966 ( .A1(MEM_stage_inst_dmem_n5836), .A2(MEM_stage_inst_dmem_n5835), .ZN(MEM_stage_inst_dmem_n5840) );
NAND2_X1 MEM_stage_inst_dmem_U5965 ( .A1(MEM_stage_inst_dmem_ram_1066), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n5835) );
NAND2_X1 MEM_stage_inst_dmem_U5964 ( .A1(MEM_stage_inst_dmem_ram_1722), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n5836) );
NAND2_X1 MEM_stage_inst_dmem_U5963 ( .A1(MEM_stage_inst_dmem_n5834), .A2(MEM_stage_inst_dmem_n5833), .ZN(MEM_stage_inst_dmem_n5850) );
NOR2_X1 MEM_stage_inst_dmem_U5962 ( .A1(MEM_stage_inst_dmem_n5832), .A2(MEM_stage_inst_dmem_n5831), .ZN(MEM_stage_inst_dmem_n5833) );
NAND2_X1 MEM_stage_inst_dmem_U5961 ( .A1(MEM_stage_inst_dmem_n5830), .A2(MEM_stage_inst_dmem_n5829), .ZN(MEM_stage_inst_dmem_n5831) );
NAND2_X1 MEM_stage_inst_dmem_U5960 ( .A1(MEM_stage_inst_dmem_ram_1530), .A2(MEM_stage_inst_dmem_n64), .ZN(MEM_stage_inst_dmem_n5829) );
NAND2_X1 MEM_stage_inst_dmem_U5959 ( .A1(MEM_stage_inst_dmem_ram_1050), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n5830) );
NAND2_X1 MEM_stage_inst_dmem_U5958 ( .A1(MEM_stage_inst_dmem_n5828), .A2(MEM_stage_inst_dmem_n5827), .ZN(MEM_stage_inst_dmem_n5832) );
NAND2_X1 MEM_stage_inst_dmem_U5957 ( .A1(MEM_stage_inst_dmem_ram_1930), .A2(MEM_stage_inst_dmem_n8193), .ZN(MEM_stage_inst_dmem_n5827) );
NAND2_X1 MEM_stage_inst_dmem_U5956 ( .A1(MEM_stage_inst_dmem_ram_1482), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n5828) );
NOR2_X1 MEM_stage_inst_dmem_U5955 ( .A1(MEM_stage_inst_dmem_n5826), .A2(MEM_stage_inst_dmem_n5825), .ZN(MEM_stage_inst_dmem_n5834) );
NAND2_X1 MEM_stage_inst_dmem_U5954 ( .A1(MEM_stage_inst_dmem_n5824), .A2(MEM_stage_inst_dmem_n5823), .ZN(MEM_stage_inst_dmem_n5825) );
NAND2_X1 MEM_stage_inst_dmem_U5953 ( .A1(MEM_stage_inst_dmem_ram_1514), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n5823) );
NAND2_X1 MEM_stage_inst_dmem_U5952 ( .A1(MEM_stage_inst_dmem_ram_1546), .A2(MEM_stage_inst_dmem_n8225), .ZN(MEM_stage_inst_dmem_n5824) );
NAND2_X1 MEM_stage_inst_dmem_U5951 ( .A1(MEM_stage_inst_dmem_n5822), .A2(MEM_stage_inst_dmem_n5821), .ZN(MEM_stage_inst_dmem_n5826) );
NAND2_X1 MEM_stage_inst_dmem_U5950 ( .A1(MEM_stage_inst_dmem_ram_2010), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n5821) );
NAND2_X1 MEM_stage_inst_dmem_U5949 ( .A1(MEM_stage_inst_dmem_ram_1562), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n5822) );
NOR2_X1 MEM_stage_inst_dmem_U5948 ( .A1(MEM_stage_inst_dmem_n5820), .A2(MEM_stage_inst_dmem_n8551), .ZN(MEM_stage_inst_dmem_n5950) );
NOR2_X1 MEM_stage_inst_dmem_U5947 ( .A1(MEM_stage_inst_dmem_n5819), .A2(MEM_stage_inst_dmem_n5818), .ZN(MEM_stage_inst_dmem_n5820) );
NAND2_X1 MEM_stage_inst_dmem_U5946 ( .A1(MEM_stage_inst_dmem_n5817), .A2(MEM_stage_inst_dmem_n5816), .ZN(MEM_stage_inst_dmem_n5818) );
NOR2_X1 MEM_stage_inst_dmem_U5945 ( .A1(MEM_stage_inst_dmem_n5815), .A2(MEM_stage_inst_dmem_n5814), .ZN(MEM_stage_inst_dmem_n5816) );
NAND2_X1 MEM_stage_inst_dmem_U5944 ( .A1(MEM_stage_inst_dmem_n5813), .A2(MEM_stage_inst_dmem_n5812), .ZN(MEM_stage_inst_dmem_n5814) );
NOR2_X1 MEM_stage_inst_dmem_U5943 ( .A1(MEM_stage_inst_dmem_n5811), .A2(MEM_stage_inst_dmem_n5810), .ZN(MEM_stage_inst_dmem_n5812) );
NAND2_X1 MEM_stage_inst_dmem_U5942 ( .A1(MEM_stage_inst_dmem_n5809), .A2(MEM_stage_inst_dmem_n5808), .ZN(MEM_stage_inst_dmem_n5810) );
NAND2_X1 MEM_stage_inst_dmem_U5941 ( .A1(MEM_stage_inst_dmem_ram_154), .A2(MEM_stage_inst_dmem_n5807), .ZN(MEM_stage_inst_dmem_n5808) );
NAND2_X1 MEM_stage_inst_dmem_U5940 ( .A1(MEM_stage_inst_dmem_ram_186), .A2(MEM_stage_inst_dmem_n55), .ZN(MEM_stage_inst_dmem_n5809) );
NAND2_X1 MEM_stage_inst_dmem_U5939 ( .A1(MEM_stage_inst_dmem_n5806), .A2(MEM_stage_inst_dmem_n5805), .ZN(MEM_stage_inst_dmem_n5811) );
NAND2_X1 MEM_stage_inst_dmem_U5938 ( .A1(MEM_stage_inst_dmem_ram_762), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n5805) );
NAND2_X1 MEM_stage_inst_dmem_U5937 ( .A1(MEM_stage_inst_dmem_ram_266), .A2(MEM_stage_inst_dmem_n7898), .ZN(MEM_stage_inst_dmem_n5806) );
NOR2_X1 MEM_stage_inst_dmem_U5936 ( .A1(MEM_stage_inst_dmem_n5804), .A2(MEM_stage_inst_dmem_n5803), .ZN(MEM_stage_inst_dmem_n5813) );
NAND2_X1 MEM_stage_inst_dmem_U5935 ( .A1(MEM_stage_inst_dmem_n5802), .A2(MEM_stage_inst_dmem_n5801), .ZN(MEM_stage_inst_dmem_n5803) );
NAND2_X1 MEM_stage_inst_dmem_U5934 ( .A1(MEM_stage_inst_dmem_ram_378), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n5801) );
NAND2_X1 MEM_stage_inst_dmem_U5933 ( .A1(MEM_stage_inst_dmem_ram_666), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n5802) );
NAND2_X1 MEM_stage_inst_dmem_U5932 ( .A1(MEM_stage_inst_dmem_n5800), .A2(MEM_stage_inst_dmem_n5799), .ZN(MEM_stage_inst_dmem_n5804) );
NAND2_X1 MEM_stage_inst_dmem_U5931 ( .A1(MEM_stage_inst_dmem_ram_234), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n5799) );
NAND2_X1 MEM_stage_inst_dmem_U5930 ( .A1(MEM_stage_inst_dmem_ram_1018), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n5800) );
NAND2_X1 MEM_stage_inst_dmem_U5929 ( .A1(MEM_stage_inst_dmem_n5798), .A2(MEM_stage_inst_dmem_n5797), .ZN(MEM_stage_inst_dmem_n5815) );
NOR2_X1 MEM_stage_inst_dmem_U5928 ( .A1(MEM_stage_inst_dmem_n5796), .A2(MEM_stage_inst_dmem_n5795), .ZN(MEM_stage_inst_dmem_n5797) );
NAND2_X1 MEM_stage_inst_dmem_U5927 ( .A1(MEM_stage_inst_dmem_n5794), .A2(MEM_stage_inst_dmem_n5793), .ZN(MEM_stage_inst_dmem_n5795) );
NAND2_X1 MEM_stage_inst_dmem_U5926 ( .A1(MEM_stage_inst_dmem_ram_474), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n5793) );
NAND2_X1 MEM_stage_inst_dmem_U5925 ( .A1(MEM_stage_inst_dmem_ram_458), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n5794) );
NAND2_X1 MEM_stage_inst_dmem_U5924 ( .A1(MEM_stage_inst_dmem_n5792), .A2(MEM_stage_inst_dmem_n5791), .ZN(MEM_stage_inst_dmem_n5796) );
NAND2_X1 MEM_stage_inst_dmem_U5923 ( .A1(MEM_stage_inst_dmem_ram_90), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n5791) );
NAND2_X1 MEM_stage_inst_dmem_U5922 ( .A1(MEM_stage_inst_dmem_ram_794), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n5792) );
NOR2_X1 MEM_stage_inst_dmem_U5921 ( .A1(MEM_stage_inst_dmem_n5790), .A2(MEM_stage_inst_dmem_n5789), .ZN(MEM_stage_inst_dmem_n5798) );
NAND2_X1 MEM_stage_inst_dmem_U5920 ( .A1(MEM_stage_inst_dmem_n5788), .A2(MEM_stage_inst_dmem_n5787), .ZN(MEM_stage_inst_dmem_n5789) );
NAND2_X1 MEM_stage_inst_dmem_U5919 ( .A1(MEM_stage_inst_dmem_ram_58), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n5787) );
NAND2_X1 MEM_stage_inst_dmem_U5918 ( .A1(MEM_stage_inst_dmem_ram_10), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n5788) );
NAND2_X1 MEM_stage_inst_dmem_U5917 ( .A1(MEM_stage_inst_dmem_n5786), .A2(MEM_stage_inst_dmem_n5785), .ZN(MEM_stage_inst_dmem_n5790) );
NAND2_X1 MEM_stage_inst_dmem_U5916 ( .A1(MEM_stage_inst_dmem_ram_842), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n5785) );
NAND2_X1 MEM_stage_inst_dmem_U5915 ( .A1(MEM_stage_inst_dmem_ram_538), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n5786) );
NOR2_X1 MEM_stage_inst_dmem_U5914 ( .A1(MEM_stage_inst_dmem_n5784), .A2(MEM_stage_inst_dmem_n5783), .ZN(MEM_stage_inst_dmem_n5817) );
NAND2_X1 MEM_stage_inst_dmem_U5913 ( .A1(MEM_stage_inst_dmem_n5782), .A2(MEM_stage_inst_dmem_n5781), .ZN(MEM_stage_inst_dmem_n5783) );
NOR2_X1 MEM_stage_inst_dmem_U5912 ( .A1(MEM_stage_inst_dmem_n5780), .A2(MEM_stage_inst_dmem_n5779), .ZN(MEM_stage_inst_dmem_n5781) );
NAND2_X1 MEM_stage_inst_dmem_U5911 ( .A1(MEM_stage_inst_dmem_n5778), .A2(MEM_stage_inst_dmem_n5777), .ZN(MEM_stage_inst_dmem_n5779) );
NAND2_X1 MEM_stage_inst_dmem_U5910 ( .A1(MEM_stage_inst_dmem_ram_362), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n5777) );
NAND2_X1 MEM_stage_inst_dmem_U5909 ( .A1(MEM_stage_inst_dmem_ram_42), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n5778) );
NAND2_X1 MEM_stage_inst_dmem_U5908 ( .A1(MEM_stage_inst_dmem_n5776), .A2(MEM_stage_inst_dmem_n5775), .ZN(MEM_stage_inst_dmem_n5780) );
NAND2_X1 MEM_stage_inst_dmem_U5907 ( .A1(MEM_stage_inst_dmem_ram_394), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n5775) );
NAND2_X1 MEM_stage_inst_dmem_U5906 ( .A1(MEM_stage_inst_dmem_ram_938), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n5776) );
NOR2_X1 MEM_stage_inst_dmem_U5905 ( .A1(MEM_stage_inst_dmem_n5774), .A2(MEM_stage_inst_dmem_n5773), .ZN(MEM_stage_inst_dmem_n5782) );
NAND2_X1 MEM_stage_inst_dmem_U5904 ( .A1(MEM_stage_inst_dmem_n5772), .A2(MEM_stage_inst_dmem_n5771), .ZN(MEM_stage_inst_dmem_n5773) );
NAND2_X1 MEM_stage_inst_dmem_U5903 ( .A1(MEM_stage_inst_dmem_ram_874), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n5771) );
NAND2_X1 MEM_stage_inst_dmem_U5902 ( .A1(MEM_stage_inst_dmem_ram_250), .A2(MEM_stage_inst_dmem_n39), .ZN(MEM_stage_inst_dmem_n5772) );
NAND2_X1 MEM_stage_inst_dmem_U5901 ( .A1(MEM_stage_inst_dmem_n5770), .A2(MEM_stage_inst_dmem_n5769), .ZN(MEM_stage_inst_dmem_n5774) );
NAND2_X1 MEM_stage_inst_dmem_U5900 ( .A1(MEM_stage_inst_dmem_ram_314), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n5769) );
NAND2_X1 MEM_stage_inst_dmem_U5899 ( .A1(MEM_stage_inst_dmem_ram_986), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n5770) );
NAND2_X1 MEM_stage_inst_dmem_U5898 ( .A1(MEM_stage_inst_dmem_n5768), .A2(MEM_stage_inst_dmem_n5767), .ZN(MEM_stage_inst_dmem_n5784) );
NOR2_X1 MEM_stage_inst_dmem_U5897 ( .A1(MEM_stage_inst_dmem_n5766), .A2(MEM_stage_inst_dmem_n5765), .ZN(MEM_stage_inst_dmem_n5767) );
NAND2_X1 MEM_stage_inst_dmem_U5896 ( .A1(MEM_stage_inst_dmem_n5764), .A2(MEM_stage_inst_dmem_n5763), .ZN(MEM_stage_inst_dmem_n5765) );
NAND2_X1 MEM_stage_inst_dmem_U5895 ( .A1(MEM_stage_inst_dmem_ram_858), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n5763) );
NAND2_X1 MEM_stage_inst_dmem_U5894 ( .A1(MEM_stage_inst_dmem_ram_682), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n5764) );
NAND2_X1 MEM_stage_inst_dmem_U5893 ( .A1(MEM_stage_inst_dmem_n5762), .A2(MEM_stage_inst_dmem_n5761), .ZN(MEM_stage_inst_dmem_n5766) );
NAND2_X1 MEM_stage_inst_dmem_U5892 ( .A1(MEM_stage_inst_dmem_ram_506), .A2(MEM_stage_inst_dmem_n64), .ZN(MEM_stage_inst_dmem_n5761) );
NAND2_X1 MEM_stage_inst_dmem_U5891 ( .A1(MEM_stage_inst_dmem_ram_26), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n5762) );
NOR2_X1 MEM_stage_inst_dmem_U5890 ( .A1(MEM_stage_inst_dmem_n5760), .A2(MEM_stage_inst_dmem_n5759), .ZN(MEM_stage_inst_dmem_n5768) );
NAND2_X1 MEM_stage_inst_dmem_U5889 ( .A1(MEM_stage_inst_dmem_n5758), .A2(MEM_stage_inst_dmem_n5757), .ZN(MEM_stage_inst_dmem_n5759) );
NAND2_X1 MEM_stage_inst_dmem_U5888 ( .A1(MEM_stage_inst_dmem_ram_634), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n5757) );
NAND2_X1 MEM_stage_inst_dmem_U5887 ( .A1(MEM_stage_inst_dmem_ram_106), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n5758) );
NAND2_X1 MEM_stage_inst_dmem_U5886 ( .A1(MEM_stage_inst_dmem_n5756), .A2(MEM_stage_inst_dmem_n5755), .ZN(MEM_stage_inst_dmem_n5760) );
NAND2_X1 MEM_stage_inst_dmem_U5885 ( .A1(MEM_stage_inst_dmem_ram_522), .A2(MEM_stage_inst_dmem_n8225), .ZN(MEM_stage_inst_dmem_n5755) );
NAND2_X1 MEM_stage_inst_dmem_U5884 ( .A1(MEM_stage_inst_dmem_ram_730), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n5756) );
NAND2_X1 MEM_stage_inst_dmem_U5883 ( .A1(MEM_stage_inst_dmem_n5754), .A2(MEM_stage_inst_dmem_n5753), .ZN(MEM_stage_inst_dmem_n5819) );
NOR2_X1 MEM_stage_inst_dmem_U5882 ( .A1(MEM_stage_inst_dmem_n5752), .A2(MEM_stage_inst_dmem_n5751), .ZN(MEM_stage_inst_dmem_n5753) );
NAND2_X1 MEM_stage_inst_dmem_U5881 ( .A1(MEM_stage_inst_dmem_n5750), .A2(MEM_stage_inst_dmem_n5749), .ZN(MEM_stage_inst_dmem_n5751) );
NOR2_X1 MEM_stage_inst_dmem_U5880 ( .A1(MEM_stage_inst_dmem_n5748), .A2(MEM_stage_inst_dmem_n5747), .ZN(MEM_stage_inst_dmem_n5749) );
NAND2_X1 MEM_stage_inst_dmem_U5879 ( .A1(MEM_stage_inst_dmem_n5746), .A2(MEM_stage_inst_dmem_n5745), .ZN(MEM_stage_inst_dmem_n5747) );
NAND2_X1 MEM_stage_inst_dmem_U5878 ( .A1(MEM_stage_inst_dmem_ram_570), .A2(MEM_stage_inst_dmem_n8169), .ZN(MEM_stage_inst_dmem_n5745) );
NAND2_X1 MEM_stage_inst_dmem_U5877 ( .A1(MEM_stage_inst_dmem_ram_346), .A2(MEM_stage_inst_dmem_n3216), .ZN(MEM_stage_inst_dmem_n5746) );
NAND2_X1 MEM_stage_inst_dmem_U5876 ( .A1(MEM_stage_inst_dmem_n5744), .A2(MEM_stage_inst_dmem_n5743), .ZN(MEM_stage_inst_dmem_n5748) );
NAND2_X1 MEM_stage_inst_dmem_U5875 ( .A1(MEM_stage_inst_dmem_ram_922), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n5743) );
NAND2_X1 MEM_stage_inst_dmem_U5874 ( .A1(MEM_stage_inst_dmem_ram_970), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n5744) );
NOR2_X1 MEM_stage_inst_dmem_U5873 ( .A1(MEM_stage_inst_dmem_n5742), .A2(MEM_stage_inst_dmem_n5741), .ZN(MEM_stage_inst_dmem_n5750) );
NAND2_X1 MEM_stage_inst_dmem_U5872 ( .A1(MEM_stage_inst_dmem_n5740), .A2(MEM_stage_inst_dmem_n5739), .ZN(MEM_stage_inst_dmem_n5741) );
NAND2_X1 MEM_stage_inst_dmem_U5871 ( .A1(MEM_stage_inst_dmem_ram_138), .A2(MEM_stage_inst_dmem_n8174), .ZN(MEM_stage_inst_dmem_n5739) );
NAND2_X1 MEM_stage_inst_dmem_U5870 ( .A1(MEM_stage_inst_dmem_ram_586), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n5740) );
NAND2_X1 MEM_stage_inst_dmem_U5869 ( .A1(MEM_stage_inst_dmem_n5738), .A2(MEM_stage_inst_dmem_n5737), .ZN(MEM_stage_inst_dmem_n5742) );
NAND2_X1 MEM_stage_inst_dmem_U5868 ( .A1(MEM_stage_inst_dmem_ram_1002), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n5737) );
NAND2_X1 MEM_stage_inst_dmem_U5867 ( .A1(MEM_stage_inst_dmem_ram_602), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n5738) );
NAND2_X1 MEM_stage_inst_dmem_U5866 ( .A1(MEM_stage_inst_dmem_n5736), .A2(MEM_stage_inst_dmem_n5735), .ZN(MEM_stage_inst_dmem_n5752) );
NOR2_X1 MEM_stage_inst_dmem_U5865 ( .A1(MEM_stage_inst_dmem_n5734), .A2(MEM_stage_inst_dmem_n5733), .ZN(MEM_stage_inst_dmem_n5735) );
NAND2_X1 MEM_stage_inst_dmem_U5864 ( .A1(MEM_stage_inst_dmem_n5732), .A2(MEM_stage_inst_dmem_n5731), .ZN(MEM_stage_inst_dmem_n5733) );
NAND2_X1 MEM_stage_inst_dmem_U5863 ( .A1(MEM_stage_inst_dmem_ram_714), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n5731) );
NAND2_X1 MEM_stage_inst_dmem_U5862 ( .A1(MEM_stage_inst_dmem_ram_698), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n5732) );
NAND2_X1 MEM_stage_inst_dmem_U5861 ( .A1(MEM_stage_inst_dmem_n5730), .A2(MEM_stage_inst_dmem_n5729), .ZN(MEM_stage_inst_dmem_n5734) );
NAND2_X1 MEM_stage_inst_dmem_U5860 ( .A1(MEM_stage_inst_dmem_ram_202), .A2(MEM_stage_inst_dmem_n8256), .ZN(MEM_stage_inst_dmem_n5729) );
NAND2_X1 MEM_stage_inst_dmem_U5859 ( .A1(MEM_stage_inst_dmem_ram_778), .A2(MEM_stage_inst_dmem_n37), .ZN(MEM_stage_inst_dmem_n5730) );
NOR2_X1 MEM_stage_inst_dmem_U5858 ( .A1(MEM_stage_inst_dmem_n5728), .A2(MEM_stage_inst_dmem_n5727), .ZN(MEM_stage_inst_dmem_n5736) );
NAND2_X1 MEM_stage_inst_dmem_U5857 ( .A1(MEM_stage_inst_dmem_n5726), .A2(MEM_stage_inst_dmem_n5725), .ZN(MEM_stage_inst_dmem_n5727) );
NAND2_X1 MEM_stage_inst_dmem_U5856 ( .A1(MEM_stage_inst_dmem_ram_410), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n5725) );
NAND2_X1 MEM_stage_inst_dmem_U5855 ( .A1(MEM_stage_inst_dmem_ram_426), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n5726) );
NAND2_X1 MEM_stage_inst_dmem_U5854 ( .A1(MEM_stage_inst_dmem_n5724), .A2(MEM_stage_inst_dmem_n5723), .ZN(MEM_stage_inst_dmem_n5728) );
NAND2_X1 MEM_stage_inst_dmem_U5853 ( .A1(MEM_stage_inst_dmem_ram_554), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n5723) );
NAND2_X1 MEM_stage_inst_dmem_U5852 ( .A1(MEM_stage_inst_dmem_ram_826), .A2(MEM_stage_inst_dmem_n46), .ZN(MEM_stage_inst_dmem_n5724) );
NOR2_X1 MEM_stage_inst_dmem_U5851 ( .A1(MEM_stage_inst_dmem_n5722), .A2(MEM_stage_inst_dmem_n5721), .ZN(MEM_stage_inst_dmem_n5754) );
NAND2_X1 MEM_stage_inst_dmem_U5850 ( .A1(MEM_stage_inst_dmem_n5720), .A2(MEM_stage_inst_dmem_n5719), .ZN(MEM_stage_inst_dmem_n5721) );
NOR2_X1 MEM_stage_inst_dmem_U5849 ( .A1(MEM_stage_inst_dmem_n5718), .A2(MEM_stage_inst_dmem_n5717), .ZN(MEM_stage_inst_dmem_n5719) );
NAND2_X1 MEM_stage_inst_dmem_U5848 ( .A1(MEM_stage_inst_dmem_n5716), .A2(MEM_stage_inst_dmem_n5715), .ZN(MEM_stage_inst_dmem_n5717) );
NAND2_X1 MEM_stage_inst_dmem_U5847 ( .A1(MEM_stage_inst_dmem_ram_122), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n5715) );
NAND2_X1 MEM_stage_inst_dmem_U5846 ( .A1(MEM_stage_inst_dmem_ram_746), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n5716) );
NAND2_X1 MEM_stage_inst_dmem_U5845 ( .A1(MEM_stage_inst_dmem_n5714), .A2(MEM_stage_inst_dmem_n5713), .ZN(MEM_stage_inst_dmem_n5718) );
NAND2_X1 MEM_stage_inst_dmem_U5844 ( .A1(MEM_stage_inst_dmem_ram_650), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n5713) );
NAND2_X1 MEM_stage_inst_dmem_U5843 ( .A1(MEM_stage_inst_dmem_ram_170), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n5714) );
NOR2_X1 MEM_stage_inst_dmem_U5842 ( .A1(MEM_stage_inst_dmem_n5712), .A2(MEM_stage_inst_dmem_n5711), .ZN(MEM_stage_inst_dmem_n5720) );
NAND2_X1 MEM_stage_inst_dmem_U5841 ( .A1(MEM_stage_inst_dmem_n5710), .A2(MEM_stage_inst_dmem_n5709), .ZN(MEM_stage_inst_dmem_n5711) );
NAND2_X1 MEM_stage_inst_dmem_U5840 ( .A1(MEM_stage_inst_dmem_ram_954), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n5709) );
NAND2_X1 MEM_stage_inst_dmem_U5839 ( .A1(MEM_stage_inst_dmem_ram_810), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n5710) );
NAND2_X1 MEM_stage_inst_dmem_U5838 ( .A1(MEM_stage_inst_dmem_n5708), .A2(MEM_stage_inst_dmem_n5707), .ZN(MEM_stage_inst_dmem_n5712) );
NAND2_X1 MEM_stage_inst_dmem_U5837 ( .A1(MEM_stage_inst_dmem_ram_282), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n5707) );
NAND2_X1 MEM_stage_inst_dmem_U5836 ( .A1(MEM_stage_inst_dmem_ram_218), .A2(MEM_stage_inst_dmem_n8206), .ZN(MEM_stage_inst_dmem_n5708) );
NAND2_X1 MEM_stage_inst_dmem_U5835 ( .A1(MEM_stage_inst_dmem_n5706), .A2(MEM_stage_inst_dmem_n5705), .ZN(MEM_stage_inst_dmem_n5722) );
NOR2_X1 MEM_stage_inst_dmem_U5834 ( .A1(MEM_stage_inst_dmem_n5704), .A2(MEM_stage_inst_dmem_n5703), .ZN(MEM_stage_inst_dmem_n5705) );
NAND2_X1 MEM_stage_inst_dmem_U5833 ( .A1(MEM_stage_inst_dmem_n5702), .A2(MEM_stage_inst_dmem_n5701), .ZN(MEM_stage_inst_dmem_n5703) );
NAND2_X1 MEM_stage_inst_dmem_U5832 ( .A1(MEM_stage_inst_dmem_ram_490), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n5701) );
NAND2_X1 MEM_stage_inst_dmem_U5831 ( .A1(MEM_stage_inst_dmem_ram_906), .A2(MEM_stage_inst_dmem_n8193), .ZN(MEM_stage_inst_dmem_n5702) );
NAND2_X1 MEM_stage_inst_dmem_U5830 ( .A1(MEM_stage_inst_dmem_n5700), .A2(MEM_stage_inst_dmem_n5699), .ZN(MEM_stage_inst_dmem_n5704) );
NAND2_X1 MEM_stage_inst_dmem_U5829 ( .A1(MEM_stage_inst_dmem_ram_618), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n5699) );
NAND2_X1 MEM_stage_inst_dmem_U5828 ( .A1(MEM_stage_inst_dmem_ram_298), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n5700) );
NOR2_X1 MEM_stage_inst_dmem_U5827 ( .A1(MEM_stage_inst_dmem_n5698), .A2(MEM_stage_inst_dmem_n5697), .ZN(MEM_stage_inst_dmem_n5706) );
NAND2_X1 MEM_stage_inst_dmem_U5826 ( .A1(MEM_stage_inst_dmem_n5696), .A2(MEM_stage_inst_dmem_n5695), .ZN(MEM_stage_inst_dmem_n5697) );
NAND2_X1 MEM_stage_inst_dmem_U5825 ( .A1(MEM_stage_inst_dmem_ram_442), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n5695) );
NAND2_X1 MEM_stage_inst_dmem_U5824 ( .A1(MEM_stage_inst_dmem_ram_74), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n5696) );
NAND2_X1 MEM_stage_inst_dmem_U5823 ( .A1(MEM_stage_inst_dmem_n5694), .A2(MEM_stage_inst_dmem_n5693), .ZN(MEM_stage_inst_dmem_n5698) );
NAND2_X1 MEM_stage_inst_dmem_U5822 ( .A1(MEM_stage_inst_dmem_ram_890), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n5693) );
NAND2_X1 MEM_stage_inst_dmem_U5821 ( .A1(MEM_stage_inst_dmem_ram_330), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n5694) );
NOR2_X1 MEM_stage_inst_dmem_U5820 ( .A1(MEM_stage_inst_dmem_n5692), .A2(MEM_stage_inst_dmem_n5691), .ZN(MEM_stage_inst_dmem_n5952) );
NOR2_X1 MEM_stage_inst_dmem_U5819 ( .A1(MEM_stage_inst_dmem_n5690), .A2(MEM_stage_inst_dmem_n8286), .ZN(MEM_stage_inst_dmem_n5691) );
NOR2_X1 MEM_stage_inst_dmem_U5818 ( .A1(MEM_stage_inst_dmem_n5689), .A2(MEM_stage_inst_dmem_n5688), .ZN(MEM_stage_inst_dmem_n5690) );
NAND2_X1 MEM_stage_inst_dmem_U5817 ( .A1(MEM_stage_inst_dmem_n5687), .A2(MEM_stage_inst_dmem_n5686), .ZN(MEM_stage_inst_dmem_n5688) );
NOR2_X1 MEM_stage_inst_dmem_U5816 ( .A1(MEM_stage_inst_dmem_n5685), .A2(MEM_stage_inst_dmem_n5684), .ZN(MEM_stage_inst_dmem_n5686) );
NAND2_X1 MEM_stage_inst_dmem_U5815 ( .A1(MEM_stage_inst_dmem_n5683), .A2(MEM_stage_inst_dmem_n5682), .ZN(MEM_stage_inst_dmem_n5684) );
NOR2_X1 MEM_stage_inst_dmem_U5814 ( .A1(MEM_stage_inst_dmem_n5681), .A2(MEM_stage_inst_dmem_n5680), .ZN(MEM_stage_inst_dmem_n5682) );
NAND2_X1 MEM_stage_inst_dmem_U5813 ( .A1(MEM_stage_inst_dmem_n5679), .A2(MEM_stage_inst_dmem_n5678), .ZN(MEM_stage_inst_dmem_n5680) );
NAND2_X1 MEM_stage_inst_dmem_U5812 ( .A1(MEM_stage_inst_dmem_ram_2746), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n5678) );
NAND2_X1 MEM_stage_inst_dmem_U5811 ( .A1(MEM_stage_inst_dmem_ram_2986), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n5679) );
NAND2_X1 MEM_stage_inst_dmem_U5810 ( .A1(MEM_stage_inst_dmem_n5677), .A2(MEM_stage_inst_dmem_n5676), .ZN(MEM_stage_inst_dmem_n5681) );
NAND2_X1 MEM_stage_inst_dmem_U5809 ( .A1(MEM_stage_inst_dmem_ram_2938), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n5676) );
NAND2_X1 MEM_stage_inst_dmem_U5808 ( .A1(MEM_stage_inst_dmem_ram_2970), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n5677) );
NOR2_X1 MEM_stage_inst_dmem_U5807 ( .A1(MEM_stage_inst_dmem_n5675), .A2(MEM_stage_inst_dmem_n5674), .ZN(MEM_stage_inst_dmem_n5683) );
NAND2_X1 MEM_stage_inst_dmem_U5806 ( .A1(MEM_stage_inst_dmem_n5673), .A2(MEM_stage_inst_dmem_n5672), .ZN(MEM_stage_inst_dmem_n5674) );
NAND2_X1 MEM_stage_inst_dmem_U5805 ( .A1(MEM_stage_inst_dmem_ram_3034), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n5672) );
NAND2_X1 MEM_stage_inst_dmem_U5804 ( .A1(MEM_stage_inst_dmem_ram_2346), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n5673) );
NAND2_X1 MEM_stage_inst_dmem_U5803 ( .A1(MEM_stage_inst_dmem_n5671), .A2(MEM_stage_inst_dmem_n5670), .ZN(MEM_stage_inst_dmem_n5675) );
NAND2_X1 MEM_stage_inst_dmem_U5802 ( .A1(MEM_stage_inst_dmem_ram_2282), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n5670) );
NAND2_X1 MEM_stage_inst_dmem_U5801 ( .A1(MEM_stage_inst_dmem_ram_2330), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n5671) );
NAND2_X1 MEM_stage_inst_dmem_U5800 ( .A1(MEM_stage_inst_dmem_n5669), .A2(MEM_stage_inst_dmem_n5668), .ZN(MEM_stage_inst_dmem_n5685) );
NOR2_X1 MEM_stage_inst_dmem_U5799 ( .A1(MEM_stage_inst_dmem_n5667), .A2(MEM_stage_inst_dmem_n5666), .ZN(MEM_stage_inst_dmem_n5668) );
NAND2_X1 MEM_stage_inst_dmem_U5798 ( .A1(MEM_stage_inst_dmem_n5665), .A2(MEM_stage_inst_dmem_n5664), .ZN(MEM_stage_inst_dmem_n5666) );
NAND2_X1 MEM_stage_inst_dmem_U5797 ( .A1(MEM_stage_inst_dmem_ram_2410), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n5664) );
NAND2_X1 MEM_stage_inst_dmem_U5796 ( .A1(MEM_stage_inst_dmem_ram_2714), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n5665) );
NAND2_X1 MEM_stage_inst_dmem_U5795 ( .A1(MEM_stage_inst_dmem_n5663), .A2(MEM_stage_inst_dmem_n5662), .ZN(MEM_stage_inst_dmem_n5667) );
NAND2_X1 MEM_stage_inst_dmem_U5794 ( .A1(MEM_stage_inst_dmem_ram_2826), .A2(MEM_stage_inst_dmem_n8472), .ZN(MEM_stage_inst_dmem_n5662) );
NAND2_X1 MEM_stage_inst_dmem_U5793 ( .A1(MEM_stage_inst_dmem_ram_2890), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n5663) );
NOR2_X1 MEM_stage_inst_dmem_U5792 ( .A1(MEM_stage_inst_dmem_n5661), .A2(MEM_stage_inst_dmem_n5660), .ZN(MEM_stage_inst_dmem_n5669) );
NAND2_X1 MEM_stage_inst_dmem_U5791 ( .A1(MEM_stage_inst_dmem_n5659), .A2(MEM_stage_inst_dmem_n5658), .ZN(MEM_stage_inst_dmem_n5660) );
NAND2_X1 MEM_stage_inst_dmem_U5790 ( .A1(MEM_stage_inst_dmem_ram_2074), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n5658) );
NAND2_X1 MEM_stage_inst_dmem_U5789 ( .A1(MEM_stage_inst_dmem_ram_2314), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n5659) );
NAND2_X1 MEM_stage_inst_dmem_U5788 ( .A1(MEM_stage_inst_dmem_n5657), .A2(MEM_stage_inst_dmem_n5656), .ZN(MEM_stage_inst_dmem_n5661) );
NAND2_X1 MEM_stage_inst_dmem_U5787 ( .A1(MEM_stage_inst_dmem_ram_2730), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n5656) );
NAND2_X1 MEM_stage_inst_dmem_U5786 ( .A1(MEM_stage_inst_dmem_ram_2586), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n5657) );
NOR2_X1 MEM_stage_inst_dmem_U5785 ( .A1(MEM_stage_inst_dmem_n5655), .A2(MEM_stage_inst_dmem_n5654), .ZN(MEM_stage_inst_dmem_n5687) );
NAND2_X1 MEM_stage_inst_dmem_U5784 ( .A1(MEM_stage_inst_dmem_n5653), .A2(MEM_stage_inst_dmem_n5652), .ZN(MEM_stage_inst_dmem_n5654) );
NOR2_X1 MEM_stage_inst_dmem_U5783 ( .A1(MEM_stage_inst_dmem_n5651), .A2(MEM_stage_inst_dmem_n5650), .ZN(MEM_stage_inst_dmem_n5652) );
NAND2_X1 MEM_stage_inst_dmem_U5782 ( .A1(MEM_stage_inst_dmem_n5649), .A2(MEM_stage_inst_dmem_n5648), .ZN(MEM_stage_inst_dmem_n5650) );
NAND2_X1 MEM_stage_inst_dmem_U5781 ( .A1(MEM_stage_inst_dmem_ram_2666), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n5648) );
NAND2_X1 MEM_stage_inst_dmem_U5780 ( .A1(MEM_stage_inst_dmem_ram_2794), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n5649) );
NAND2_X1 MEM_stage_inst_dmem_U5779 ( .A1(MEM_stage_inst_dmem_n5647), .A2(MEM_stage_inst_dmem_n5646), .ZN(MEM_stage_inst_dmem_n5651) );
NAND2_X1 MEM_stage_inst_dmem_U5778 ( .A1(MEM_stage_inst_dmem_ram_2554), .A2(MEM_stage_inst_dmem_n64), .ZN(MEM_stage_inst_dmem_n5646) );
NAND2_X1 MEM_stage_inst_dmem_U5777 ( .A1(MEM_stage_inst_dmem_ram_3066), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n5647) );
NOR2_X1 MEM_stage_inst_dmem_U5776 ( .A1(MEM_stage_inst_dmem_n5645), .A2(MEM_stage_inst_dmem_n5644), .ZN(MEM_stage_inst_dmem_n5653) );
NAND2_X1 MEM_stage_inst_dmem_U5775 ( .A1(MEM_stage_inst_dmem_n5643), .A2(MEM_stage_inst_dmem_n5642), .ZN(MEM_stage_inst_dmem_n5644) );
NAND2_X1 MEM_stage_inst_dmem_U5774 ( .A1(MEM_stage_inst_dmem_ram_2522), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n5642) );
NAND2_X1 MEM_stage_inst_dmem_U5773 ( .A1(MEM_stage_inst_dmem_ram_2650), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n5643) );
NAND2_X1 MEM_stage_inst_dmem_U5772 ( .A1(MEM_stage_inst_dmem_n5641), .A2(MEM_stage_inst_dmem_n5640), .ZN(MEM_stage_inst_dmem_n5645) );
NAND2_X1 MEM_stage_inst_dmem_U5771 ( .A1(MEM_stage_inst_dmem_ram_2618), .A2(MEM_stage_inst_dmem_n8169), .ZN(MEM_stage_inst_dmem_n5640) );
NAND2_X1 MEM_stage_inst_dmem_U5770 ( .A1(MEM_stage_inst_dmem_ram_2762), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n5641) );
NAND2_X1 MEM_stage_inst_dmem_U5769 ( .A1(MEM_stage_inst_dmem_n5639), .A2(MEM_stage_inst_dmem_n5638), .ZN(MEM_stage_inst_dmem_n5655) );
NOR2_X1 MEM_stage_inst_dmem_U5768 ( .A1(MEM_stage_inst_dmem_n5637), .A2(MEM_stage_inst_dmem_n5636), .ZN(MEM_stage_inst_dmem_n5638) );
NAND2_X1 MEM_stage_inst_dmem_U5767 ( .A1(MEM_stage_inst_dmem_n5635), .A2(MEM_stage_inst_dmem_n5634), .ZN(MEM_stage_inst_dmem_n5636) );
NAND2_X1 MEM_stage_inst_dmem_U5766 ( .A1(MEM_stage_inst_dmem_ram_3050), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n5634) );
NAND2_X1 MEM_stage_inst_dmem_U5765 ( .A1(MEM_stage_inst_dmem_ram_2602), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n5635) );
NAND2_X1 MEM_stage_inst_dmem_U5764 ( .A1(MEM_stage_inst_dmem_n5633), .A2(MEM_stage_inst_dmem_n5632), .ZN(MEM_stage_inst_dmem_n5637) );
NAND2_X1 MEM_stage_inst_dmem_U5763 ( .A1(MEM_stage_inst_dmem_ram_2106), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n5632) );
NAND2_X1 MEM_stage_inst_dmem_U5762 ( .A1(MEM_stage_inst_dmem_ram_2810), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n5633) );
NOR2_X1 MEM_stage_inst_dmem_U5761 ( .A1(MEM_stage_inst_dmem_n5631), .A2(MEM_stage_inst_dmem_n5630), .ZN(MEM_stage_inst_dmem_n5639) );
NAND2_X1 MEM_stage_inst_dmem_U5760 ( .A1(MEM_stage_inst_dmem_n5629), .A2(MEM_stage_inst_dmem_n5628), .ZN(MEM_stage_inst_dmem_n5630) );
NAND2_X1 MEM_stage_inst_dmem_U5759 ( .A1(MEM_stage_inst_dmem_ram_2538), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n5628) );
NAND2_X1 MEM_stage_inst_dmem_U5758 ( .A1(MEM_stage_inst_dmem_ram_2202), .A2(MEM_stage_inst_dmem_n44), .ZN(MEM_stage_inst_dmem_n5629) );
NAND2_X1 MEM_stage_inst_dmem_U5757 ( .A1(MEM_stage_inst_dmem_n5627), .A2(MEM_stage_inst_dmem_n5626), .ZN(MEM_stage_inst_dmem_n5631) );
NAND2_X1 MEM_stage_inst_dmem_U5756 ( .A1(MEM_stage_inst_dmem_ram_2682), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n5626) );
NAND2_X1 MEM_stage_inst_dmem_U5755 ( .A1(MEM_stage_inst_dmem_ram_2154), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n5627) );
NAND2_X1 MEM_stage_inst_dmem_U5754 ( .A1(MEM_stage_inst_dmem_n5625), .A2(MEM_stage_inst_dmem_n5624), .ZN(MEM_stage_inst_dmem_n5689) );
NOR2_X1 MEM_stage_inst_dmem_U5753 ( .A1(MEM_stage_inst_dmem_n5623), .A2(MEM_stage_inst_dmem_n5622), .ZN(MEM_stage_inst_dmem_n5624) );
NAND2_X1 MEM_stage_inst_dmem_U5752 ( .A1(MEM_stage_inst_dmem_n5621), .A2(MEM_stage_inst_dmem_n5620), .ZN(MEM_stage_inst_dmem_n5622) );
NOR2_X1 MEM_stage_inst_dmem_U5751 ( .A1(MEM_stage_inst_dmem_n5619), .A2(MEM_stage_inst_dmem_n5618), .ZN(MEM_stage_inst_dmem_n5620) );
NAND2_X1 MEM_stage_inst_dmem_U5750 ( .A1(MEM_stage_inst_dmem_n5617), .A2(MEM_stage_inst_dmem_n5616), .ZN(MEM_stage_inst_dmem_n5618) );
NAND2_X1 MEM_stage_inst_dmem_U5749 ( .A1(MEM_stage_inst_dmem_ram_2122), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n5616) );
NAND2_X1 MEM_stage_inst_dmem_U5748 ( .A1(MEM_stage_inst_dmem_ram_2186), .A2(MEM_stage_inst_dmem_n8174), .ZN(MEM_stage_inst_dmem_n5617) );
NAND2_X1 MEM_stage_inst_dmem_U5747 ( .A1(MEM_stage_inst_dmem_n5615), .A2(MEM_stage_inst_dmem_n5614), .ZN(MEM_stage_inst_dmem_n5619) );
NAND2_X1 MEM_stage_inst_dmem_U5746 ( .A1(MEM_stage_inst_dmem_ram_2378), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n5614) );
NAND2_X1 MEM_stage_inst_dmem_U5745 ( .A1(MEM_stage_inst_dmem_ram_2458), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n5615) );
NOR2_X1 MEM_stage_inst_dmem_U5744 ( .A1(MEM_stage_inst_dmem_n5613), .A2(MEM_stage_inst_dmem_n5612), .ZN(MEM_stage_inst_dmem_n5621) );
NAND2_X1 MEM_stage_inst_dmem_U5743 ( .A1(MEM_stage_inst_dmem_n5611), .A2(MEM_stage_inst_dmem_n5610), .ZN(MEM_stage_inst_dmem_n5612) );
NAND2_X1 MEM_stage_inst_dmem_U5742 ( .A1(MEM_stage_inst_dmem_ram_2170), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n5610) );
NAND2_X1 MEM_stage_inst_dmem_U5741 ( .A1(MEM_stage_inst_dmem_ram_2778), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n5611) );
NAND2_X1 MEM_stage_inst_dmem_U5740 ( .A1(MEM_stage_inst_dmem_n5609), .A2(MEM_stage_inst_dmem_n5608), .ZN(MEM_stage_inst_dmem_n5613) );
NAND2_X1 MEM_stage_inst_dmem_U5739 ( .A1(MEM_stage_inst_dmem_ram_3002), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n5608) );
NAND2_X1 MEM_stage_inst_dmem_U5738 ( .A1(MEM_stage_inst_dmem_ram_2394), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n5609) );
NAND2_X1 MEM_stage_inst_dmem_U5737 ( .A1(MEM_stage_inst_dmem_n5607), .A2(MEM_stage_inst_dmem_n5606), .ZN(MEM_stage_inst_dmem_n5623) );
NOR2_X1 MEM_stage_inst_dmem_U5736 ( .A1(MEM_stage_inst_dmem_n5605), .A2(MEM_stage_inst_dmem_n5604), .ZN(MEM_stage_inst_dmem_n5606) );
NAND2_X1 MEM_stage_inst_dmem_U5735 ( .A1(MEM_stage_inst_dmem_n5603), .A2(MEM_stage_inst_dmem_n5602), .ZN(MEM_stage_inst_dmem_n5604) );
NAND2_X1 MEM_stage_inst_dmem_U5734 ( .A1(MEM_stage_inst_dmem_ram_2906), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n5602) );
NAND2_X1 MEM_stage_inst_dmem_U5733 ( .A1(MEM_stage_inst_dmem_ram_2298), .A2(MEM_stage_inst_dmem_n39), .ZN(MEM_stage_inst_dmem_n5603) );
NAND2_X1 MEM_stage_inst_dmem_U5732 ( .A1(MEM_stage_inst_dmem_n5601), .A2(MEM_stage_inst_dmem_n5600), .ZN(MEM_stage_inst_dmem_n5605) );
NAND2_X1 MEM_stage_inst_dmem_U5731 ( .A1(MEM_stage_inst_dmem_ram_2138), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n5600) );
NAND2_X1 MEM_stage_inst_dmem_U5730 ( .A1(MEM_stage_inst_dmem_ram_2842), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n5601) );
NOR2_X1 MEM_stage_inst_dmem_U5729 ( .A1(MEM_stage_inst_dmem_n5599), .A2(MEM_stage_inst_dmem_n5598), .ZN(MEM_stage_inst_dmem_n5607) );
NAND2_X1 MEM_stage_inst_dmem_U5728 ( .A1(MEM_stage_inst_dmem_n5597), .A2(MEM_stage_inst_dmem_n5596), .ZN(MEM_stage_inst_dmem_n5598) );
NAND2_X1 MEM_stage_inst_dmem_U5727 ( .A1(MEM_stage_inst_dmem_ram_2570), .A2(MEM_stage_inst_dmem_n8225), .ZN(MEM_stage_inst_dmem_n5596) );
NAND2_X1 MEM_stage_inst_dmem_U5726 ( .A1(MEM_stage_inst_dmem_ram_2058), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n5597) );
NAND2_X1 MEM_stage_inst_dmem_U5725 ( .A1(MEM_stage_inst_dmem_n5595), .A2(MEM_stage_inst_dmem_n5594), .ZN(MEM_stage_inst_dmem_n5599) );
NAND2_X1 MEM_stage_inst_dmem_U5724 ( .A1(MEM_stage_inst_dmem_ram_2858), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n5594) );
NAND2_X1 MEM_stage_inst_dmem_U5723 ( .A1(MEM_stage_inst_dmem_ram_2426), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n5595) );
NOR2_X1 MEM_stage_inst_dmem_U5722 ( .A1(MEM_stage_inst_dmem_n5593), .A2(MEM_stage_inst_dmem_n5592), .ZN(MEM_stage_inst_dmem_n5625) );
NAND2_X1 MEM_stage_inst_dmem_U5721 ( .A1(MEM_stage_inst_dmem_n5591), .A2(MEM_stage_inst_dmem_n5590), .ZN(MEM_stage_inst_dmem_n5592) );
NOR2_X1 MEM_stage_inst_dmem_U5720 ( .A1(MEM_stage_inst_dmem_n5589), .A2(MEM_stage_inst_dmem_n5588), .ZN(MEM_stage_inst_dmem_n5590) );
NAND2_X1 MEM_stage_inst_dmem_U5719 ( .A1(MEM_stage_inst_dmem_n5587), .A2(MEM_stage_inst_dmem_n5586), .ZN(MEM_stage_inst_dmem_n5588) );
NAND2_X1 MEM_stage_inst_dmem_U5718 ( .A1(MEM_stage_inst_dmem_ram_2954), .A2(MEM_stage_inst_dmem_n8193), .ZN(MEM_stage_inst_dmem_n5586) );
NAND2_X1 MEM_stage_inst_dmem_U5717 ( .A1(MEM_stage_inst_dmem_ram_2506), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n5587) );
NAND2_X1 MEM_stage_inst_dmem_U5716 ( .A1(MEM_stage_inst_dmem_n5585), .A2(MEM_stage_inst_dmem_n5584), .ZN(MEM_stage_inst_dmem_n5589) );
NAND2_X1 MEM_stage_inst_dmem_U5715 ( .A1(MEM_stage_inst_dmem_ram_3018), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n5584) );
NAND2_X1 MEM_stage_inst_dmem_U5714 ( .A1(MEM_stage_inst_dmem_ram_2474), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n5585) );
NOR2_X1 MEM_stage_inst_dmem_U5713 ( .A1(MEM_stage_inst_dmem_n5583), .A2(MEM_stage_inst_dmem_n5582), .ZN(MEM_stage_inst_dmem_n5591) );
NAND2_X1 MEM_stage_inst_dmem_U5712 ( .A1(MEM_stage_inst_dmem_n5581), .A2(MEM_stage_inst_dmem_n5580), .ZN(MEM_stage_inst_dmem_n5582) );
NAND2_X1 MEM_stage_inst_dmem_U5711 ( .A1(MEM_stage_inst_dmem_ram_2362), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n5580) );
NAND2_X1 MEM_stage_inst_dmem_U5710 ( .A1(MEM_stage_inst_dmem_ram_2634), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n5581) );
NAND2_X1 MEM_stage_inst_dmem_U5709 ( .A1(MEM_stage_inst_dmem_n5579), .A2(MEM_stage_inst_dmem_n5578), .ZN(MEM_stage_inst_dmem_n5583) );
NAND2_X1 MEM_stage_inst_dmem_U5708 ( .A1(MEM_stage_inst_dmem_ram_2922), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n5578) );
NAND2_X1 MEM_stage_inst_dmem_U5707 ( .A1(MEM_stage_inst_dmem_ram_2490), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n5579) );
NAND2_X1 MEM_stage_inst_dmem_U5706 ( .A1(MEM_stage_inst_dmem_n5577), .A2(MEM_stage_inst_dmem_n5576), .ZN(MEM_stage_inst_dmem_n5593) );
NOR2_X1 MEM_stage_inst_dmem_U5705 ( .A1(MEM_stage_inst_dmem_n5575), .A2(MEM_stage_inst_dmem_n5574), .ZN(MEM_stage_inst_dmem_n5576) );
NAND2_X1 MEM_stage_inst_dmem_U5704 ( .A1(MEM_stage_inst_dmem_n5573), .A2(MEM_stage_inst_dmem_n5572), .ZN(MEM_stage_inst_dmem_n5574) );
NAND2_X1 MEM_stage_inst_dmem_U5703 ( .A1(MEM_stage_inst_dmem_ram_2090), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n5572) );
NAND2_X1 MEM_stage_inst_dmem_U5702 ( .A1(MEM_stage_inst_dmem_ram_2442), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n5573) );
NAND2_X1 MEM_stage_inst_dmem_U5701 ( .A1(MEM_stage_inst_dmem_n5571), .A2(MEM_stage_inst_dmem_n5570), .ZN(MEM_stage_inst_dmem_n5575) );
NAND2_X1 MEM_stage_inst_dmem_U5700 ( .A1(MEM_stage_inst_dmem_ram_2250), .A2(MEM_stage_inst_dmem_n8256), .ZN(MEM_stage_inst_dmem_n5570) );
NAND2_X1 MEM_stage_inst_dmem_U5699 ( .A1(MEM_stage_inst_dmem_ram_2234), .A2(MEM_stage_inst_dmem_n8434), .ZN(MEM_stage_inst_dmem_n5571) );
NOR2_X1 MEM_stage_inst_dmem_U5698 ( .A1(MEM_stage_inst_dmem_n5569), .A2(MEM_stage_inst_dmem_n5568), .ZN(MEM_stage_inst_dmem_n5577) );
NAND2_X1 MEM_stage_inst_dmem_U5697 ( .A1(MEM_stage_inst_dmem_n5567), .A2(MEM_stage_inst_dmem_n5566), .ZN(MEM_stage_inst_dmem_n5568) );
NAND2_X1 MEM_stage_inst_dmem_U5696 ( .A1(MEM_stage_inst_dmem_ram_2874), .A2(MEM_stage_inst_dmem_n46), .ZN(MEM_stage_inst_dmem_n5566) );
NAND2_X1 MEM_stage_inst_dmem_U5695 ( .A1(MEM_stage_inst_dmem_ram_2266), .A2(MEM_stage_inst_dmem_n8206), .ZN(MEM_stage_inst_dmem_n5567) );
NAND2_X1 MEM_stage_inst_dmem_U5694 ( .A1(MEM_stage_inst_dmem_n5565), .A2(MEM_stage_inst_dmem_n5564), .ZN(MEM_stage_inst_dmem_n5569) );
NAND2_X1 MEM_stage_inst_dmem_U5693 ( .A1(MEM_stage_inst_dmem_ram_2698), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n5564) );
NAND2_X1 MEM_stage_inst_dmem_U5692 ( .A1(MEM_stage_inst_dmem_ram_2218), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n5565) );
NOR2_X1 MEM_stage_inst_dmem_U5691 ( .A1(MEM_stage_inst_dmem_n5563), .A2(MEM_stage_inst_dmem_n8417), .ZN(MEM_stage_inst_dmem_n5692) );
NOR2_X1 MEM_stage_inst_dmem_U5690 ( .A1(MEM_stage_inst_dmem_n5562), .A2(MEM_stage_inst_dmem_n5561), .ZN(MEM_stage_inst_dmem_n5563) );
NAND2_X1 MEM_stage_inst_dmem_U5689 ( .A1(MEM_stage_inst_dmem_n5560), .A2(MEM_stage_inst_dmem_n5559), .ZN(MEM_stage_inst_dmem_n5561) );
NOR2_X1 MEM_stage_inst_dmem_U5688 ( .A1(MEM_stage_inst_dmem_n5558), .A2(MEM_stage_inst_dmem_n5557), .ZN(MEM_stage_inst_dmem_n5559) );
NAND2_X1 MEM_stage_inst_dmem_U5687 ( .A1(MEM_stage_inst_dmem_n5556), .A2(MEM_stage_inst_dmem_n5555), .ZN(MEM_stage_inst_dmem_n5557) );
NOR2_X1 MEM_stage_inst_dmem_U5686 ( .A1(MEM_stage_inst_dmem_n5554), .A2(MEM_stage_inst_dmem_n5553), .ZN(MEM_stage_inst_dmem_n5555) );
NAND2_X1 MEM_stage_inst_dmem_U5685 ( .A1(MEM_stage_inst_dmem_n5552), .A2(MEM_stage_inst_dmem_n5551), .ZN(MEM_stage_inst_dmem_n5553) );
NAND2_X1 MEM_stage_inst_dmem_U5684 ( .A1(MEM_stage_inst_dmem_ram_3802), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n5551) );
NAND2_X1 MEM_stage_inst_dmem_U5683 ( .A1(MEM_stage_inst_dmem_ram_3738), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n5552) );
NAND2_X1 MEM_stage_inst_dmem_U5682 ( .A1(MEM_stage_inst_dmem_n5550), .A2(MEM_stage_inst_dmem_n5549), .ZN(MEM_stage_inst_dmem_n5554) );
NAND2_X1 MEM_stage_inst_dmem_U5681 ( .A1(MEM_stage_inst_dmem_ram_3850), .A2(MEM_stage_inst_dmem_n8472), .ZN(MEM_stage_inst_dmem_n5549) );
NAND2_X1 MEM_stage_inst_dmem_U5680 ( .A1(MEM_stage_inst_dmem_ram_3674), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n5550) );
NOR2_X1 MEM_stage_inst_dmem_U5679 ( .A1(MEM_stage_inst_dmem_n5548), .A2(MEM_stage_inst_dmem_n5547), .ZN(MEM_stage_inst_dmem_n5556) );
NAND2_X1 MEM_stage_inst_dmem_U5678 ( .A1(MEM_stage_inst_dmem_n5546), .A2(MEM_stage_inst_dmem_n5545), .ZN(MEM_stage_inst_dmem_n5547) );
NAND2_X1 MEM_stage_inst_dmem_U5677 ( .A1(MEM_stage_inst_dmem_ram_3322), .A2(MEM_stage_inst_dmem_n39), .ZN(MEM_stage_inst_dmem_n5545) );
NAND2_X1 MEM_stage_inst_dmem_U5676 ( .A1(MEM_stage_inst_dmem_ram_3706), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n5546) );
NAND2_X1 MEM_stage_inst_dmem_U5675 ( .A1(MEM_stage_inst_dmem_n5544), .A2(MEM_stage_inst_dmem_n5543), .ZN(MEM_stage_inst_dmem_n5548) );
NAND2_X1 MEM_stage_inst_dmem_U5674 ( .A1(MEM_stage_inst_dmem_ram_3402), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n5543) );
NAND2_X1 MEM_stage_inst_dmem_U5673 ( .A1(MEM_stage_inst_dmem_ram_3242), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n5544) );
NAND2_X1 MEM_stage_inst_dmem_U5672 ( .A1(MEM_stage_inst_dmem_n5542), .A2(MEM_stage_inst_dmem_n5541), .ZN(MEM_stage_inst_dmem_n5558) );
NOR2_X1 MEM_stage_inst_dmem_U5671 ( .A1(MEM_stage_inst_dmem_n5540), .A2(MEM_stage_inst_dmem_n5539), .ZN(MEM_stage_inst_dmem_n5541) );
NAND2_X1 MEM_stage_inst_dmem_U5670 ( .A1(MEM_stage_inst_dmem_n5538), .A2(MEM_stage_inst_dmem_n5537), .ZN(MEM_stage_inst_dmem_n5539) );
NAND2_X1 MEM_stage_inst_dmem_U5669 ( .A1(MEM_stage_inst_dmem_ram_3274), .A2(MEM_stage_inst_dmem_n8256), .ZN(MEM_stage_inst_dmem_n5537) );
NAND2_X1 MEM_stage_inst_dmem_U5668 ( .A1(MEM_stage_inst_dmem_ram_3898), .A2(MEM_stage_inst_dmem_n46), .ZN(MEM_stage_inst_dmem_n5538) );
NAND2_X1 MEM_stage_inst_dmem_U5667 ( .A1(MEM_stage_inst_dmem_n5536), .A2(MEM_stage_inst_dmem_n5535), .ZN(MEM_stage_inst_dmem_n5540) );
NAND2_X1 MEM_stage_inst_dmem_U5666 ( .A1(MEM_stage_inst_dmem_ram_3562), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n5535) );
NAND2_X1 MEM_stage_inst_dmem_U5665 ( .A1(MEM_stage_inst_dmem_ram_3690), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n5536) );
NOR2_X1 MEM_stage_inst_dmem_U5664 ( .A1(MEM_stage_inst_dmem_n5534), .A2(MEM_stage_inst_dmem_n5533), .ZN(MEM_stage_inst_dmem_n5542) );
NAND2_X1 MEM_stage_inst_dmem_U5663 ( .A1(MEM_stage_inst_dmem_n5532), .A2(MEM_stage_inst_dmem_n5531), .ZN(MEM_stage_inst_dmem_n5533) );
NAND2_X1 MEM_stage_inst_dmem_U5662 ( .A1(MEM_stage_inst_dmem_ram_3978), .A2(MEM_stage_inst_dmem_n8193), .ZN(MEM_stage_inst_dmem_n5531) );
NAND2_X1 MEM_stage_inst_dmem_U5661 ( .A1(MEM_stage_inst_dmem_ram_3770), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n5532) );
NAND2_X1 MEM_stage_inst_dmem_U5660 ( .A1(MEM_stage_inst_dmem_n5530), .A2(MEM_stage_inst_dmem_n5529), .ZN(MEM_stage_inst_dmem_n5534) );
NAND2_X1 MEM_stage_inst_dmem_U5659 ( .A1(MEM_stage_inst_dmem_ram_3098), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n5529) );
NAND2_X1 MEM_stage_inst_dmem_U5658 ( .A1(MEM_stage_inst_dmem_ram_3866), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n5530) );
NOR2_X1 MEM_stage_inst_dmem_U5657 ( .A1(MEM_stage_inst_dmem_n5528), .A2(MEM_stage_inst_dmem_n5527), .ZN(MEM_stage_inst_dmem_n5560) );
NAND2_X1 MEM_stage_inst_dmem_U5656 ( .A1(MEM_stage_inst_dmem_n5526), .A2(MEM_stage_inst_dmem_n5525), .ZN(MEM_stage_inst_dmem_n5527) );
NOR2_X1 MEM_stage_inst_dmem_U5655 ( .A1(MEM_stage_inst_dmem_n5524), .A2(MEM_stage_inst_dmem_n5523), .ZN(MEM_stage_inst_dmem_n5525) );
NAND2_X1 MEM_stage_inst_dmem_U5654 ( .A1(MEM_stage_inst_dmem_n5522), .A2(MEM_stage_inst_dmem_n5521), .ZN(MEM_stage_inst_dmem_n5523) );
NAND2_X1 MEM_stage_inst_dmem_U5653 ( .A1(MEM_stage_inst_dmem_ram_3434), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n5521) );
NAND2_X1 MEM_stage_inst_dmem_U5652 ( .A1(MEM_stage_inst_dmem_ram_3818), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n5522) );
NAND2_X1 MEM_stage_inst_dmem_U5651 ( .A1(MEM_stage_inst_dmem_n5520), .A2(MEM_stage_inst_dmem_n5519), .ZN(MEM_stage_inst_dmem_n5524) );
NAND2_X1 MEM_stage_inst_dmem_U5650 ( .A1(MEM_stage_inst_dmem_ram_3882), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n5519) );
NAND2_X1 MEM_stage_inst_dmem_U5649 ( .A1(MEM_stage_inst_dmem_ram_3530), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n5520) );
NOR2_X1 MEM_stage_inst_dmem_U5648 ( .A1(MEM_stage_inst_dmem_n5518), .A2(MEM_stage_inst_dmem_n5517), .ZN(MEM_stage_inst_dmem_n5526) );
NAND2_X1 MEM_stage_inst_dmem_U5647 ( .A1(MEM_stage_inst_dmem_n5516), .A2(MEM_stage_inst_dmem_n5515), .ZN(MEM_stage_inst_dmem_n5517) );
NAND2_X1 MEM_stage_inst_dmem_U5646 ( .A1(MEM_stage_inst_dmem_ram_3578), .A2(MEM_stage_inst_dmem_n64), .ZN(MEM_stage_inst_dmem_n5515) );
NAND2_X1 MEM_stage_inst_dmem_U5645 ( .A1(MEM_stage_inst_dmem_ram_4058), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n5516) );
NAND2_X1 MEM_stage_inst_dmem_U5644 ( .A1(MEM_stage_inst_dmem_n5514), .A2(MEM_stage_inst_dmem_n5513), .ZN(MEM_stage_inst_dmem_n5518) );
NAND2_X1 MEM_stage_inst_dmem_U5643 ( .A1(MEM_stage_inst_dmem_ram_3946), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n5513) );
NAND2_X1 MEM_stage_inst_dmem_U5642 ( .A1(MEM_stage_inst_dmem_ram_3482), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n5514) );
NAND2_X1 MEM_stage_inst_dmem_U5641 ( .A1(MEM_stage_inst_dmem_n5512), .A2(MEM_stage_inst_dmem_n5511), .ZN(MEM_stage_inst_dmem_n5528) );
NOR2_X1 MEM_stage_inst_dmem_U5640 ( .A1(MEM_stage_inst_dmem_n5510), .A2(MEM_stage_inst_dmem_n5509), .ZN(MEM_stage_inst_dmem_n5511) );
NAND2_X1 MEM_stage_inst_dmem_U5639 ( .A1(MEM_stage_inst_dmem_n5508), .A2(MEM_stage_inst_dmem_n5507), .ZN(MEM_stage_inst_dmem_n5509) );
NAND2_X1 MEM_stage_inst_dmem_U5638 ( .A1(MEM_stage_inst_dmem_ram_3642), .A2(MEM_stage_inst_dmem_n8169), .ZN(MEM_stage_inst_dmem_n5507) );
NAND2_X1 MEM_stage_inst_dmem_U5637 ( .A1(MEM_stage_inst_dmem_ram_3418), .A2(MEM_stage_inst_dmem_n3216), .ZN(MEM_stage_inst_dmem_n5508) );
NAND2_X1 MEM_stage_inst_dmem_U5636 ( .A1(MEM_stage_inst_dmem_n5506), .A2(MEM_stage_inst_dmem_n5505), .ZN(MEM_stage_inst_dmem_n5510) );
NAND2_X1 MEM_stage_inst_dmem_U5635 ( .A1(MEM_stage_inst_dmem_ram_3626), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n5505) );
NAND2_X1 MEM_stage_inst_dmem_U5634 ( .A1(MEM_stage_inst_dmem_ram_3658), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n5506) );
NOR2_X1 MEM_stage_inst_dmem_U5633 ( .A1(MEM_stage_inst_dmem_n5504), .A2(MEM_stage_inst_dmem_n5503), .ZN(MEM_stage_inst_dmem_n5512) );
NAND2_X1 MEM_stage_inst_dmem_U5632 ( .A1(MEM_stage_inst_dmem_n5502), .A2(MEM_stage_inst_dmem_n5501), .ZN(MEM_stage_inst_dmem_n5503) );
NAND2_X1 MEM_stage_inst_dmem_U5631 ( .A1(MEM_stage_inst_dmem_ram_3466), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n5501) );
NAND2_X1 MEM_stage_inst_dmem_U5630 ( .A1(MEM_stage_inst_dmem_ram_3450), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n5502) );
NAND2_X1 MEM_stage_inst_dmem_U5629 ( .A1(MEM_stage_inst_dmem_n5500), .A2(MEM_stage_inst_dmem_n5499), .ZN(MEM_stage_inst_dmem_n5504) );
NAND2_X1 MEM_stage_inst_dmem_U5628 ( .A1(MEM_stage_inst_dmem_ram_3786), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n5499) );
NAND2_X1 MEM_stage_inst_dmem_U5627 ( .A1(MEM_stage_inst_dmem_ram_3594), .A2(MEM_stage_inst_dmem_n8225), .ZN(MEM_stage_inst_dmem_n5500) );
NAND2_X1 MEM_stage_inst_dmem_U5626 ( .A1(MEM_stage_inst_dmem_n5498), .A2(MEM_stage_inst_dmem_n5497), .ZN(MEM_stage_inst_dmem_n5562) );
NOR2_X1 MEM_stage_inst_dmem_U5625 ( .A1(MEM_stage_inst_dmem_n5496), .A2(MEM_stage_inst_dmem_n5495), .ZN(MEM_stage_inst_dmem_n5497) );
NAND2_X1 MEM_stage_inst_dmem_U5624 ( .A1(MEM_stage_inst_dmem_n5494), .A2(MEM_stage_inst_dmem_n5493), .ZN(MEM_stage_inst_dmem_n5495) );
NOR2_X1 MEM_stage_inst_dmem_U5623 ( .A1(MEM_stage_inst_dmem_n5492), .A2(MEM_stage_inst_dmem_n5491), .ZN(MEM_stage_inst_dmem_n5493) );
NAND2_X1 MEM_stage_inst_dmem_U5622 ( .A1(MEM_stage_inst_dmem_n5490), .A2(MEM_stage_inst_dmem_n5489), .ZN(MEM_stage_inst_dmem_n5491) );
NAND2_X1 MEM_stage_inst_dmem_U5621 ( .A1(MEM_stage_inst_dmem_ram_3114), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n5489) );
NAND2_X1 MEM_stage_inst_dmem_U5620 ( .A1(MEM_stage_inst_dmem_ram_3354), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n5490) );
NAND2_X1 MEM_stage_inst_dmem_U5619 ( .A1(MEM_stage_inst_dmem_n5488), .A2(MEM_stage_inst_dmem_n5487), .ZN(MEM_stage_inst_dmem_n5492) );
NAND2_X1 MEM_stage_inst_dmem_U5618 ( .A1(MEM_stage_inst_dmem_ram_3834), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n5487) );
NAND2_X1 MEM_stage_inst_dmem_U5617 ( .A1(MEM_stage_inst_dmem_ram_3370), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n5488) );
NOR2_X1 MEM_stage_inst_dmem_U5616 ( .A1(MEM_stage_inst_dmem_n5486), .A2(MEM_stage_inst_dmem_n5485), .ZN(MEM_stage_inst_dmem_n5494) );
NAND2_X1 MEM_stage_inst_dmem_U5615 ( .A1(MEM_stage_inst_dmem_n5484), .A2(MEM_stage_inst_dmem_n5483), .ZN(MEM_stage_inst_dmem_n5485) );
NAND2_X1 MEM_stage_inst_dmem_U5614 ( .A1(MEM_stage_inst_dmem_ram_3994), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n5483) );
NAND2_X1 MEM_stage_inst_dmem_U5613 ( .A1(MEM_stage_inst_dmem_ram_3498), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n5484) );
NAND2_X1 MEM_stage_inst_dmem_U5612 ( .A1(MEM_stage_inst_dmem_n5482), .A2(MEM_stage_inst_dmem_n5481), .ZN(MEM_stage_inst_dmem_n5486) );
NAND2_X1 MEM_stage_inst_dmem_U5611 ( .A1(MEM_stage_inst_dmem_ram_3930), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n5481) );
NAND2_X1 MEM_stage_inst_dmem_U5610 ( .A1(MEM_stage_inst_dmem_ram_4042), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n5482) );
NAND2_X1 MEM_stage_inst_dmem_U5609 ( .A1(MEM_stage_inst_dmem_n5480), .A2(MEM_stage_inst_dmem_n5479), .ZN(MEM_stage_inst_dmem_n5496) );
NOR2_X1 MEM_stage_inst_dmem_U5608 ( .A1(MEM_stage_inst_dmem_n5478), .A2(MEM_stage_inst_dmem_n5477), .ZN(MEM_stage_inst_dmem_n5479) );
NAND2_X1 MEM_stage_inst_dmem_U5607 ( .A1(MEM_stage_inst_dmem_n5476), .A2(MEM_stage_inst_dmem_n5475), .ZN(MEM_stage_inst_dmem_n5477) );
NAND2_X1 MEM_stage_inst_dmem_U5606 ( .A1(MEM_stage_inst_dmem_ram_3962), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n5475) );
NAND2_X1 MEM_stage_inst_dmem_U5605 ( .A1(MEM_stage_inst_dmem_ram_3146), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n5476) );
NAND2_X1 MEM_stage_inst_dmem_U5604 ( .A1(MEM_stage_inst_dmem_n5474), .A2(MEM_stage_inst_dmem_n5473), .ZN(MEM_stage_inst_dmem_n5478) );
NAND2_X1 MEM_stage_inst_dmem_U5603 ( .A1(MEM_stage_inst_dmem_ram_3514), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n5473) );
NAND2_X1 MEM_stage_inst_dmem_U5602 ( .A1(MEM_stage_inst_dmem_ram_3290), .A2(MEM_stage_inst_dmem_n8206), .ZN(MEM_stage_inst_dmem_n5474) );
NOR2_X1 MEM_stage_inst_dmem_U5601 ( .A1(MEM_stage_inst_dmem_n5472), .A2(MEM_stage_inst_dmem_n5471), .ZN(MEM_stage_inst_dmem_n5480) );
NAND2_X1 MEM_stage_inst_dmem_U5600 ( .A1(MEM_stage_inst_dmem_n5470), .A2(MEM_stage_inst_dmem_n5469), .ZN(MEM_stage_inst_dmem_n5471) );
NAND2_X1 MEM_stage_inst_dmem_U5599 ( .A1(MEM_stage_inst_dmem_ram_3306), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n5469) );
NAND2_X1 MEM_stage_inst_dmem_U5598 ( .A1(MEM_stage_inst_dmem_ram_3226), .A2(MEM_stage_inst_dmem_n44), .ZN(MEM_stage_inst_dmem_n5470) );
NAND2_X1 MEM_stage_inst_dmem_U5597 ( .A1(MEM_stage_inst_dmem_n5468), .A2(MEM_stage_inst_dmem_n5467), .ZN(MEM_stage_inst_dmem_n5472) );
NAND2_X1 MEM_stage_inst_dmem_U5596 ( .A1(MEM_stage_inst_dmem_ram_4090), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n5467) );
NAND2_X1 MEM_stage_inst_dmem_U5595 ( .A1(MEM_stage_inst_dmem_ram_3178), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n5468) );
NOR2_X1 MEM_stage_inst_dmem_U5594 ( .A1(MEM_stage_inst_dmem_n5466), .A2(MEM_stage_inst_dmem_n5465), .ZN(MEM_stage_inst_dmem_n5498) );
NAND2_X1 MEM_stage_inst_dmem_U5593 ( .A1(MEM_stage_inst_dmem_n5464), .A2(MEM_stage_inst_dmem_n5463), .ZN(MEM_stage_inst_dmem_n5465) );
NOR2_X1 MEM_stage_inst_dmem_U5592 ( .A1(MEM_stage_inst_dmem_n5462), .A2(MEM_stage_inst_dmem_n5461), .ZN(MEM_stage_inst_dmem_n5463) );
NAND2_X1 MEM_stage_inst_dmem_U5591 ( .A1(MEM_stage_inst_dmem_n5460), .A2(MEM_stage_inst_dmem_n5459), .ZN(MEM_stage_inst_dmem_n5461) );
NAND2_X1 MEM_stage_inst_dmem_U5590 ( .A1(MEM_stage_inst_dmem_ram_3722), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n5459) );
NAND2_X1 MEM_stage_inst_dmem_U5589 ( .A1(MEM_stage_inst_dmem_ram_4010), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n5460) );
NAND2_X1 MEM_stage_inst_dmem_U5588 ( .A1(MEM_stage_inst_dmem_n5458), .A2(MEM_stage_inst_dmem_n5457), .ZN(MEM_stage_inst_dmem_n5462) );
NAND2_X1 MEM_stage_inst_dmem_U5587 ( .A1(MEM_stage_inst_dmem_ram_3194), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n5457) );
NAND2_X1 MEM_stage_inst_dmem_U5586 ( .A1(MEM_stage_inst_dmem_ram_3610), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n5458) );
NOR2_X1 MEM_stage_inst_dmem_U5585 ( .A1(MEM_stage_inst_dmem_n5456), .A2(MEM_stage_inst_dmem_n5455), .ZN(MEM_stage_inst_dmem_n5464) );
NAND2_X1 MEM_stage_inst_dmem_U5584 ( .A1(MEM_stage_inst_dmem_n5454), .A2(MEM_stage_inst_dmem_n5453), .ZN(MEM_stage_inst_dmem_n5455) );
NAND2_X1 MEM_stage_inst_dmem_U5583 ( .A1(MEM_stage_inst_dmem_ram_3386), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n5453) );
NAND2_X1 MEM_stage_inst_dmem_U5582 ( .A1(MEM_stage_inst_dmem_ram_3162), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n5454) );
NAND2_X1 MEM_stage_inst_dmem_U5581 ( .A1(MEM_stage_inst_dmem_n5452), .A2(MEM_stage_inst_dmem_n5451), .ZN(MEM_stage_inst_dmem_n5456) );
NAND2_X1 MEM_stage_inst_dmem_U5580 ( .A1(MEM_stage_inst_dmem_ram_3546), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n5451) );
NAND2_X1 MEM_stage_inst_dmem_U5579 ( .A1(MEM_stage_inst_dmem_ram_3338), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n5452) );
NAND2_X1 MEM_stage_inst_dmem_U5578 ( .A1(MEM_stage_inst_dmem_n5450), .A2(MEM_stage_inst_dmem_n5449), .ZN(MEM_stage_inst_dmem_n5466) );
NOR2_X1 MEM_stage_inst_dmem_U5577 ( .A1(MEM_stage_inst_dmem_n5448), .A2(MEM_stage_inst_dmem_n5447), .ZN(MEM_stage_inst_dmem_n5449) );
NAND2_X1 MEM_stage_inst_dmem_U5576 ( .A1(MEM_stage_inst_dmem_n5446), .A2(MEM_stage_inst_dmem_n5445), .ZN(MEM_stage_inst_dmem_n5447) );
NAND2_X1 MEM_stage_inst_dmem_U5575 ( .A1(MEM_stage_inst_dmem_ram_3130), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n5445) );
NAND2_X1 MEM_stage_inst_dmem_U5574 ( .A1(MEM_stage_inst_dmem_ram_3210), .A2(MEM_stage_inst_dmem_n8174), .ZN(MEM_stage_inst_dmem_n5446) );
NAND2_X1 MEM_stage_inst_dmem_U5573 ( .A1(MEM_stage_inst_dmem_n5444), .A2(MEM_stage_inst_dmem_n5443), .ZN(MEM_stage_inst_dmem_n5448) );
NAND2_X1 MEM_stage_inst_dmem_U5572 ( .A1(MEM_stage_inst_dmem_ram_4074), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n5443) );
NAND2_X1 MEM_stage_inst_dmem_U5571 ( .A1(MEM_stage_inst_dmem_ram_3258), .A2(MEM_stage_inst_dmem_n8434), .ZN(MEM_stage_inst_dmem_n5444) );
NOR2_X1 MEM_stage_inst_dmem_U5570 ( .A1(MEM_stage_inst_dmem_n5442), .A2(MEM_stage_inst_dmem_n5441), .ZN(MEM_stage_inst_dmem_n5450) );
NAND2_X1 MEM_stage_inst_dmem_U5569 ( .A1(MEM_stage_inst_dmem_n5440), .A2(MEM_stage_inst_dmem_n5439), .ZN(MEM_stage_inst_dmem_n5441) );
NAND2_X1 MEM_stage_inst_dmem_U5568 ( .A1(MEM_stage_inst_dmem_ram_3754), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n5439) );
NAND2_X1 MEM_stage_inst_dmem_U5567 ( .A1(MEM_stage_inst_dmem_ram_3082), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n5440) );
NAND2_X1 MEM_stage_inst_dmem_U5566 ( .A1(MEM_stage_inst_dmem_n5438), .A2(MEM_stage_inst_dmem_n5437), .ZN(MEM_stage_inst_dmem_n5442) );
NAND2_X1 MEM_stage_inst_dmem_U5565 ( .A1(MEM_stage_inst_dmem_ram_3914), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n5437) );
NAND2_X1 MEM_stage_inst_dmem_U5564 ( .A1(MEM_stage_inst_dmem_ram_4026), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n5438) );
NAND2_X1 MEM_stage_inst_dmem_U5563 ( .A1(MEM_stage_inst_dmem_n5436), .A2(MEM_stage_inst_dmem_n5435), .ZN(MEM_stage_inst_mem_read_data_9) );
NOR2_X1 MEM_stage_inst_dmem_U5562 ( .A1(MEM_stage_inst_dmem_n5434), .A2(MEM_stage_inst_dmem_n5433), .ZN(MEM_stage_inst_dmem_n5435) );
NOR2_X1 MEM_stage_inst_dmem_U5561 ( .A1(MEM_stage_inst_dmem_n5432), .A2(MEM_stage_inst_dmem_n8551), .ZN(MEM_stage_inst_dmem_n5433) );
NOR2_X1 MEM_stage_inst_dmem_U5560 ( .A1(MEM_stage_inst_dmem_n5431), .A2(MEM_stage_inst_dmem_n5430), .ZN(MEM_stage_inst_dmem_n5432) );
NAND2_X1 MEM_stage_inst_dmem_U5559 ( .A1(MEM_stage_inst_dmem_n5429), .A2(MEM_stage_inst_dmem_n5428), .ZN(MEM_stage_inst_dmem_n5430) );
NOR2_X1 MEM_stage_inst_dmem_U5558 ( .A1(MEM_stage_inst_dmem_n5427), .A2(MEM_stage_inst_dmem_n5426), .ZN(MEM_stage_inst_dmem_n5428) );
NAND2_X1 MEM_stage_inst_dmem_U5557 ( .A1(MEM_stage_inst_dmem_n5425), .A2(MEM_stage_inst_dmem_n5424), .ZN(MEM_stage_inst_dmem_n5426) );
NOR2_X1 MEM_stage_inst_dmem_U5556 ( .A1(MEM_stage_inst_dmem_n5423), .A2(MEM_stage_inst_dmem_n5422), .ZN(MEM_stage_inst_dmem_n5424) );
NAND2_X1 MEM_stage_inst_dmem_U5555 ( .A1(MEM_stage_inst_dmem_n5421), .A2(MEM_stage_inst_dmem_n5420), .ZN(MEM_stage_inst_dmem_n5422) );
NAND2_X1 MEM_stage_inst_dmem_U5554 ( .A1(MEM_stage_inst_dmem_ram_425), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n5420) );
NAND2_X1 MEM_stage_inst_dmem_U5553 ( .A1(MEM_stage_inst_dmem_ram_217), .A2(MEM_stage_inst_dmem_n51), .ZN(MEM_stage_inst_dmem_n5421) );
NAND2_X1 MEM_stage_inst_dmem_U5552 ( .A1(MEM_stage_inst_dmem_n5419), .A2(MEM_stage_inst_dmem_n5418), .ZN(MEM_stage_inst_dmem_n5423) );
NAND2_X1 MEM_stage_inst_dmem_U5551 ( .A1(MEM_stage_inst_dmem_ram_457), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n5418) );
NAND2_X1 MEM_stage_inst_dmem_U5550 ( .A1(MEM_stage_inst_dmem_ram_617), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n5419) );
NOR2_X1 MEM_stage_inst_dmem_U5549 ( .A1(MEM_stage_inst_dmem_n5417), .A2(MEM_stage_inst_dmem_n5416), .ZN(MEM_stage_inst_dmem_n5425) );
NAND2_X1 MEM_stage_inst_dmem_U5548 ( .A1(MEM_stage_inst_dmem_n5415), .A2(MEM_stage_inst_dmem_n5414), .ZN(MEM_stage_inst_dmem_n5416) );
NAND2_X1 MEM_stage_inst_dmem_U5547 ( .A1(MEM_stage_inst_dmem_ram_681), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n5414) );
NAND2_X1 MEM_stage_inst_dmem_U5546 ( .A1(MEM_stage_inst_dmem_ram_169), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n5415) );
NAND2_X1 MEM_stage_inst_dmem_U5545 ( .A1(MEM_stage_inst_dmem_n5413), .A2(MEM_stage_inst_dmem_n5412), .ZN(MEM_stage_inst_dmem_n5417) );
NAND2_X1 MEM_stage_inst_dmem_U5544 ( .A1(MEM_stage_inst_dmem_ram_777), .A2(MEM_stage_inst_dmem_n37), .ZN(MEM_stage_inst_dmem_n5412) );
NAND2_X1 MEM_stage_inst_dmem_U5543 ( .A1(MEM_stage_inst_dmem_ram_985), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n5413) );
NAND2_X1 MEM_stage_inst_dmem_U5542 ( .A1(MEM_stage_inst_dmem_n5411), .A2(MEM_stage_inst_dmem_n5410), .ZN(MEM_stage_inst_dmem_n5427) );
NOR2_X1 MEM_stage_inst_dmem_U5541 ( .A1(MEM_stage_inst_dmem_n5409), .A2(MEM_stage_inst_dmem_n5408), .ZN(MEM_stage_inst_dmem_n5410) );
NAND2_X1 MEM_stage_inst_dmem_U5540 ( .A1(MEM_stage_inst_dmem_n5407), .A2(MEM_stage_inst_dmem_n5406), .ZN(MEM_stage_inst_dmem_n5408) );
NAND2_X1 MEM_stage_inst_dmem_U5539 ( .A1(MEM_stage_inst_dmem_ram_393), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n5406) );
NAND2_X1 MEM_stage_inst_dmem_U5538 ( .A1(MEM_stage_inst_dmem_ram_345), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n5407) );
NAND2_X1 MEM_stage_inst_dmem_U5537 ( .A1(MEM_stage_inst_dmem_n5405), .A2(MEM_stage_inst_dmem_n5404), .ZN(MEM_stage_inst_dmem_n5409) );
NAND2_X1 MEM_stage_inst_dmem_U5536 ( .A1(MEM_stage_inst_dmem_ram_921), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n5404) );
NAND2_X1 MEM_stage_inst_dmem_U5535 ( .A1(MEM_stage_inst_dmem_ram_281), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n5405) );
NOR2_X1 MEM_stage_inst_dmem_U5534 ( .A1(MEM_stage_inst_dmem_n5403), .A2(MEM_stage_inst_dmem_n5402), .ZN(MEM_stage_inst_dmem_n5411) );
NAND2_X1 MEM_stage_inst_dmem_U5533 ( .A1(MEM_stage_inst_dmem_n5401), .A2(MEM_stage_inst_dmem_n5400), .ZN(MEM_stage_inst_dmem_n5402) );
NAND2_X1 MEM_stage_inst_dmem_U5532 ( .A1(MEM_stage_inst_dmem_ram_233), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n5400) );
NAND2_X1 MEM_stage_inst_dmem_U5531 ( .A1(MEM_stage_inst_dmem_ram_105), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n5401) );
NAND2_X1 MEM_stage_inst_dmem_U5530 ( .A1(MEM_stage_inst_dmem_n5399), .A2(MEM_stage_inst_dmem_n5398), .ZN(MEM_stage_inst_dmem_n5403) );
NAND2_X1 MEM_stage_inst_dmem_U5529 ( .A1(MEM_stage_inst_dmem_ram_201), .A2(MEM_stage_inst_dmem_n36), .ZN(MEM_stage_inst_dmem_n5398) );
NAND2_X1 MEM_stage_inst_dmem_U5528 ( .A1(MEM_stage_inst_dmem_ram_585), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n5399) );
NOR2_X1 MEM_stage_inst_dmem_U5527 ( .A1(MEM_stage_inst_dmem_n5397), .A2(MEM_stage_inst_dmem_n5396), .ZN(MEM_stage_inst_dmem_n5429) );
NAND2_X1 MEM_stage_inst_dmem_U5526 ( .A1(MEM_stage_inst_dmem_n5395), .A2(MEM_stage_inst_dmem_n5394), .ZN(MEM_stage_inst_dmem_n5396) );
NOR2_X1 MEM_stage_inst_dmem_U5525 ( .A1(MEM_stage_inst_dmem_n5393), .A2(MEM_stage_inst_dmem_n5392), .ZN(MEM_stage_inst_dmem_n5394) );
NAND2_X1 MEM_stage_inst_dmem_U5524 ( .A1(MEM_stage_inst_dmem_n5391), .A2(MEM_stage_inst_dmem_n5390), .ZN(MEM_stage_inst_dmem_n5392) );
NAND2_X1 MEM_stage_inst_dmem_U5523 ( .A1(MEM_stage_inst_dmem_ram_649), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n5390) );
NAND2_X1 MEM_stage_inst_dmem_U5522 ( .A1(MEM_stage_inst_dmem_ram_665), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n5391) );
NAND2_X1 MEM_stage_inst_dmem_U5521 ( .A1(MEM_stage_inst_dmem_n5389), .A2(MEM_stage_inst_dmem_n5388), .ZN(MEM_stage_inst_dmem_n5393) );
NAND2_X1 MEM_stage_inst_dmem_U5520 ( .A1(MEM_stage_inst_dmem_ram_409), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n5388) );
NAND2_X1 MEM_stage_inst_dmem_U5519 ( .A1(MEM_stage_inst_dmem_ram_1017), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n5389) );
NOR2_X1 MEM_stage_inst_dmem_U5518 ( .A1(MEM_stage_inst_dmem_n5387), .A2(MEM_stage_inst_dmem_n5386), .ZN(MEM_stage_inst_dmem_n5395) );
NAND2_X1 MEM_stage_inst_dmem_U5517 ( .A1(MEM_stage_inst_dmem_n5385), .A2(MEM_stage_inst_dmem_n5384), .ZN(MEM_stage_inst_dmem_n5386) );
NAND2_X1 MEM_stage_inst_dmem_U5516 ( .A1(MEM_stage_inst_dmem_ram_553), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n5384) );
NAND2_X1 MEM_stage_inst_dmem_U5515 ( .A1(MEM_stage_inst_dmem_ram_793), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n5385) );
NAND2_X1 MEM_stage_inst_dmem_U5514 ( .A1(MEM_stage_inst_dmem_n5383), .A2(MEM_stage_inst_dmem_n5382), .ZN(MEM_stage_inst_dmem_n5387) );
NAND2_X1 MEM_stage_inst_dmem_U5513 ( .A1(MEM_stage_inst_dmem_ram_841), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n5382) );
NAND2_X1 MEM_stage_inst_dmem_U5512 ( .A1(MEM_stage_inst_dmem_ram_937), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n5383) );
NAND2_X1 MEM_stage_inst_dmem_U5511 ( .A1(MEM_stage_inst_dmem_n5381), .A2(MEM_stage_inst_dmem_n5380), .ZN(MEM_stage_inst_dmem_n5397) );
NOR2_X1 MEM_stage_inst_dmem_U5510 ( .A1(MEM_stage_inst_dmem_n5379), .A2(MEM_stage_inst_dmem_n5378), .ZN(MEM_stage_inst_dmem_n5380) );
NAND2_X1 MEM_stage_inst_dmem_U5509 ( .A1(MEM_stage_inst_dmem_n5377), .A2(MEM_stage_inst_dmem_n5376), .ZN(MEM_stage_inst_dmem_n5378) );
NAND2_X1 MEM_stage_inst_dmem_U5508 ( .A1(MEM_stage_inst_dmem_ram_713), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n5376) );
NAND2_X1 MEM_stage_inst_dmem_U5507 ( .A1(MEM_stage_inst_dmem_ram_377), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n5377) );
NAND2_X1 MEM_stage_inst_dmem_U5506 ( .A1(MEM_stage_inst_dmem_n5375), .A2(MEM_stage_inst_dmem_n5374), .ZN(MEM_stage_inst_dmem_n5379) );
NAND2_X1 MEM_stage_inst_dmem_U5505 ( .A1(MEM_stage_inst_dmem_ram_569), .A2(MEM_stage_inst_dmem_n41), .ZN(MEM_stage_inst_dmem_n5374) );
NAND2_X1 MEM_stage_inst_dmem_U5504 ( .A1(MEM_stage_inst_dmem_ram_601), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n5375) );
NOR2_X1 MEM_stage_inst_dmem_U5503 ( .A1(MEM_stage_inst_dmem_n5373), .A2(MEM_stage_inst_dmem_n5372), .ZN(MEM_stage_inst_dmem_n5381) );
NAND2_X1 MEM_stage_inst_dmem_U5502 ( .A1(MEM_stage_inst_dmem_n5371), .A2(MEM_stage_inst_dmem_n5370), .ZN(MEM_stage_inst_dmem_n5372) );
NAND2_X1 MEM_stage_inst_dmem_U5501 ( .A1(MEM_stage_inst_dmem_ram_361), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n5370) );
NAND2_X1 MEM_stage_inst_dmem_U5500 ( .A1(MEM_stage_inst_dmem_ram_953), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n5371) );
NAND2_X1 MEM_stage_inst_dmem_U5499 ( .A1(MEM_stage_inst_dmem_n5369), .A2(MEM_stage_inst_dmem_n5368), .ZN(MEM_stage_inst_dmem_n5373) );
NAND2_X1 MEM_stage_inst_dmem_U5498 ( .A1(MEM_stage_inst_dmem_ram_505), .A2(MEM_stage_inst_dmem_n64), .ZN(MEM_stage_inst_dmem_n5368) );
NAND2_X1 MEM_stage_inst_dmem_U5497 ( .A1(MEM_stage_inst_dmem_ram_329), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n5369) );
NAND2_X1 MEM_stage_inst_dmem_U5496 ( .A1(MEM_stage_inst_dmem_n5367), .A2(MEM_stage_inst_dmem_n5366), .ZN(MEM_stage_inst_dmem_n5431) );
NOR2_X1 MEM_stage_inst_dmem_U5495 ( .A1(MEM_stage_inst_dmem_n5365), .A2(MEM_stage_inst_dmem_n5364), .ZN(MEM_stage_inst_dmem_n5366) );
NAND2_X1 MEM_stage_inst_dmem_U5494 ( .A1(MEM_stage_inst_dmem_n5363), .A2(MEM_stage_inst_dmem_n5362), .ZN(MEM_stage_inst_dmem_n5364) );
NOR2_X1 MEM_stage_inst_dmem_U5493 ( .A1(MEM_stage_inst_dmem_n5361), .A2(MEM_stage_inst_dmem_n5360), .ZN(MEM_stage_inst_dmem_n5362) );
NAND2_X1 MEM_stage_inst_dmem_U5492 ( .A1(MEM_stage_inst_dmem_n5359), .A2(MEM_stage_inst_dmem_n5358), .ZN(MEM_stage_inst_dmem_n5360) );
NAND2_X1 MEM_stage_inst_dmem_U5491 ( .A1(MEM_stage_inst_dmem_ram_761), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n5358) );
NAND2_X1 MEM_stage_inst_dmem_U5490 ( .A1(MEM_stage_inst_dmem_ram_25), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n5359) );
NAND2_X1 MEM_stage_inst_dmem_U5489 ( .A1(MEM_stage_inst_dmem_n5357), .A2(MEM_stage_inst_dmem_n5356), .ZN(MEM_stage_inst_dmem_n5361) );
NAND2_X1 MEM_stage_inst_dmem_U5488 ( .A1(MEM_stage_inst_dmem_ram_969), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n5356) );
NAND2_X1 MEM_stage_inst_dmem_U5487 ( .A1(MEM_stage_inst_dmem_ram_825), .A2(MEM_stage_inst_dmem_n46), .ZN(MEM_stage_inst_dmem_n5357) );
NOR2_X1 MEM_stage_inst_dmem_U5486 ( .A1(MEM_stage_inst_dmem_n5355), .A2(MEM_stage_inst_dmem_n5354), .ZN(MEM_stage_inst_dmem_n5363) );
NAND2_X1 MEM_stage_inst_dmem_U5485 ( .A1(MEM_stage_inst_dmem_n5353), .A2(MEM_stage_inst_dmem_n5352), .ZN(MEM_stage_inst_dmem_n5354) );
NAND2_X1 MEM_stage_inst_dmem_U5484 ( .A1(MEM_stage_inst_dmem_ram_185), .A2(MEM_stage_inst_dmem_n55), .ZN(MEM_stage_inst_dmem_n5352) );
NAND2_X1 MEM_stage_inst_dmem_U5483 ( .A1(MEM_stage_inst_dmem_ram_9), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n5353) );
NAND2_X1 MEM_stage_inst_dmem_U5482 ( .A1(MEM_stage_inst_dmem_n5351), .A2(MEM_stage_inst_dmem_n5350), .ZN(MEM_stage_inst_dmem_n5355) );
NAND2_X1 MEM_stage_inst_dmem_U5481 ( .A1(MEM_stage_inst_dmem_ram_57), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n5350) );
NAND2_X1 MEM_stage_inst_dmem_U5480 ( .A1(MEM_stage_inst_dmem_ram_745), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n5351) );
NAND2_X1 MEM_stage_inst_dmem_U5479 ( .A1(MEM_stage_inst_dmem_n5349), .A2(MEM_stage_inst_dmem_n5348), .ZN(MEM_stage_inst_dmem_n5365) );
NOR2_X1 MEM_stage_inst_dmem_U5478 ( .A1(MEM_stage_inst_dmem_n5347), .A2(MEM_stage_inst_dmem_n5346), .ZN(MEM_stage_inst_dmem_n5348) );
NAND2_X1 MEM_stage_inst_dmem_U5477 ( .A1(MEM_stage_inst_dmem_n5345), .A2(MEM_stage_inst_dmem_n5344), .ZN(MEM_stage_inst_dmem_n5346) );
NAND2_X1 MEM_stage_inst_dmem_U5476 ( .A1(MEM_stage_inst_dmem_ram_313), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n5344) );
NAND2_X1 MEM_stage_inst_dmem_U5475 ( .A1(MEM_stage_inst_dmem_ram_249), .A2(MEM_stage_inst_dmem_n39), .ZN(MEM_stage_inst_dmem_n5345) );
NAND2_X1 MEM_stage_inst_dmem_U5474 ( .A1(MEM_stage_inst_dmem_n5343), .A2(MEM_stage_inst_dmem_n5342), .ZN(MEM_stage_inst_dmem_n5347) );
NAND2_X1 MEM_stage_inst_dmem_U5473 ( .A1(MEM_stage_inst_dmem_ram_633), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n5342) );
NAND2_X1 MEM_stage_inst_dmem_U5472 ( .A1(MEM_stage_inst_dmem_ram_729), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n5343) );
NOR2_X1 MEM_stage_inst_dmem_U5471 ( .A1(MEM_stage_inst_dmem_n5341), .A2(MEM_stage_inst_dmem_n5340), .ZN(MEM_stage_inst_dmem_n5349) );
NAND2_X1 MEM_stage_inst_dmem_U5470 ( .A1(MEM_stage_inst_dmem_n5339), .A2(MEM_stage_inst_dmem_n5338), .ZN(MEM_stage_inst_dmem_n5340) );
NAND2_X1 MEM_stage_inst_dmem_U5469 ( .A1(MEM_stage_inst_dmem_ram_41), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n5338) );
NAND2_X1 MEM_stage_inst_dmem_U5468 ( .A1(MEM_stage_inst_dmem_ram_265), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n5339) );
NAND2_X1 MEM_stage_inst_dmem_U5467 ( .A1(MEM_stage_inst_dmem_n5337), .A2(MEM_stage_inst_dmem_n5336), .ZN(MEM_stage_inst_dmem_n5341) );
NAND2_X1 MEM_stage_inst_dmem_U5466 ( .A1(MEM_stage_inst_dmem_ram_873), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n5336) );
NAND2_X1 MEM_stage_inst_dmem_U5465 ( .A1(MEM_stage_inst_dmem_ram_697), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n5337) );
NOR2_X1 MEM_stage_inst_dmem_U5464 ( .A1(MEM_stage_inst_dmem_n5335), .A2(MEM_stage_inst_dmem_n5334), .ZN(MEM_stage_inst_dmem_n5367) );
NAND2_X1 MEM_stage_inst_dmem_U5463 ( .A1(MEM_stage_inst_dmem_n5333), .A2(MEM_stage_inst_dmem_n5332), .ZN(MEM_stage_inst_dmem_n5334) );
NOR2_X1 MEM_stage_inst_dmem_U5462 ( .A1(MEM_stage_inst_dmem_n5331), .A2(MEM_stage_inst_dmem_n5330), .ZN(MEM_stage_inst_dmem_n5332) );
NAND2_X1 MEM_stage_inst_dmem_U5461 ( .A1(MEM_stage_inst_dmem_n5329), .A2(MEM_stage_inst_dmem_n5328), .ZN(MEM_stage_inst_dmem_n5330) );
NAND2_X1 MEM_stage_inst_dmem_U5460 ( .A1(MEM_stage_inst_dmem_ram_889), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n5328) );
NAND2_X1 MEM_stage_inst_dmem_U5459 ( .A1(MEM_stage_inst_dmem_ram_521), .A2(MEM_stage_inst_dmem_n71), .ZN(MEM_stage_inst_dmem_n5329) );
NAND2_X1 MEM_stage_inst_dmem_U5458 ( .A1(MEM_stage_inst_dmem_n5327), .A2(MEM_stage_inst_dmem_n5326), .ZN(MEM_stage_inst_dmem_n5331) );
NAND2_X1 MEM_stage_inst_dmem_U5457 ( .A1(MEM_stage_inst_dmem_ram_441), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n5326) );
NAND2_X1 MEM_stage_inst_dmem_U5456 ( .A1(MEM_stage_inst_dmem_ram_89), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n5327) );
NOR2_X1 MEM_stage_inst_dmem_U5455 ( .A1(MEM_stage_inst_dmem_n5325), .A2(MEM_stage_inst_dmem_n5324), .ZN(MEM_stage_inst_dmem_n5333) );
NAND2_X1 MEM_stage_inst_dmem_U5454 ( .A1(MEM_stage_inst_dmem_n5323), .A2(MEM_stage_inst_dmem_n5322), .ZN(MEM_stage_inst_dmem_n5324) );
NAND2_X1 MEM_stage_inst_dmem_U5453 ( .A1(MEM_stage_inst_dmem_ram_489), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n5322) );
NAND2_X1 MEM_stage_inst_dmem_U5452 ( .A1(MEM_stage_inst_dmem_ram_121), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n5323) );
NAND2_X1 MEM_stage_inst_dmem_U5451 ( .A1(MEM_stage_inst_dmem_n5321), .A2(MEM_stage_inst_dmem_n5320), .ZN(MEM_stage_inst_dmem_n5325) );
NAND2_X1 MEM_stage_inst_dmem_U5450 ( .A1(MEM_stage_inst_dmem_ram_857), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n5320) );
NAND2_X1 MEM_stage_inst_dmem_U5449 ( .A1(MEM_stage_inst_dmem_ram_73), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n5321) );
NAND2_X1 MEM_stage_inst_dmem_U5448 ( .A1(MEM_stage_inst_dmem_n5319), .A2(MEM_stage_inst_dmem_n5318), .ZN(MEM_stage_inst_dmem_n5335) );
NOR2_X1 MEM_stage_inst_dmem_U5447 ( .A1(MEM_stage_inst_dmem_n5317), .A2(MEM_stage_inst_dmem_n5316), .ZN(MEM_stage_inst_dmem_n5318) );
NAND2_X1 MEM_stage_inst_dmem_U5446 ( .A1(MEM_stage_inst_dmem_n5315), .A2(MEM_stage_inst_dmem_n5314), .ZN(MEM_stage_inst_dmem_n5316) );
NAND2_X1 MEM_stage_inst_dmem_U5445 ( .A1(MEM_stage_inst_dmem_ram_905), .A2(MEM_stage_inst_dmem_n72), .ZN(MEM_stage_inst_dmem_n5314) );
NAND2_X1 MEM_stage_inst_dmem_U5444 ( .A1(MEM_stage_inst_dmem_ram_297), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n5315) );
NAND2_X1 MEM_stage_inst_dmem_U5443 ( .A1(MEM_stage_inst_dmem_n5313), .A2(MEM_stage_inst_dmem_n5312), .ZN(MEM_stage_inst_dmem_n5317) );
NAND2_X1 MEM_stage_inst_dmem_U5442 ( .A1(MEM_stage_inst_dmem_ram_137), .A2(MEM_stage_inst_dmem_n61), .ZN(MEM_stage_inst_dmem_n5312) );
NAND2_X1 MEM_stage_inst_dmem_U5441 ( .A1(MEM_stage_inst_dmem_ram_537), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n5313) );
NOR2_X1 MEM_stage_inst_dmem_U5440 ( .A1(MEM_stage_inst_dmem_n5311), .A2(MEM_stage_inst_dmem_n5310), .ZN(MEM_stage_inst_dmem_n5319) );
NAND2_X1 MEM_stage_inst_dmem_U5439 ( .A1(MEM_stage_inst_dmem_n5309), .A2(MEM_stage_inst_dmem_n5308), .ZN(MEM_stage_inst_dmem_n5310) );
NAND2_X1 MEM_stage_inst_dmem_U5438 ( .A1(MEM_stage_inst_dmem_ram_809), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n5308) );
NAND2_X1 MEM_stage_inst_dmem_U5437 ( .A1(MEM_stage_inst_dmem_ram_153), .A2(MEM_stage_inst_dmem_n44), .ZN(MEM_stage_inst_dmem_n5309) );
NAND2_X1 MEM_stage_inst_dmem_U5436 ( .A1(MEM_stage_inst_dmem_n5307), .A2(MEM_stage_inst_dmem_n5306), .ZN(MEM_stage_inst_dmem_n5311) );
NAND2_X1 MEM_stage_inst_dmem_U5435 ( .A1(MEM_stage_inst_dmem_ram_1001), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n5306) );
NAND2_X1 MEM_stage_inst_dmem_U5434 ( .A1(MEM_stage_inst_dmem_ram_473), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n5307) );
NOR2_X1 MEM_stage_inst_dmem_U5433 ( .A1(MEM_stage_inst_dmem_n5305), .A2(MEM_stage_inst_dmem_n8417), .ZN(MEM_stage_inst_dmem_n5434) );
NOR2_X1 MEM_stage_inst_dmem_U5432 ( .A1(MEM_stage_inst_dmem_n5304), .A2(MEM_stage_inst_dmem_n5303), .ZN(MEM_stage_inst_dmem_n5305) );
NAND2_X1 MEM_stage_inst_dmem_U5431 ( .A1(MEM_stage_inst_dmem_n5302), .A2(MEM_stage_inst_dmem_n5301), .ZN(MEM_stage_inst_dmem_n5303) );
NOR2_X1 MEM_stage_inst_dmem_U5430 ( .A1(MEM_stage_inst_dmem_n5300), .A2(MEM_stage_inst_dmem_n5299), .ZN(MEM_stage_inst_dmem_n5301) );
NAND2_X1 MEM_stage_inst_dmem_U5429 ( .A1(MEM_stage_inst_dmem_n5298), .A2(MEM_stage_inst_dmem_n5297), .ZN(MEM_stage_inst_dmem_n5299) );
NOR2_X1 MEM_stage_inst_dmem_U5428 ( .A1(MEM_stage_inst_dmem_n5296), .A2(MEM_stage_inst_dmem_n5295), .ZN(MEM_stage_inst_dmem_n5297) );
NAND2_X1 MEM_stage_inst_dmem_U5427 ( .A1(MEM_stage_inst_dmem_n5294), .A2(MEM_stage_inst_dmem_n5293), .ZN(MEM_stage_inst_dmem_n5295) );
NAND2_X1 MEM_stage_inst_dmem_U5426 ( .A1(MEM_stage_inst_dmem_ram_3721), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n5293) );
NAND2_X1 MEM_stage_inst_dmem_U5425 ( .A1(MEM_stage_inst_dmem_ram_3753), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n5294) );
NAND2_X1 MEM_stage_inst_dmem_U5424 ( .A1(MEM_stage_inst_dmem_n5292), .A2(MEM_stage_inst_dmem_n5291), .ZN(MEM_stage_inst_dmem_n5296) );
NAND2_X1 MEM_stage_inst_dmem_U5423 ( .A1(MEM_stage_inst_dmem_ram_3321), .A2(MEM_stage_inst_dmem_n39), .ZN(MEM_stage_inst_dmem_n5291) );
NAND2_X1 MEM_stage_inst_dmem_U5422 ( .A1(MEM_stage_inst_dmem_ram_3113), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n5292) );
NOR2_X1 MEM_stage_inst_dmem_U5421 ( .A1(MEM_stage_inst_dmem_n5290), .A2(MEM_stage_inst_dmem_n5289), .ZN(MEM_stage_inst_dmem_n5298) );
NAND2_X1 MEM_stage_inst_dmem_U5420 ( .A1(MEM_stage_inst_dmem_n5288), .A2(MEM_stage_inst_dmem_n5287), .ZN(MEM_stage_inst_dmem_n5289) );
NAND2_X1 MEM_stage_inst_dmem_U5419 ( .A1(MEM_stage_inst_dmem_ram_3353), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n5287) );
NAND2_X1 MEM_stage_inst_dmem_U5418 ( .A1(MEM_stage_inst_dmem_ram_3817), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n5288) );
NAND2_X1 MEM_stage_inst_dmem_U5417 ( .A1(MEM_stage_inst_dmem_n5286), .A2(MEM_stage_inst_dmem_n5285), .ZN(MEM_stage_inst_dmem_n5290) );
NAND2_X1 MEM_stage_inst_dmem_U5416 ( .A1(MEM_stage_inst_dmem_ram_3385), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n5285) );
NAND2_X1 MEM_stage_inst_dmem_U5415 ( .A1(MEM_stage_inst_dmem_ram_3497), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n5286) );
NAND2_X1 MEM_stage_inst_dmem_U5414 ( .A1(MEM_stage_inst_dmem_n5284), .A2(MEM_stage_inst_dmem_n5283), .ZN(MEM_stage_inst_dmem_n5300) );
NOR2_X1 MEM_stage_inst_dmem_U5413 ( .A1(MEM_stage_inst_dmem_n5282), .A2(MEM_stage_inst_dmem_n5281), .ZN(MEM_stage_inst_dmem_n5283) );
NAND2_X1 MEM_stage_inst_dmem_U5412 ( .A1(MEM_stage_inst_dmem_n5280), .A2(MEM_stage_inst_dmem_n5279), .ZN(MEM_stage_inst_dmem_n5281) );
NAND2_X1 MEM_stage_inst_dmem_U5411 ( .A1(MEM_stage_inst_dmem_ram_4073), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n5279) );
NAND2_X1 MEM_stage_inst_dmem_U5410 ( .A1(MEM_stage_inst_dmem_ram_3209), .A2(MEM_stage_inst_dmem_n61), .ZN(MEM_stage_inst_dmem_n5280) );
NAND2_X1 MEM_stage_inst_dmem_U5409 ( .A1(MEM_stage_inst_dmem_n5278), .A2(MEM_stage_inst_dmem_n5277), .ZN(MEM_stage_inst_dmem_n5282) );
NAND2_X1 MEM_stage_inst_dmem_U5408 ( .A1(MEM_stage_inst_dmem_ram_3945), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n5277) );
NAND2_X1 MEM_stage_inst_dmem_U5407 ( .A1(MEM_stage_inst_dmem_ram_3737), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n5278) );
NOR2_X1 MEM_stage_inst_dmem_U5406 ( .A1(MEM_stage_inst_dmem_n5276), .A2(MEM_stage_inst_dmem_n5275), .ZN(MEM_stage_inst_dmem_n5284) );
NAND2_X1 MEM_stage_inst_dmem_U5405 ( .A1(MEM_stage_inst_dmem_n5274), .A2(MEM_stage_inst_dmem_n5273), .ZN(MEM_stage_inst_dmem_n5275) );
NAND2_X1 MEM_stage_inst_dmem_U5404 ( .A1(MEM_stage_inst_dmem_ram_3961), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n5273) );
NAND2_X1 MEM_stage_inst_dmem_U5403 ( .A1(MEM_stage_inst_dmem_ram_3881), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n5274) );
NAND2_X1 MEM_stage_inst_dmem_U5402 ( .A1(MEM_stage_inst_dmem_n5272), .A2(MEM_stage_inst_dmem_n5271), .ZN(MEM_stage_inst_dmem_n5276) );
NAND2_X1 MEM_stage_inst_dmem_U5401 ( .A1(MEM_stage_inst_dmem_ram_3433), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n5271) );
NAND2_X1 MEM_stage_inst_dmem_U5400 ( .A1(MEM_stage_inst_dmem_ram_3977), .A2(MEM_stage_inst_dmem_n72), .ZN(MEM_stage_inst_dmem_n5272) );
NOR2_X1 MEM_stage_inst_dmem_U5399 ( .A1(MEM_stage_inst_dmem_n5270), .A2(MEM_stage_inst_dmem_n5269), .ZN(MEM_stage_inst_dmem_n5302) );
NAND2_X1 MEM_stage_inst_dmem_U5398 ( .A1(MEM_stage_inst_dmem_n5268), .A2(MEM_stage_inst_dmem_n5267), .ZN(MEM_stage_inst_dmem_n5269) );
NOR2_X1 MEM_stage_inst_dmem_U5397 ( .A1(MEM_stage_inst_dmem_n5266), .A2(MEM_stage_inst_dmem_n5265), .ZN(MEM_stage_inst_dmem_n5267) );
NAND2_X1 MEM_stage_inst_dmem_U5396 ( .A1(MEM_stage_inst_dmem_n5264), .A2(MEM_stage_inst_dmem_n5263), .ZN(MEM_stage_inst_dmem_n5265) );
NAND2_X1 MEM_stage_inst_dmem_U5395 ( .A1(MEM_stage_inst_dmem_ram_3929), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n5263) );
NAND2_X1 MEM_stage_inst_dmem_U5394 ( .A1(MEM_stage_inst_dmem_ram_3417), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n5264) );
NAND2_X1 MEM_stage_inst_dmem_U5393 ( .A1(MEM_stage_inst_dmem_n5262), .A2(MEM_stage_inst_dmem_n5261), .ZN(MEM_stage_inst_dmem_n5266) );
NAND2_X1 MEM_stage_inst_dmem_U5392 ( .A1(MEM_stage_inst_dmem_ram_3401), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n5261) );
NAND2_X1 MEM_stage_inst_dmem_U5391 ( .A1(MEM_stage_inst_dmem_ram_3241), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n5262) );
NOR2_X1 MEM_stage_inst_dmem_U5390 ( .A1(MEM_stage_inst_dmem_n5260), .A2(MEM_stage_inst_dmem_n5259), .ZN(MEM_stage_inst_dmem_n5268) );
NAND2_X1 MEM_stage_inst_dmem_U5389 ( .A1(MEM_stage_inst_dmem_n5258), .A2(MEM_stage_inst_dmem_n5257), .ZN(MEM_stage_inst_dmem_n5259) );
NAND2_X1 MEM_stage_inst_dmem_U5388 ( .A1(MEM_stage_inst_dmem_ram_3849), .A2(MEM_stage_inst_dmem_n37), .ZN(MEM_stage_inst_dmem_n5257) );
NAND2_X1 MEM_stage_inst_dmem_U5387 ( .A1(MEM_stage_inst_dmem_ram_3657), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n5258) );
NAND2_X1 MEM_stage_inst_dmem_U5386 ( .A1(MEM_stage_inst_dmem_n5256), .A2(MEM_stage_inst_dmem_n5255), .ZN(MEM_stage_inst_dmem_n5260) );
NAND2_X1 MEM_stage_inst_dmem_U5385 ( .A1(MEM_stage_inst_dmem_ram_3625), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n5255) );
NAND2_X1 MEM_stage_inst_dmem_U5384 ( .A1(MEM_stage_inst_dmem_ram_3081), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n5256) );
NAND2_X1 MEM_stage_inst_dmem_U5383 ( .A1(MEM_stage_inst_dmem_n5254), .A2(MEM_stage_inst_dmem_n5253), .ZN(MEM_stage_inst_dmem_n5270) );
NOR2_X1 MEM_stage_inst_dmem_U5382 ( .A1(MEM_stage_inst_dmem_n5252), .A2(MEM_stage_inst_dmem_n5251), .ZN(MEM_stage_inst_dmem_n5253) );
NAND2_X1 MEM_stage_inst_dmem_U5381 ( .A1(MEM_stage_inst_dmem_n5250), .A2(MEM_stage_inst_dmem_n5249), .ZN(MEM_stage_inst_dmem_n5251) );
NAND2_X1 MEM_stage_inst_dmem_U5380 ( .A1(MEM_stage_inst_dmem_ram_3273), .A2(MEM_stage_inst_dmem_n36), .ZN(MEM_stage_inst_dmem_n5249) );
NAND2_X1 MEM_stage_inst_dmem_U5379 ( .A1(MEM_stage_inst_dmem_ram_4057), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n5250) );
NAND2_X1 MEM_stage_inst_dmem_U5378 ( .A1(MEM_stage_inst_dmem_n5248), .A2(MEM_stage_inst_dmem_n5247), .ZN(MEM_stage_inst_dmem_n5252) );
NAND2_X1 MEM_stage_inst_dmem_U5377 ( .A1(MEM_stage_inst_dmem_ram_3161), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n5247) );
NAND2_X1 MEM_stage_inst_dmem_U5376 ( .A1(MEM_stage_inst_dmem_ram_3673), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n5248) );
NOR2_X1 MEM_stage_inst_dmem_U5375 ( .A1(MEM_stage_inst_dmem_n5246), .A2(MEM_stage_inst_dmem_n5245), .ZN(MEM_stage_inst_dmem_n5254) );
NAND2_X1 MEM_stage_inst_dmem_U5374 ( .A1(MEM_stage_inst_dmem_n5244), .A2(MEM_stage_inst_dmem_n5243), .ZN(MEM_stage_inst_dmem_n5245) );
NAND2_X1 MEM_stage_inst_dmem_U5373 ( .A1(MEM_stage_inst_dmem_ram_3225), .A2(MEM_stage_inst_dmem_n5807), .ZN(MEM_stage_inst_dmem_n5243) );
NAND2_X1 MEM_stage_inst_dmem_U5372 ( .A1(MEM_stage_inst_dmem_ram_3801), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n5244) );
NAND2_X1 MEM_stage_inst_dmem_U5371 ( .A1(MEM_stage_inst_dmem_n5242), .A2(MEM_stage_inst_dmem_n5241), .ZN(MEM_stage_inst_dmem_n5246) );
NAND2_X1 MEM_stage_inst_dmem_U5370 ( .A1(MEM_stage_inst_dmem_ram_3545), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n5241) );
NAND2_X1 MEM_stage_inst_dmem_U5369 ( .A1(MEM_stage_inst_dmem_ram_4009), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n5242) );
NAND2_X1 MEM_stage_inst_dmem_U5368 ( .A1(MEM_stage_inst_dmem_n5240), .A2(MEM_stage_inst_dmem_n5239), .ZN(MEM_stage_inst_dmem_n5304) );
NOR2_X1 MEM_stage_inst_dmem_U5367 ( .A1(MEM_stage_inst_dmem_n5238), .A2(MEM_stage_inst_dmem_n5237), .ZN(MEM_stage_inst_dmem_n5239) );
NAND2_X1 MEM_stage_inst_dmem_U5366 ( .A1(MEM_stage_inst_dmem_n5236), .A2(MEM_stage_inst_dmem_n5235), .ZN(MEM_stage_inst_dmem_n5237) );
NOR2_X1 MEM_stage_inst_dmem_U5365 ( .A1(MEM_stage_inst_dmem_n5234), .A2(MEM_stage_inst_dmem_n5233), .ZN(MEM_stage_inst_dmem_n5235) );
NAND2_X1 MEM_stage_inst_dmem_U5364 ( .A1(MEM_stage_inst_dmem_n5232), .A2(MEM_stage_inst_dmem_n5231), .ZN(MEM_stage_inst_dmem_n5233) );
NAND2_X1 MEM_stage_inst_dmem_U5363 ( .A1(MEM_stage_inst_dmem_ram_3785), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n5231) );
NAND2_X1 MEM_stage_inst_dmem_U5362 ( .A1(MEM_stage_inst_dmem_ram_3865), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n5232) );
NAND2_X1 MEM_stage_inst_dmem_U5361 ( .A1(MEM_stage_inst_dmem_n5230), .A2(MEM_stage_inst_dmem_n5229), .ZN(MEM_stage_inst_dmem_n5234) );
NAND2_X1 MEM_stage_inst_dmem_U5360 ( .A1(MEM_stage_inst_dmem_ram_3993), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n5229) );
NAND2_X1 MEM_stage_inst_dmem_U5359 ( .A1(MEM_stage_inst_dmem_ram_3193), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n5230) );
NOR2_X1 MEM_stage_inst_dmem_U5358 ( .A1(MEM_stage_inst_dmem_n5228), .A2(MEM_stage_inst_dmem_n5227), .ZN(MEM_stage_inst_dmem_n5236) );
NAND2_X1 MEM_stage_inst_dmem_U5357 ( .A1(MEM_stage_inst_dmem_n5226), .A2(MEM_stage_inst_dmem_n5225), .ZN(MEM_stage_inst_dmem_n5227) );
NAND2_X1 MEM_stage_inst_dmem_U5356 ( .A1(MEM_stage_inst_dmem_ram_3513), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n5225) );
NAND2_X1 MEM_stage_inst_dmem_U5355 ( .A1(MEM_stage_inst_dmem_ram_3769), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n5226) );
NAND2_X1 MEM_stage_inst_dmem_U5354 ( .A1(MEM_stage_inst_dmem_n5224), .A2(MEM_stage_inst_dmem_n5223), .ZN(MEM_stage_inst_dmem_n5228) );
NAND2_X1 MEM_stage_inst_dmem_U5353 ( .A1(MEM_stage_inst_dmem_ram_3305), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n5223) );
NAND2_X1 MEM_stage_inst_dmem_U5352 ( .A1(MEM_stage_inst_dmem_ram_3705), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n5224) );
NAND2_X1 MEM_stage_inst_dmem_U5351 ( .A1(MEM_stage_inst_dmem_n5222), .A2(MEM_stage_inst_dmem_n5221), .ZN(MEM_stage_inst_dmem_n5238) );
NOR2_X1 MEM_stage_inst_dmem_U5350 ( .A1(MEM_stage_inst_dmem_n5220), .A2(MEM_stage_inst_dmem_n5219), .ZN(MEM_stage_inst_dmem_n5221) );
NAND2_X1 MEM_stage_inst_dmem_U5349 ( .A1(MEM_stage_inst_dmem_n5218), .A2(MEM_stage_inst_dmem_n5217), .ZN(MEM_stage_inst_dmem_n5219) );
NAND2_X1 MEM_stage_inst_dmem_U5348 ( .A1(MEM_stage_inst_dmem_ram_3641), .A2(MEM_stage_inst_dmem_n41), .ZN(MEM_stage_inst_dmem_n5217) );
NAND2_X1 MEM_stage_inst_dmem_U5347 ( .A1(MEM_stage_inst_dmem_ram_4089), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n5218) );
NAND2_X1 MEM_stage_inst_dmem_U5346 ( .A1(MEM_stage_inst_dmem_n5216), .A2(MEM_stage_inst_dmem_n5215), .ZN(MEM_stage_inst_dmem_n5220) );
NAND2_X1 MEM_stage_inst_dmem_U5345 ( .A1(MEM_stage_inst_dmem_ram_3833), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n5215) );
NAND2_X1 MEM_stage_inst_dmem_U5344 ( .A1(MEM_stage_inst_dmem_ram_3609), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n5216) );
NOR2_X1 MEM_stage_inst_dmem_U5343 ( .A1(MEM_stage_inst_dmem_n5214), .A2(MEM_stage_inst_dmem_n5213), .ZN(MEM_stage_inst_dmem_n5222) );
NAND2_X1 MEM_stage_inst_dmem_U5342 ( .A1(MEM_stage_inst_dmem_n5212), .A2(MEM_stage_inst_dmem_n5211), .ZN(MEM_stage_inst_dmem_n5213) );
NAND2_X1 MEM_stage_inst_dmem_U5341 ( .A1(MEM_stage_inst_dmem_ram_3897), .A2(MEM_stage_inst_dmem_n46), .ZN(MEM_stage_inst_dmem_n5211) );
NAND2_X1 MEM_stage_inst_dmem_U5340 ( .A1(MEM_stage_inst_dmem_ram_3289), .A2(MEM_stage_inst_dmem_n51), .ZN(MEM_stage_inst_dmem_n5212) );
NAND2_X1 MEM_stage_inst_dmem_U5339 ( .A1(MEM_stage_inst_dmem_n5210), .A2(MEM_stage_inst_dmem_n5209), .ZN(MEM_stage_inst_dmem_n5214) );
NAND2_X1 MEM_stage_inst_dmem_U5338 ( .A1(MEM_stage_inst_dmem_ram_3369), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n5209) );
NAND2_X1 MEM_stage_inst_dmem_U5337 ( .A1(MEM_stage_inst_dmem_ram_3449), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n5210) );
NOR2_X1 MEM_stage_inst_dmem_U5336 ( .A1(MEM_stage_inst_dmem_n5208), .A2(MEM_stage_inst_dmem_n5207), .ZN(MEM_stage_inst_dmem_n5240) );
NAND2_X1 MEM_stage_inst_dmem_U5335 ( .A1(MEM_stage_inst_dmem_n5206), .A2(MEM_stage_inst_dmem_n5205), .ZN(MEM_stage_inst_dmem_n5207) );
NOR2_X1 MEM_stage_inst_dmem_U5334 ( .A1(MEM_stage_inst_dmem_n5204), .A2(MEM_stage_inst_dmem_n5203), .ZN(MEM_stage_inst_dmem_n5205) );
NAND2_X1 MEM_stage_inst_dmem_U5333 ( .A1(MEM_stage_inst_dmem_n5202), .A2(MEM_stage_inst_dmem_n5201), .ZN(MEM_stage_inst_dmem_n5203) );
NAND2_X1 MEM_stage_inst_dmem_U5332 ( .A1(MEM_stage_inst_dmem_ram_3129), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n5201) );
NAND2_X1 MEM_stage_inst_dmem_U5331 ( .A1(MEM_stage_inst_dmem_ram_3465), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n5202) );
NAND2_X1 MEM_stage_inst_dmem_U5330 ( .A1(MEM_stage_inst_dmem_n5200), .A2(MEM_stage_inst_dmem_n5199), .ZN(MEM_stage_inst_dmem_n5204) );
NAND2_X1 MEM_stage_inst_dmem_U5329 ( .A1(MEM_stage_inst_dmem_ram_3561), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n5199) );
NAND2_X1 MEM_stage_inst_dmem_U5328 ( .A1(MEM_stage_inst_dmem_ram_3145), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n5200) );
NOR2_X1 MEM_stage_inst_dmem_U5327 ( .A1(MEM_stage_inst_dmem_n5198), .A2(MEM_stage_inst_dmem_n5197), .ZN(MEM_stage_inst_dmem_n5206) );
NAND2_X1 MEM_stage_inst_dmem_U5326 ( .A1(MEM_stage_inst_dmem_n5196), .A2(MEM_stage_inst_dmem_n5195), .ZN(MEM_stage_inst_dmem_n5197) );
NAND2_X1 MEM_stage_inst_dmem_U5325 ( .A1(MEM_stage_inst_dmem_ram_3577), .A2(MEM_stage_inst_dmem_n64), .ZN(MEM_stage_inst_dmem_n5195) );
NAND2_X1 MEM_stage_inst_dmem_U5324 ( .A1(MEM_stage_inst_dmem_ram_3913), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n5196) );
NAND2_X1 MEM_stage_inst_dmem_U5323 ( .A1(MEM_stage_inst_dmem_n5194), .A2(MEM_stage_inst_dmem_n5193), .ZN(MEM_stage_inst_dmem_n5198) );
NAND2_X1 MEM_stage_inst_dmem_U5322 ( .A1(MEM_stage_inst_dmem_ram_3593), .A2(MEM_stage_inst_dmem_n71), .ZN(MEM_stage_inst_dmem_n5193) );
NAND2_X1 MEM_stage_inst_dmem_U5321 ( .A1(MEM_stage_inst_dmem_ram_3337), .A2(MEM_stage_inst_dmem_n7898), .ZN(MEM_stage_inst_dmem_n5194) );
NAND2_X1 MEM_stage_inst_dmem_U5320 ( .A1(MEM_stage_inst_dmem_n5192), .A2(MEM_stage_inst_dmem_n5191), .ZN(MEM_stage_inst_dmem_n5208) );
NOR2_X1 MEM_stage_inst_dmem_U5319 ( .A1(MEM_stage_inst_dmem_n5190), .A2(MEM_stage_inst_dmem_n5189), .ZN(MEM_stage_inst_dmem_n5191) );
NAND2_X1 MEM_stage_inst_dmem_U5318 ( .A1(MEM_stage_inst_dmem_n5188), .A2(MEM_stage_inst_dmem_n5187), .ZN(MEM_stage_inst_dmem_n5189) );
NAND2_X1 MEM_stage_inst_dmem_U5317 ( .A1(MEM_stage_inst_dmem_ram_4041), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n5187) );
NAND2_X1 MEM_stage_inst_dmem_U5316 ( .A1(MEM_stage_inst_dmem_ram_3689), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n5188) );
NAND2_X1 MEM_stage_inst_dmem_U5315 ( .A1(MEM_stage_inst_dmem_n5186), .A2(MEM_stage_inst_dmem_n5185), .ZN(MEM_stage_inst_dmem_n5190) );
NAND2_X1 MEM_stage_inst_dmem_U5314 ( .A1(MEM_stage_inst_dmem_ram_3481), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n5185) );
NAND2_X1 MEM_stage_inst_dmem_U5313 ( .A1(MEM_stage_inst_dmem_ram_3529), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n5186) );
NOR2_X1 MEM_stage_inst_dmem_U5312 ( .A1(MEM_stage_inst_dmem_n5184), .A2(MEM_stage_inst_dmem_n5183), .ZN(MEM_stage_inst_dmem_n5192) );
NAND2_X1 MEM_stage_inst_dmem_U5311 ( .A1(MEM_stage_inst_dmem_n5182), .A2(MEM_stage_inst_dmem_n5181), .ZN(MEM_stage_inst_dmem_n5183) );
NAND2_X1 MEM_stage_inst_dmem_U5310 ( .A1(MEM_stage_inst_dmem_ram_4025), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n5181) );
NAND2_X1 MEM_stage_inst_dmem_U5309 ( .A1(MEM_stage_inst_dmem_ram_3097), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n5182) );
NAND2_X1 MEM_stage_inst_dmem_U5308 ( .A1(MEM_stage_inst_dmem_n5180), .A2(MEM_stage_inst_dmem_n5179), .ZN(MEM_stage_inst_dmem_n5184) );
NAND2_X1 MEM_stage_inst_dmem_U5307 ( .A1(MEM_stage_inst_dmem_ram_3257), .A2(MEM_stage_inst_dmem_n55), .ZN(MEM_stage_inst_dmem_n5179) );
NAND2_X1 MEM_stage_inst_dmem_U5306 ( .A1(MEM_stage_inst_dmem_ram_3177), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n5180) );
NOR2_X1 MEM_stage_inst_dmem_U5305 ( .A1(MEM_stage_inst_dmem_n5178), .A2(MEM_stage_inst_dmem_n5177), .ZN(MEM_stage_inst_dmem_n5436) );
NOR2_X1 MEM_stage_inst_dmem_U5304 ( .A1(MEM_stage_inst_dmem_n5176), .A2(MEM_stage_inst_dmem_n8286), .ZN(MEM_stage_inst_dmem_n5177) );
NOR2_X1 MEM_stage_inst_dmem_U5303 ( .A1(MEM_stage_inst_dmem_n5175), .A2(MEM_stage_inst_dmem_n5174), .ZN(MEM_stage_inst_dmem_n5176) );
NAND2_X1 MEM_stage_inst_dmem_U5302 ( .A1(MEM_stage_inst_dmem_n5173), .A2(MEM_stage_inst_dmem_n5172), .ZN(MEM_stage_inst_dmem_n5174) );
NOR2_X1 MEM_stage_inst_dmem_U5301 ( .A1(MEM_stage_inst_dmem_n5171), .A2(MEM_stage_inst_dmem_n5170), .ZN(MEM_stage_inst_dmem_n5172) );
NAND2_X1 MEM_stage_inst_dmem_U5300 ( .A1(MEM_stage_inst_dmem_n5169), .A2(MEM_stage_inst_dmem_n5168), .ZN(MEM_stage_inst_dmem_n5170) );
NOR2_X1 MEM_stage_inst_dmem_U5299 ( .A1(MEM_stage_inst_dmem_n5167), .A2(MEM_stage_inst_dmem_n5166), .ZN(MEM_stage_inst_dmem_n5168) );
NAND2_X1 MEM_stage_inst_dmem_U5298 ( .A1(MEM_stage_inst_dmem_n5165), .A2(MEM_stage_inst_dmem_n5164), .ZN(MEM_stage_inst_dmem_n5166) );
NAND2_X1 MEM_stage_inst_dmem_U5297 ( .A1(MEM_stage_inst_dmem_ram_2473), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n5164) );
NAND2_X1 MEM_stage_inst_dmem_U5296 ( .A1(MEM_stage_inst_dmem_ram_2681), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n5165) );
NAND2_X1 MEM_stage_inst_dmem_U5295 ( .A1(MEM_stage_inst_dmem_n5163), .A2(MEM_stage_inst_dmem_n5162), .ZN(MEM_stage_inst_dmem_n5167) );
NAND2_X1 MEM_stage_inst_dmem_U5294 ( .A1(MEM_stage_inst_dmem_ram_2937), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n5162) );
NAND2_X1 MEM_stage_inst_dmem_U5293 ( .A1(MEM_stage_inst_dmem_ram_2505), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n5163) );
NOR2_X1 MEM_stage_inst_dmem_U5292 ( .A1(MEM_stage_inst_dmem_n5161), .A2(MEM_stage_inst_dmem_n5160), .ZN(MEM_stage_inst_dmem_n5169) );
NAND2_X1 MEM_stage_inst_dmem_U5291 ( .A1(MEM_stage_inst_dmem_n5159), .A2(MEM_stage_inst_dmem_n5158), .ZN(MEM_stage_inst_dmem_n5160) );
NAND2_X1 MEM_stage_inst_dmem_U5290 ( .A1(MEM_stage_inst_dmem_ram_2345), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n5158) );
NAND2_X1 MEM_stage_inst_dmem_U5289 ( .A1(MEM_stage_inst_dmem_ram_2393), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n5159) );
NAND2_X1 MEM_stage_inst_dmem_U5288 ( .A1(MEM_stage_inst_dmem_n5157), .A2(MEM_stage_inst_dmem_n5156), .ZN(MEM_stage_inst_dmem_n5161) );
NAND2_X1 MEM_stage_inst_dmem_U5287 ( .A1(MEM_stage_inst_dmem_ram_2377), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n5156) );
NAND2_X1 MEM_stage_inst_dmem_U5286 ( .A1(MEM_stage_inst_dmem_ram_2441), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n5157) );
NAND2_X1 MEM_stage_inst_dmem_U5285 ( .A1(MEM_stage_inst_dmem_n5155), .A2(MEM_stage_inst_dmem_n5154), .ZN(MEM_stage_inst_dmem_n5171) );
NOR2_X1 MEM_stage_inst_dmem_U5284 ( .A1(MEM_stage_inst_dmem_n5153), .A2(MEM_stage_inst_dmem_n5152), .ZN(MEM_stage_inst_dmem_n5154) );
NAND2_X1 MEM_stage_inst_dmem_U5283 ( .A1(MEM_stage_inst_dmem_n5151), .A2(MEM_stage_inst_dmem_n5150), .ZN(MEM_stage_inst_dmem_n5152) );
NAND2_X1 MEM_stage_inst_dmem_U5282 ( .A1(MEM_stage_inst_dmem_ram_3065), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n5150) );
NAND2_X1 MEM_stage_inst_dmem_U5281 ( .A1(MEM_stage_inst_dmem_ram_2313), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n5151) );
NAND2_X1 MEM_stage_inst_dmem_U5280 ( .A1(MEM_stage_inst_dmem_n5149), .A2(MEM_stage_inst_dmem_n5148), .ZN(MEM_stage_inst_dmem_n5153) );
NAND2_X1 MEM_stage_inst_dmem_U5279 ( .A1(MEM_stage_inst_dmem_ram_2361), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n5148) );
NAND2_X1 MEM_stage_inst_dmem_U5278 ( .A1(MEM_stage_inst_dmem_ram_2073), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n5149) );
NOR2_X1 MEM_stage_inst_dmem_U5277 ( .A1(MEM_stage_inst_dmem_n5147), .A2(MEM_stage_inst_dmem_n5146), .ZN(MEM_stage_inst_dmem_n5155) );
NAND2_X1 MEM_stage_inst_dmem_U5276 ( .A1(MEM_stage_inst_dmem_n5145), .A2(MEM_stage_inst_dmem_n5144), .ZN(MEM_stage_inst_dmem_n5146) );
NAND2_X1 MEM_stage_inst_dmem_U5275 ( .A1(MEM_stage_inst_dmem_ram_2089), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n5144) );
NAND2_X1 MEM_stage_inst_dmem_U5274 ( .A1(MEM_stage_inst_dmem_ram_2729), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n5145) );
NAND2_X1 MEM_stage_inst_dmem_U5273 ( .A1(MEM_stage_inst_dmem_n5143), .A2(MEM_stage_inst_dmem_n5142), .ZN(MEM_stage_inst_dmem_n5147) );
NAND2_X1 MEM_stage_inst_dmem_U5272 ( .A1(MEM_stage_inst_dmem_ram_2761), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n5142) );
NAND2_X1 MEM_stage_inst_dmem_U5271 ( .A1(MEM_stage_inst_dmem_ram_2217), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n5143) );
NOR2_X1 MEM_stage_inst_dmem_U5270 ( .A1(MEM_stage_inst_dmem_n5141), .A2(MEM_stage_inst_dmem_n5140), .ZN(MEM_stage_inst_dmem_n5173) );
NAND2_X1 MEM_stage_inst_dmem_U5269 ( .A1(MEM_stage_inst_dmem_n5139), .A2(MEM_stage_inst_dmem_n5138), .ZN(MEM_stage_inst_dmem_n5140) );
NOR2_X1 MEM_stage_inst_dmem_U5268 ( .A1(MEM_stage_inst_dmem_n5137), .A2(MEM_stage_inst_dmem_n5136), .ZN(MEM_stage_inst_dmem_n5138) );
NAND2_X1 MEM_stage_inst_dmem_U5267 ( .A1(MEM_stage_inst_dmem_n5135), .A2(MEM_stage_inst_dmem_n5134), .ZN(MEM_stage_inst_dmem_n5136) );
NAND2_X1 MEM_stage_inst_dmem_U5266 ( .A1(MEM_stage_inst_dmem_ram_2889), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n5134) );
NAND2_X1 MEM_stage_inst_dmem_U5265 ( .A1(MEM_stage_inst_dmem_ram_2713), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n5135) );
NAND2_X1 MEM_stage_inst_dmem_U5264 ( .A1(MEM_stage_inst_dmem_n5133), .A2(MEM_stage_inst_dmem_n5132), .ZN(MEM_stage_inst_dmem_n5137) );
NAND2_X1 MEM_stage_inst_dmem_U5263 ( .A1(MEM_stage_inst_dmem_ram_2617), .A2(MEM_stage_inst_dmem_n41), .ZN(MEM_stage_inst_dmem_n5132) );
NAND2_X1 MEM_stage_inst_dmem_U5262 ( .A1(MEM_stage_inst_dmem_ram_2569), .A2(MEM_stage_inst_dmem_n71), .ZN(MEM_stage_inst_dmem_n5133) );
NOR2_X1 MEM_stage_inst_dmem_U5261 ( .A1(MEM_stage_inst_dmem_n5131), .A2(MEM_stage_inst_dmem_n5130), .ZN(MEM_stage_inst_dmem_n5139) );
NAND2_X1 MEM_stage_inst_dmem_U5260 ( .A1(MEM_stage_inst_dmem_n5129), .A2(MEM_stage_inst_dmem_n5128), .ZN(MEM_stage_inst_dmem_n5130) );
NAND2_X1 MEM_stage_inst_dmem_U5259 ( .A1(MEM_stage_inst_dmem_ram_2601), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n5128) );
NAND2_X1 MEM_stage_inst_dmem_U5258 ( .A1(MEM_stage_inst_dmem_ram_2857), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n5129) );
NAND2_X1 MEM_stage_inst_dmem_U5257 ( .A1(MEM_stage_inst_dmem_n5127), .A2(MEM_stage_inst_dmem_n5126), .ZN(MEM_stage_inst_dmem_n5131) );
NAND2_X1 MEM_stage_inst_dmem_U5256 ( .A1(MEM_stage_inst_dmem_ram_2409), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n5126) );
NAND2_X1 MEM_stage_inst_dmem_U5255 ( .A1(MEM_stage_inst_dmem_ram_2457), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n5127) );
NAND2_X1 MEM_stage_inst_dmem_U5254 ( .A1(MEM_stage_inst_dmem_n5125), .A2(MEM_stage_inst_dmem_n5124), .ZN(MEM_stage_inst_dmem_n5141) );
NOR2_X1 MEM_stage_inst_dmem_U5253 ( .A1(MEM_stage_inst_dmem_n5123), .A2(MEM_stage_inst_dmem_n5122), .ZN(MEM_stage_inst_dmem_n5124) );
NAND2_X1 MEM_stage_inst_dmem_U5252 ( .A1(MEM_stage_inst_dmem_n5121), .A2(MEM_stage_inst_dmem_n5120), .ZN(MEM_stage_inst_dmem_n5122) );
NAND2_X1 MEM_stage_inst_dmem_U5251 ( .A1(MEM_stage_inst_dmem_ram_3001), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n5120) );
NAND2_X1 MEM_stage_inst_dmem_U5250 ( .A1(MEM_stage_inst_dmem_ram_2953), .A2(MEM_stage_inst_dmem_n72), .ZN(MEM_stage_inst_dmem_n5121) );
NAND2_X1 MEM_stage_inst_dmem_U5249 ( .A1(MEM_stage_inst_dmem_n5119), .A2(MEM_stage_inst_dmem_n5118), .ZN(MEM_stage_inst_dmem_n5123) );
NAND2_X1 MEM_stage_inst_dmem_U5248 ( .A1(MEM_stage_inst_dmem_ram_2873), .A2(MEM_stage_inst_dmem_n46), .ZN(MEM_stage_inst_dmem_n5118) );
NAND2_X1 MEM_stage_inst_dmem_U5247 ( .A1(MEM_stage_inst_dmem_ram_2425), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n5119) );
NOR2_X1 MEM_stage_inst_dmem_U5246 ( .A1(MEM_stage_inst_dmem_n5117), .A2(MEM_stage_inst_dmem_n5116), .ZN(MEM_stage_inst_dmem_n5125) );
NAND2_X1 MEM_stage_inst_dmem_U5245 ( .A1(MEM_stage_inst_dmem_n5115), .A2(MEM_stage_inst_dmem_n5114), .ZN(MEM_stage_inst_dmem_n5116) );
NAND2_X1 MEM_stage_inst_dmem_U5244 ( .A1(MEM_stage_inst_dmem_ram_3017), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n5114) );
NAND2_X1 MEM_stage_inst_dmem_U5243 ( .A1(MEM_stage_inst_dmem_ram_2057), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n5115) );
NAND2_X1 MEM_stage_inst_dmem_U5242 ( .A1(MEM_stage_inst_dmem_n5113), .A2(MEM_stage_inst_dmem_n5112), .ZN(MEM_stage_inst_dmem_n5117) );
NAND2_X1 MEM_stage_inst_dmem_U5241 ( .A1(MEM_stage_inst_dmem_ram_2969), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n5112) );
NAND2_X1 MEM_stage_inst_dmem_U5240 ( .A1(MEM_stage_inst_dmem_ram_2649), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n5113) );
NAND2_X1 MEM_stage_inst_dmem_U5239 ( .A1(MEM_stage_inst_dmem_n5111), .A2(MEM_stage_inst_dmem_n5110), .ZN(MEM_stage_inst_dmem_n5175) );
NOR2_X1 MEM_stage_inst_dmem_U5238 ( .A1(MEM_stage_inst_dmem_n5109), .A2(MEM_stage_inst_dmem_n5108), .ZN(MEM_stage_inst_dmem_n5110) );
NAND2_X1 MEM_stage_inst_dmem_U5237 ( .A1(MEM_stage_inst_dmem_n5107), .A2(MEM_stage_inst_dmem_n5106), .ZN(MEM_stage_inst_dmem_n5108) );
NOR2_X1 MEM_stage_inst_dmem_U5236 ( .A1(MEM_stage_inst_dmem_n5105), .A2(MEM_stage_inst_dmem_n5104), .ZN(MEM_stage_inst_dmem_n5106) );
NAND2_X1 MEM_stage_inst_dmem_U5235 ( .A1(MEM_stage_inst_dmem_n5103), .A2(MEM_stage_inst_dmem_n5102), .ZN(MEM_stage_inst_dmem_n5104) );
NAND2_X1 MEM_stage_inst_dmem_U5234 ( .A1(MEM_stage_inst_dmem_ram_2841), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n5102) );
NAND2_X1 MEM_stage_inst_dmem_U5233 ( .A1(MEM_stage_inst_dmem_ram_2585), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n5103) );
NAND2_X1 MEM_stage_inst_dmem_U5232 ( .A1(MEM_stage_inst_dmem_n5101), .A2(MEM_stage_inst_dmem_n5100), .ZN(MEM_stage_inst_dmem_n5105) );
NAND2_X1 MEM_stage_inst_dmem_U5231 ( .A1(MEM_stage_inst_dmem_ram_2537), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n5100) );
NAND2_X1 MEM_stage_inst_dmem_U5230 ( .A1(MEM_stage_inst_dmem_ram_2777), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n5101) );
NOR2_X1 MEM_stage_inst_dmem_U5229 ( .A1(MEM_stage_inst_dmem_n5099), .A2(MEM_stage_inst_dmem_n5098), .ZN(MEM_stage_inst_dmem_n5107) );
NAND2_X1 MEM_stage_inst_dmem_U5228 ( .A1(MEM_stage_inst_dmem_n5097), .A2(MEM_stage_inst_dmem_n5096), .ZN(MEM_stage_inst_dmem_n5098) );
NAND2_X1 MEM_stage_inst_dmem_U5227 ( .A1(MEM_stage_inst_dmem_ram_2249), .A2(MEM_stage_inst_dmem_n36), .ZN(MEM_stage_inst_dmem_n5096) );
NAND2_X1 MEM_stage_inst_dmem_U5226 ( .A1(MEM_stage_inst_dmem_ram_2697), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n5097) );
NAND2_X1 MEM_stage_inst_dmem_U5225 ( .A1(MEM_stage_inst_dmem_n5095), .A2(MEM_stage_inst_dmem_n5094), .ZN(MEM_stage_inst_dmem_n5099) );
NAND2_X1 MEM_stage_inst_dmem_U5224 ( .A1(MEM_stage_inst_dmem_ram_2169), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n5094) );
NAND2_X1 MEM_stage_inst_dmem_U5223 ( .A1(MEM_stage_inst_dmem_ram_2153), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n5095) );
NAND2_X1 MEM_stage_inst_dmem_U5222 ( .A1(MEM_stage_inst_dmem_n5093), .A2(MEM_stage_inst_dmem_n5092), .ZN(MEM_stage_inst_dmem_n5109) );
NOR2_X1 MEM_stage_inst_dmem_U5221 ( .A1(MEM_stage_inst_dmem_n5091), .A2(MEM_stage_inst_dmem_n5090), .ZN(MEM_stage_inst_dmem_n5092) );
NAND2_X1 MEM_stage_inst_dmem_U5220 ( .A1(MEM_stage_inst_dmem_n5089), .A2(MEM_stage_inst_dmem_n5088), .ZN(MEM_stage_inst_dmem_n5090) );
NAND2_X1 MEM_stage_inst_dmem_U5219 ( .A1(MEM_stage_inst_dmem_ram_2825), .A2(MEM_stage_inst_dmem_n8472), .ZN(MEM_stage_inst_dmem_n5088) );
NAND2_X1 MEM_stage_inst_dmem_U5218 ( .A1(MEM_stage_inst_dmem_ram_2665), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n5089) );
NAND2_X1 MEM_stage_inst_dmem_U5217 ( .A1(MEM_stage_inst_dmem_n5087), .A2(MEM_stage_inst_dmem_n5086), .ZN(MEM_stage_inst_dmem_n5091) );
NAND2_X1 MEM_stage_inst_dmem_U5216 ( .A1(MEM_stage_inst_dmem_ram_2105), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n5086) );
NAND2_X1 MEM_stage_inst_dmem_U5215 ( .A1(MEM_stage_inst_dmem_ram_2185), .A2(MEM_stage_inst_dmem_n61), .ZN(MEM_stage_inst_dmem_n5087) );
NOR2_X1 MEM_stage_inst_dmem_U5214 ( .A1(MEM_stage_inst_dmem_n5085), .A2(MEM_stage_inst_dmem_n5084), .ZN(MEM_stage_inst_dmem_n5093) );
NAND2_X1 MEM_stage_inst_dmem_U5213 ( .A1(MEM_stage_inst_dmem_n5083), .A2(MEM_stage_inst_dmem_n5082), .ZN(MEM_stage_inst_dmem_n5084) );
NAND2_X1 MEM_stage_inst_dmem_U5212 ( .A1(MEM_stage_inst_dmem_ram_3049), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n5082) );
NAND2_X1 MEM_stage_inst_dmem_U5211 ( .A1(MEM_stage_inst_dmem_ram_2633), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n5083) );
NAND2_X1 MEM_stage_inst_dmem_U5210 ( .A1(MEM_stage_inst_dmem_n5081), .A2(MEM_stage_inst_dmem_n5080), .ZN(MEM_stage_inst_dmem_n5085) );
NAND2_X1 MEM_stage_inst_dmem_U5209 ( .A1(MEM_stage_inst_dmem_ram_3033), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n5080) );
NAND2_X1 MEM_stage_inst_dmem_U5208 ( .A1(MEM_stage_inst_dmem_ram_2201), .A2(MEM_stage_inst_dmem_n44), .ZN(MEM_stage_inst_dmem_n5081) );
NOR2_X1 MEM_stage_inst_dmem_U5207 ( .A1(MEM_stage_inst_dmem_n5079), .A2(MEM_stage_inst_dmem_n5078), .ZN(MEM_stage_inst_dmem_n5111) );
NAND2_X1 MEM_stage_inst_dmem_U5206 ( .A1(MEM_stage_inst_dmem_n5077), .A2(MEM_stage_inst_dmem_n5076), .ZN(MEM_stage_inst_dmem_n5078) );
NOR2_X1 MEM_stage_inst_dmem_U5205 ( .A1(MEM_stage_inst_dmem_n5075), .A2(MEM_stage_inst_dmem_n5074), .ZN(MEM_stage_inst_dmem_n5076) );
NAND2_X1 MEM_stage_inst_dmem_U5204 ( .A1(MEM_stage_inst_dmem_n5073), .A2(MEM_stage_inst_dmem_n5072), .ZN(MEM_stage_inst_dmem_n5074) );
NAND2_X1 MEM_stage_inst_dmem_U5203 ( .A1(MEM_stage_inst_dmem_ram_2921), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n5072) );
NAND2_X1 MEM_stage_inst_dmem_U5202 ( .A1(MEM_stage_inst_dmem_ram_2985), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n5073) );
NAND2_X1 MEM_stage_inst_dmem_U5201 ( .A1(MEM_stage_inst_dmem_n5071), .A2(MEM_stage_inst_dmem_n5070), .ZN(MEM_stage_inst_dmem_n5075) );
NAND2_X1 MEM_stage_inst_dmem_U5200 ( .A1(MEM_stage_inst_dmem_ram_2281), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n5070) );
NAND2_X1 MEM_stage_inst_dmem_U5199 ( .A1(MEM_stage_inst_dmem_ram_2233), .A2(MEM_stage_inst_dmem_n8434), .ZN(MEM_stage_inst_dmem_n5071) );
NOR2_X1 MEM_stage_inst_dmem_U5198 ( .A1(MEM_stage_inst_dmem_n5069), .A2(MEM_stage_inst_dmem_n5068), .ZN(MEM_stage_inst_dmem_n5077) );
NAND2_X1 MEM_stage_inst_dmem_U5197 ( .A1(MEM_stage_inst_dmem_n5067), .A2(MEM_stage_inst_dmem_n5066), .ZN(MEM_stage_inst_dmem_n5068) );
NAND2_X1 MEM_stage_inst_dmem_U5196 ( .A1(MEM_stage_inst_dmem_ram_2905), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n5066) );
NAND2_X1 MEM_stage_inst_dmem_U5195 ( .A1(MEM_stage_inst_dmem_ram_2329), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n5067) );
NAND2_X1 MEM_stage_inst_dmem_U5194 ( .A1(MEM_stage_inst_dmem_n5065), .A2(MEM_stage_inst_dmem_n5064), .ZN(MEM_stage_inst_dmem_n5069) );
NAND2_X1 MEM_stage_inst_dmem_U5193 ( .A1(MEM_stage_inst_dmem_ram_2553), .A2(MEM_stage_inst_dmem_n64), .ZN(MEM_stage_inst_dmem_n5064) );
NAND2_X1 MEM_stage_inst_dmem_U5192 ( .A1(MEM_stage_inst_dmem_ram_2809), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n5065) );
NAND2_X1 MEM_stage_inst_dmem_U5191 ( .A1(MEM_stage_inst_dmem_n5063), .A2(MEM_stage_inst_dmem_n5062), .ZN(MEM_stage_inst_dmem_n5079) );
NOR2_X1 MEM_stage_inst_dmem_U5190 ( .A1(MEM_stage_inst_dmem_n5061), .A2(MEM_stage_inst_dmem_n5060), .ZN(MEM_stage_inst_dmem_n5062) );
NAND2_X1 MEM_stage_inst_dmem_U5189 ( .A1(MEM_stage_inst_dmem_n5059), .A2(MEM_stage_inst_dmem_n5058), .ZN(MEM_stage_inst_dmem_n5060) );
NAND2_X1 MEM_stage_inst_dmem_U5188 ( .A1(MEM_stage_inst_dmem_ram_2745), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n5058) );
NAND2_X1 MEM_stage_inst_dmem_U5187 ( .A1(MEM_stage_inst_dmem_ram_2793), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n5059) );
NAND2_X1 MEM_stage_inst_dmem_U5186 ( .A1(MEM_stage_inst_dmem_n5057), .A2(MEM_stage_inst_dmem_n5056), .ZN(MEM_stage_inst_dmem_n5061) );
NAND2_X1 MEM_stage_inst_dmem_U5185 ( .A1(MEM_stage_inst_dmem_ram_2137), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n5056) );
NAND2_X1 MEM_stage_inst_dmem_U5184 ( .A1(MEM_stage_inst_dmem_ram_2521), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n5057) );
NOR2_X1 MEM_stage_inst_dmem_U5183 ( .A1(MEM_stage_inst_dmem_n5055), .A2(MEM_stage_inst_dmem_n5054), .ZN(MEM_stage_inst_dmem_n5063) );
NAND2_X1 MEM_stage_inst_dmem_U5182 ( .A1(MEM_stage_inst_dmem_n5053), .A2(MEM_stage_inst_dmem_n5052), .ZN(MEM_stage_inst_dmem_n5054) );
NAND2_X1 MEM_stage_inst_dmem_U5181 ( .A1(MEM_stage_inst_dmem_ram_2489), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n5052) );
NAND2_X1 MEM_stage_inst_dmem_U5180 ( .A1(MEM_stage_inst_dmem_ram_2121), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n5053) );
NAND2_X1 MEM_stage_inst_dmem_U5179 ( .A1(MEM_stage_inst_dmem_n5051), .A2(MEM_stage_inst_dmem_n5050), .ZN(MEM_stage_inst_dmem_n5055) );
NAND2_X1 MEM_stage_inst_dmem_U5178 ( .A1(MEM_stage_inst_dmem_ram_2297), .A2(MEM_stage_inst_dmem_n39), .ZN(MEM_stage_inst_dmem_n5050) );
NAND2_X1 MEM_stage_inst_dmem_U5177 ( .A1(MEM_stage_inst_dmem_ram_2265), .A2(MEM_stage_inst_dmem_n51), .ZN(MEM_stage_inst_dmem_n5051) );
NOR2_X1 MEM_stage_inst_dmem_U5176 ( .A1(MEM_stage_inst_dmem_n5049), .A2(MEM_stage_inst_dmem_n8152), .ZN(MEM_stage_inst_dmem_n5178) );
NOR2_X1 MEM_stage_inst_dmem_U5175 ( .A1(MEM_stage_inst_dmem_n5048), .A2(MEM_stage_inst_dmem_n5047), .ZN(MEM_stage_inst_dmem_n5049) );
NAND2_X1 MEM_stage_inst_dmem_U5174 ( .A1(MEM_stage_inst_dmem_n5046), .A2(MEM_stage_inst_dmem_n5045), .ZN(MEM_stage_inst_dmem_n5047) );
NOR2_X1 MEM_stage_inst_dmem_U5173 ( .A1(MEM_stage_inst_dmem_n5044), .A2(MEM_stage_inst_dmem_n5043), .ZN(MEM_stage_inst_dmem_n5045) );
NAND2_X1 MEM_stage_inst_dmem_U5172 ( .A1(MEM_stage_inst_dmem_n5042), .A2(MEM_stage_inst_dmem_n5041), .ZN(MEM_stage_inst_dmem_n5043) );
NOR2_X1 MEM_stage_inst_dmem_U5171 ( .A1(MEM_stage_inst_dmem_n5040), .A2(MEM_stage_inst_dmem_n5039), .ZN(MEM_stage_inst_dmem_n5041) );
NAND2_X1 MEM_stage_inst_dmem_U5170 ( .A1(MEM_stage_inst_dmem_n5038), .A2(MEM_stage_inst_dmem_n5037), .ZN(MEM_stage_inst_dmem_n5039) );
NAND2_X1 MEM_stage_inst_dmem_U5169 ( .A1(MEM_stage_inst_dmem_ram_1273), .A2(MEM_stage_inst_dmem_n39), .ZN(MEM_stage_inst_dmem_n5037) );
NAND2_X1 MEM_stage_inst_dmem_U5168 ( .A1(MEM_stage_inst_dmem_ram_1545), .A2(MEM_stage_inst_dmem_n71), .ZN(MEM_stage_inst_dmem_n5038) );
NAND2_X1 MEM_stage_inst_dmem_U5167 ( .A1(MEM_stage_inst_dmem_n5036), .A2(MEM_stage_inst_dmem_n5035), .ZN(MEM_stage_inst_dmem_n5040) );
NAND2_X1 MEM_stage_inst_dmem_U5166 ( .A1(MEM_stage_inst_dmem_ram_1801), .A2(MEM_stage_inst_dmem_n7992), .ZN(MEM_stage_inst_dmem_n5035) );
NAND2_X1 MEM_stage_inst_dmem_U5165 ( .A1(MEM_stage_inst_dmem_ram_1977), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n5036) );
NOR2_X1 MEM_stage_inst_dmem_U5164 ( .A1(MEM_stage_inst_dmem_n5034), .A2(MEM_stage_inst_dmem_n5033), .ZN(MEM_stage_inst_dmem_n5042) );
NAND2_X1 MEM_stage_inst_dmem_U5163 ( .A1(MEM_stage_inst_dmem_n5032), .A2(MEM_stage_inst_dmem_n5031), .ZN(MEM_stage_inst_dmem_n5033) );
NAND2_X1 MEM_stage_inst_dmem_U5162 ( .A1(MEM_stage_inst_dmem_ram_1049), .A2(MEM_stage_inst_dmem_n7887), .ZN(MEM_stage_inst_dmem_n5031) );
NAND2_X1 MEM_stage_inst_dmem_U5161 ( .A1(MEM_stage_inst_dmem_ram_1241), .A2(MEM_stage_inst_dmem_n51), .ZN(MEM_stage_inst_dmem_n5032) );
NAND2_X1 MEM_stage_inst_dmem_U5160 ( .A1(MEM_stage_inst_dmem_n5030), .A2(MEM_stage_inst_dmem_n5029), .ZN(MEM_stage_inst_dmem_n5034) );
NAND2_X1 MEM_stage_inst_dmem_U5159 ( .A1(MEM_stage_inst_dmem_ram_1209), .A2(MEM_stage_inst_dmem_n7937), .ZN(MEM_stage_inst_dmem_n5029) );
NAND2_X1 MEM_stage_inst_dmem_U5158 ( .A1(MEM_stage_inst_dmem_ram_1401), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n5030) );
NAND2_X1 MEM_stage_inst_dmem_U5157 ( .A1(MEM_stage_inst_dmem_n5028), .A2(MEM_stage_inst_dmem_n5027), .ZN(MEM_stage_inst_dmem_n5044) );
NOR2_X1 MEM_stage_inst_dmem_U5156 ( .A1(MEM_stage_inst_dmem_n5026), .A2(MEM_stage_inst_dmem_n5025), .ZN(MEM_stage_inst_dmem_n5027) );
NAND2_X1 MEM_stage_inst_dmem_U5155 ( .A1(MEM_stage_inst_dmem_n5024), .A2(MEM_stage_inst_dmem_n5023), .ZN(MEM_stage_inst_dmem_n5025) );
NAND2_X1 MEM_stage_inst_dmem_U5154 ( .A1(MEM_stage_inst_dmem_ram_1673), .A2(MEM_stage_inst_dmem_n7960), .ZN(MEM_stage_inst_dmem_n5023) );
NAND2_X1 MEM_stage_inst_dmem_U5153 ( .A1(MEM_stage_inst_dmem_ram_2041), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n5024) );
NAND2_X1 MEM_stage_inst_dmem_U5152 ( .A1(MEM_stage_inst_dmem_n5022), .A2(MEM_stage_inst_dmem_n5021), .ZN(MEM_stage_inst_dmem_n5026) );
NAND2_X1 MEM_stage_inst_dmem_U5151 ( .A1(MEM_stage_inst_dmem_ram_1929), .A2(MEM_stage_inst_dmem_n72), .ZN(MEM_stage_inst_dmem_n5021) );
NAND2_X1 MEM_stage_inst_dmem_U5150 ( .A1(MEM_stage_inst_dmem_ram_1657), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n5022) );
NOR2_X1 MEM_stage_inst_dmem_U5149 ( .A1(MEM_stage_inst_dmem_n5020), .A2(MEM_stage_inst_dmem_n5019), .ZN(MEM_stage_inst_dmem_n5028) );
NAND2_X1 MEM_stage_inst_dmem_U5148 ( .A1(MEM_stage_inst_dmem_n5018), .A2(MEM_stage_inst_dmem_n5017), .ZN(MEM_stage_inst_dmem_n5019) );
NAND2_X1 MEM_stage_inst_dmem_U5147 ( .A1(MEM_stage_inst_dmem_ram_1257), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n5017) );
NAND2_X1 MEM_stage_inst_dmem_U5146 ( .A1(MEM_stage_inst_dmem_ram_1321), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n5018) );
NAND2_X1 MEM_stage_inst_dmem_U5145 ( .A1(MEM_stage_inst_dmem_n5016), .A2(MEM_stage_inst_dmem_n5015), .ZN(MEM_stage_inst_dmem_n5020) );
NAND2_X1 MEM_stage_inst_dmem_U5144 ( .A1(MEM_stage_inst_dmem_ram_1465), .A2(MEM_stage_inst_dmem_n7888), .ZN(MEM_stage_inst_dmem_n5015) );
NAND2_X1 MEM_stage_inst_dmem_U5143 ( .A1(MEM_stage_inst_dmem_ram_1641), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n5016) );
NOR2_X1 MEM_stage_inst_dmem_U5142 ( .A1(MEM_stage_inst_dmem_n5014), .A2(MEM_stage_inst_dmem_n5013), .ZN(MEM_stage_inst_dmem_n5046) );
NAND2_X1 MEM_stage_inst_dmem_U5141 ( .A1(MEM_stage_inst_dmem_n5012), .A2(MEM_stage_inst_dmem_n5011), .ZN(MEM_stage_inst_dmem_n5013) );
NOR2_X1 MEM_stage_inst_dmem_U5140 ( .A1(MEM_stage_inst_dmem_n5010), .A2(MEM_stage_inst_dmem_n5009), .ZN(MEM_stage_inst_dmem_n5011) );
NAND2_X1 MEM_stage_inst_dmem_U5139 ( .A1(MEM_stage_inst_dmem_n5008), .A2(MEM_stage_inst_dmem_n5007), .ZN(MEM_stage_inst_dmem_n5009) );
NAND2_X1 MEM_stage_inst_dmem_U5138 ( .A1(MEM_stage_inst_dmem_ram_1913), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n5007) );
NAND2_X1 MEM_stage_inst_dmem_U5137 ( .A1(MEM_stage_inst_dmem_ram_1849), .A2(MEM_stage_inst_dmem_n46), .ZN(MEM_stage_inst_dmem_n5008) );
NAND2_X1 MEM_stage_inst_dmem_U5136 ( .A1(MEM_stage_inst_dmem_n5006), .A2(MEM_stage_inst_dmem_n5005), .ZN(MEM_stage_inst_dmem_n5010) );
NAND2_X1 MEM_stage_inst_dmem_U5135 ( .A1(MEM_stage_inst_dmem_ram_1433), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n5005) );
NAND2_X1 MEM_stage_inst_dmem_U5134 ( .A1(MEM_stage_inst_dmem_ram_1833), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n5006) );
NOR2_X1 MEM_stage_inst_dmem_U5133 ( .A1(MEM_stage_inst_dmem_n5004), .A2(MEM_stage_inst_dmem_n5003), .ZN(MEM_stage_inst_dmem_n5012) );
NAND2_X1 MEM_stage_inst_dmem_U5132 ( .A1(MEM_stage_inst_dmem_n5002), .A2(MEM_stage_inst_dmem_n5001), .ZN(MEM_stage_inst_dmem_n5003) );
NAND2_X1 MEM_stage_inst_dmem_U5131 ( .A1(MEM_stage_inst_dmem_ram_2009), .A2(MEM_stage_inst_dmem_n7895), .ZN(MEM_stage_inst_dmem_n5001) );
NAND2_X1 MEM_stage_inst_dmem_U5130 ( .A1(MEM_stage_inst_dmem_ram_1129), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n5002) );
NAND2_X1 MEM_stage_inst_dmem_U5129 ( .A1(MEM_stage_inst_dmem_n5000), .A2(MEM_stage_inst_dmem_n4999), .ZN(MEM_stage_inst_dmem_n5004) );
NAND2_X1 MEM_stage_inst_dmem_U5128 ( .A1(MEM_stage_inst_dmem_ram_1705), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n4999) );
NAND2_X1 MEM_stage_inst_dmem_U5127 ( .A1(MEM_stage_inst_dmem_ram_1753), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n5000) );
NAND2_X1 MEM_stage_inst_dmem_U5126 ( .A1(MEM_stage_inst_dmem_n4998), .A2(MEM_stage_inst_dmem_n4997), .ZN(MEM_stage_inst_dmem_n5014) );
NOR2_X1 MEM_stage_inst_dmem_U5125 ( .A1(MEM_stage_inst_dmem_n4996), .A2(MEM_stage_inst_dmem_n4995), .ZN(MEM_stage_inst_dmem_n4997) );
NAND2_X1 MEM_stage_inst_dmem_U5124 ( .A1(MEM_stage_inst_dmem_n4994), .A2(MEM_stage_inst_dmem_n4993), .ZN(MEM_stage_inst_dmem_n4995) );
NAND2_X1 MEM_stage_inst_dmem_U5123 ( .A1(MEM_stage_inst_dmem_ram_1993), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n4993) );
NAND2_X1 MEM_stage_inst_dmem_U5122 ( .A1(MEM_stage_inst_dmem_ram_1625), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n4994) );
NAND2_X1 MEM_stage_inst_dmem_U5121 ( .A1(MEM_stage_inst_dmem_n4992), .A2(MEM_stage_inst_dmem_n4991), .ZN(MEM_stage_inst_dmem_n4996) );
NAND2_X1 MEM_stage_inst_dmem_U5120 ( .A1(MEM_stage_inst_dmem_ram_1513), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n4991) );
NAND2_X1 MEM_stage_inst_dmem_U5119 ( .A1(MEM_stage_inst_dmem_ram_1177), .A2(MEM_stage_inst_dmem_n7903), .ZN(MEM_stage_inst_dmem_n4992) );
NOR2_X1 MEM_stage_inst_dmem_U5118 ( .A1(MEM_stage_inst_dmem_n4990), .A2(MEM_stage_inst_dmem_n4989), .ZN(MEM_stage_inst_dmem_n4998) );
NAND2_X1 MEM_stage_inst_dmem_U5117 ( .A1(MEM_stage_inst_dmem_n4988), .A2(MEM_stage_inst_dmem_n4987), .ZN(MEM_stage_inst_dmem_n4989) );
NAND2_X1 MEM_stage_inst_dmem_U5116 ( .A1(MEM_stage_inst_dmem_ram_1881), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n4987) );
NAND2_X1 MEM_stage_inst_dmem_U5115 ( .A1(MEM_stage_inst_dmem_ram_1593), .A2(MEM_stage_inst_dmem_n41), .ZN(MEM_stage_inst_dmem_n4988) );
NAND2_X1 MEM_stage_inst_dmem_U5114 ( .A1(MEM_stage_inst_dmem_n4986), .A2(MEM_stage_inst_dmem_n4985), .ZN(MEM_stage_inst_dmem_n4990) );
NAND2_X1 MEM_stage_inst_dmem_U5113 ( .A1(MEM_stage_inst_dmem_ram_1865), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n4985) );
NAND2_X1 MEM_stage_inst_dmem_U5112 ( .A1(MEM_stage_inst_dmem_ram_1145), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n4986) );
NAND2_X1 MEM_stage_inst_dmem_U5111 ( .A1(MEM_stage_inst_dmem_n4984), .A2(MEM_stage_inst_dmem_n4983), .ZN(MEM_stage_inst_dmem_n5048) );
NOR2_X1 MEM_stage_inst_dmem_U5110 ( .A1(MEM_stage_inst_dmem_n4982), .A2(MEM_stage_inst_dmem_n4981), .ZN(MEM_stage_inst_dmem_n4983) );
NAND2_X1 MEM_stage_inst_dmem_U5109 ( .A1(MEM_stage_inst_dmem_n4980), .A2(MEM_stage_inst_dmem_n4979), .ZN(MEM_stage_inst_dmem_n4981) );
NOR2_X1 MEM_stage_inst_dmem_U5108 ( .A1(MEM_stage_inst_dmem_n4978), .A2(MEM_stage_inst_dmem_n4977), .ZN(MEM_stage_inst_dmem_n4979) );
NAND2_X1 MEM_stage_inst_dmem_U5107 ( .A1(MEM_stage_inst_dmem_n4976), .A2(MEM_stage_inst_dmem_n4975), .ZN(MEM_stage_inst_dmem_n4977) );
NAND2_X1 MEM_stage_inst_dmem_U5106 ( .A1(MEM_stage_inst_dmem_ram_1897), .A2(MEM_stage_inst_dmem_n7923), .ZN(MEM_stage_inst_dmem_n4975) );
NAND2_X1 MEM_stage_inst_dmem_U5105 ( .A1(MEM_stage_inst_dmem_ram_1065), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n4976) );
NAND2_X1 MEM_stage_inst_dmem_U5104 ( .A1(MEM_stage_inst_dmem_n4974), .A2(MEM_stage_inst_dmem_n4973), .ZN(MEM_stage_inst_dmem_n4978) );
NAND2_X1 MEM_stage_inst_dmem_U5103 ( .A1(MEM_stage_inst_dmem_ram_1529), .A2(MEM_stage_inst_dmem_n64), .ZN(MEM_stage_inst_dmem_n4973) );
NAND2_X1 MEM_stage_inst_dmem_U5102 ( .A1(MEM_stage_inst_dmem_ram_1961), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n4974) );
NOR2_X1 MEM_stage_inst_dmem_U5101 ( .A1(MEM_stage_inst_dmem_n4972), .A2(MEM_stage_inst_dmem_n4971), .ZN(MEM_stage_inst_dmem_n4980) );
NAND2_X1 MEM_stage_inst_dmem_U5100 ( .A1(MEM_stage_inst_dmem_n4970), .A2(MEM_stage_inst_dmem_n4969), .ZN(MEM_stage_inst_dmem_n4971) );
NAND2_X1 MEM_stage_inst_dmem_U5099 ( .A1(MEM_stage_inst_dmem_ram_1721), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n4969) );
NAND2_X1 MEM_stage_inst_dmem_U5098 ( .A1(MEM_stage_inst_dmem_ram_1689), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n4970) );
NAND2_X1 MEM_stage_inst_dmem_U5097 ( .A1(MEM_stage_inst_dmem_n4968), .A2(MEM_stage_inst_dmem_n4967), .ZN(MEM_stage_inst_dmem_n4972) );
NAND2_X1 MEM_stage_inst_dmem_U5096 ( .A1(MEM_stage_inst_dmem_ram_1945), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n4967) );
NAND2_X1 MEM_stage_inst_dmem_U5095 ( .A1(MEM_stage_inst_dmem_ram_1481), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n4968) );
NAND2_X1 MEM_stage_inst_dmem_U5094 ( .A1(MEM_stage_inst_dmem_n4966), .A2(MEM_stage_inst_dmem_n4965), .ZN(MEM_stage_inst_dmem_n4982) );
NOR2_X1 MEM_stage_inst_dmem_U5093 ( .A1(MEM_stage_inst_dmem_n4964), .A2(MEM_stage_inst_dmem_n4963), .ZN(MEM_stage_inst_dmem_n4965) );
NAND2_X1 MEM_stage_inst_dmem_U5092 ( .A1(MEM_stage_inst_dmem_n4962), .A2(MEM_stage_inst_dmem_n4961), .ZN(MEM_stage_inst_dmem_n4963) );
NAND2_X1 MEM_stage_inst_dmem_U5091 ( .A1(MEM_stage_inst_dmem_ram_1449), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n4961) );
NAND2_X1 MEM_stage_inst_dmem_U5090 ( .A1(MEM_stage_inst_dmem_ram_1033), .A2(MEM_stage_inst_dmem_n7953), .ZN(MEM_stage_inst_dmem_n4962) );
NAND2_X1 MEM_stage_inst_dmem_U5089 ( .A1(MEM_stage_inst_dmem_n4960), .A2(MEM_stage_inst_dmem_n4959), .ZN(MEM_stage_inst_dmem_n4964) );
NAND2_X1 MEM_stage_inst_dmem_U5088 ( .A1(MEM_stage_inst_dmem_ram_1737), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n4959) );
NAND2_X1 MEM_stage_inst_dmem_U5087 ( .A1(MEM_stage_inst_dmem_ram_1369), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n4960) );
NOR2_X1 MEM_stage_inst_dmem_U5086 ( .A1(MEM_stage_inst_dmem_n4958), .A2(MEM_stage_inst_dmem_n4957), .ZN(MEM_stage_inst_dmem_n4966) );
NAND2_X1 MEM_stage_inst_dmem_U5085 ( .A1(MEM_stage_inst_dmem_n4956), .A2(MEM_stage_inst_dmem_n4955), .ZN(MEM_stage_inst_dmem_n4957) );
NAND2_X1 MEM_stage_inst_dmem_U5084 ( .A1(MEM_stage_inst_dmem_ram_1225), .A2(MEM_stage_inst_dmem_n36), .ZN(MEM_stage_inst_dmem_n4955) );
NAND2_X1 MEM_stage_inst_dmem_U5083 ( .A1(MEM_stage_inst_dmem_ram_1289), .A2(MEM_stage_inst_dmem_n7898), .ZN(MEM_stage_inst_dmem_n4956) );
NAND2_X1 MEM_stage_inst_dmem_U5082 ( .A1(MEM_stage_inst_dmem_n4954), .A2(MEM_stage_inst_dmem_n4953), .ZN(MEM_stage_inst_dmem_n4958) );
NAND2_X1 MEM_stage_inst_dmem_U5081 ( .A1(MEM_stage_inst_dmem_ram_1785), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n4953) );
NAND2_X1 MEM_stage_inst_dmem_U5080 ( .A1(MEM_stage_inst_dmem_ram_1577), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n4954) );
NOR2_X1 MEM_stage_inst_dmem_U5079 ( .A1(MEM_stage_inst_dmem_n4952), .A2(MEM_stage_inst_dmem_n4951), .ZN(MEM_stage_inst_dmem_n4984) );
NAND2_X1 MEM_stage_inst_dmem_U5078 ( .A1(MEM_stage_inst_dmem_n4950), .A2(MEM_stage_inst_dmem_n4949), .ZN(MEM_stage_inst_dmem_n4951) );
NOR2_X1 MEM_stage_inst_dmem_U5077 ( .A1(MEM_stage_inst_dmem_n4948), .A2(MEM_stage_inst_dmem_n4947), .ZN(MEM_stage_inst_dmem_n4949) );
NAND2_X1 MEM_stage_inst_dmem_U5076 ( .A1(MEM_stage_inst_dmem_n4946), .A2(MEM_stage_inst_dmem_n4945), .ZN(MEM_stage_inst_dmem_n4947) );
NAND2_X1 MEM_stage_inst_dmem_U5075 ( .A1(MEM_stage_inst_dmem_ram_1097), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n4945) );
NAND2_X1 MEM_stage_inst_dmem_U5074 ( .A1(MEM_stage_inst_dmem_ram_1609), .A2(MEM_stage_inst_dmem_n7973), .ZN(MEM_stage_inst_dmem_n4946) );
NAND2_X1 MEM_stage_inst_dmem_U5073 ( .A1(MEM_stage_inst_dmem_n4944), .A2(MEM_stage_inst_dmem_n4943), .ZN(MEM_stage_inst_dmem_n4948) );
NAND2_X1 MEM_stage_inst_dmem_U5072 ( .A1(MEM_stage_inst_dmem_ram_1081), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n4943) );
NAND2_X1 MEM_stage_inst_dmem_U5071 ( .A1(MEM_stage_inst_dmem_ram_1417), .A2(MEM_stage_inst_dmem_n7930), .ZN(MEM_stage_inst_dmem_n4944) );
NOR2_X1 MEM_stage_inst_dmem_U5070 ( .A1(MEM_stage_inst_dmem_n4942), .A2(MEM_stage_inst_dmem_n4941), .ZN(MEM_stage_inst_dmem_n4950) );
NAND2_X1 MEM_stage_inst_dmem_U5069 ( .A1(MEM_stage_inst_dmem_n4940), .A2(MEM_stage_inst_dmem_n4939), .ZN(MEM_stage_inst_dmem_n4941) );
NAND2_X1 MEM_stage_inst_dmem_U5068 ( .A1(MEM_stage_inst_dmem_ram_1161), .A2(MEM_stage_inst_dmem_n61), .ZN(MEM_stage_inst_dmem_n4939) );
NAND2_X1 MEM_stage_inst_dmem_U5067 ( .A1(MEM_stage_inst_dmem_ram_1817), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n4940) );
NAND2_X1 MEM_stage_inst_dmem_U5066 ( .A1(MEM_stage_inst_dmem_n4938), .A2(MEM_stage_inst_dmem_n4937), .ZN(MEM_stage_inst_dmem_n4942) );
NAND2_X1 MEM_stage_inst_dmem_U5065 ( .A1(MEM_stage_inst_dmem_ram_1353), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n4937) );
NAND2_X1 MEM_stage_inst_dmem_U5064 ( .A1(MEM_stage_inst_dmem_ram_1305), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n4938) );
NAND2_X1 MEM_stage_inst_dmem_U5063 ( .A1(MEM_stage_inst_dmem_n4936), .A2(MEM_stage_inst_dmem_n4935), .ZN(MEM_stage_inst_dmem_n4952) );
NOR2_X1 MEM_stage_inst_dmem_U5062 ( .A1(MEM_stage_inst_dmem_n4934), .A2(MEM_stage_inst_dmem_n4933), .ZN(MEM_stage_inst_dmem_n4935) );
NAND2_X1 MEM_stage_inst_dmem_U5061 ( .A1(MEM_stage_inst_dmem_n4932), .A2(MEM_stage_inst_dmem_n4931), .ZN(MEM_stage_inst_dmem_n4933) );
NAND2_X1 MEM_stage_inst_dmem_U5060 ( .A1(MEM_stage_inst_dmem_ram_1337), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n4931) );
NAND2_X1 MEM_stage_inst_dmem_U5059 ( .A1(MEM_stage_inst_dmem_ram_1497), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n4932) );
NAND2_X1 MEM_stage_inst_dmem_U5058 ( .A1(MEM_stage_inst_dmem_n4930), .A2(MEM_stage_inst_dmem_n4929), .ZN(MEM_stage_inst_dmem_n4934) );
NAND2_X1 MEM_stage_inst_dmem_U5057 ( .A1(MEM_stage_inst_dmem_ram_1561), .A2(MEM_stage_inst_dmem_n7884), .ZN(MEM_stage_inst_dmem_n4929) );
NAND2_X1 MEM_stage_inst_dmem_U5056 ( .A1(MEM_stage_inst_dmem_ram_1769), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n4930) );
NOR2_X1 MEM_stage_inst_dmem_U5055 ( .A1(MEM_stage_inst_dmem_n4928), .A2(MEM_stage_inst_dmem_n4927), .ZN(MEM_stage_inst_dmem_n4936) );
NAND2_X1 MEM_stage_inst_dmem_U5054 ( .A1(MEM_stage_inst_dmem_n4926), .A2(MEM_stage_inst_dmem_n4925), .ZN(MEM_stage_inst_dmem_n4927) );
NAND2_X1 MEM_stage_inst_dmem_U5053 ( .A1(MEM_stage_inst_dmem_ram_2025), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n4925) );
NAND2_X1 MEM_stage_inst_dmem_U5052 ( .A1(MEM_stage_inst_dmem_ram_1193), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n4926) );
NAND2_X1 MEM_stage_inst_dmem_U5051 ( .A1(MEM_stage_inst_dmem_n4924), .A2(MEM_stage_inst_dmem_n4923), .ZN(MEM_stage_inst_dmem_n4928) );
NAND2_X1 MEM_stage_inst_dmem_U5050 ( .A1(MEM_stage_inst_dmem_ram_1385), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n4923) );
NAND2_X1 MEM_stage_inst_dmem_U5049 ( .A1(MEM_stage_inst_dmem_ram_1113), .A2(MEM_stage_inst_dmem_n7938), .ZN(MEM_stage_inst_dmem_n4924) );
NAND2_X1 MEM_stage_inst_dmem_U5048 ( .A1(MEM_stage_inst_dmem_n4922), .A2(MEM_stage_inst_dmem_n4921), .ZN(MEM_stage_inst_mem_read_data_8) );
NOR2_X1 MEM_stage_inst_dmem_U5047 ( .A1(MEM_stage_inst_dmem_n4920), .A2(MEM_stage_inst_dmem_n4919), .ZN(MEM_stage_inst_dmem_n4921) );
NOR2_X1 MEM_stage_inst_dmem_U5046 ( .A1(MEM_stage_inst_dmem_n4918), .A2(MEM_stage_inst_dmem_n8551), .ZN(MEM_stage_inst_dmem_n4919) );
NOR2_X1 MEM_stage_inst_dmem_U5045 ( .A1(MEM_stage_inst_dmem_n4917), .A2(MEM_stage_inst_dmem_n4916), .ZN(MEM_stage_inst_dmem_n4918) );
NAND2_X1 MEM_stage_inst_dmem_U5044 ( .A1(MEM_stage_inst_dmem_n4915), .A2(MEM_stage_inst_dmem_n4914), .ZN(MEM_stage_inst_dmem_n4916) );
NOR2_X1 MEM_stage_inst_dmem_U5043 ( .A1(MEM_stage_inst_dmem_n4913), .A2(MEM_stage_inst_dmem_n4912), .ZN(MEM_stage_inst_dmem_n4914) );
NAND2_X1 MEM_stage_inst_dmem_U5042 ( .A1(MEM_stage_inst_dmem_n4911), .A2(MEM_stage_inst_dmem_n4910), .ZN(MEM_stage_inst_dmem_n4912) );
NOR2_X1 MEM_stage_inst_dmem_U5041 ( .A1(MEM_stage_inst_dmem_n4909), .A2(MEM_stage_inst_dmem_n4908), .ZN(MEM_stage_inst_dmem_n4910) );
NAND2_X1 MEM_stage_inst_dmem_U5040 ( .A1(MEM_stage_inst_dmem_n4907), .A2(MEM_stage_inst_dmem_n4906), .ZN(MEM_stage_inst_dmem_n4908) );
NAND2_X1 MEM_stage_inst_dmem_U5039 ( .A1(MEM_stage_inst_dmem_ram_840), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n4906) );
NAND2_X1 MEM_stage_inst_dmem_U5038 ( .A1(MEM_stage_inst_dmem_ram_744), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n4907) );
NAND2_X1 MEM_stage_inst_dmem_U5037 ( .A1(MEM_stage_inst_dmem_n4905), .A2(MEM_stage_inst_dmem_n4904), .ZN(MEM_stage_inst_dmem_n4909) );
NAND2_X1 MEM_stage_inst_dmem_U5036 ( .A1(MEM_stage_inst_dmem_ram_24), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n4904) );
NAND2_X1 MEM_stage_inst_dmem_U5035 ( .A1(MEM_stage_inst_dmem_ram_1016), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n4905) );
NOR2_X1 MEM_stage_inst_dmem_U5034 ( .A1(MEM_stage_inst_dmem_n4903), .A2(MEM_stage_inst_dmem_n4902), .ZN(MEM_stage_inst_dmem_n4911) );
NAND2_X1 MEM_stage_inst_dmem_U5033 ( .A1(MEM_stage_inst_dmem_n4901), .A2(MEM_stage_inst_dmem_n4900), .ZN(MEM_stage_inst_dmem_n4902) );
NAND2_X1 MEM_stage_inst_dmem_U5032 ( .A1(MEM_stage_inst_dmem_ram_856), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n4900) );
NAND2_X1 MEM_stage_inst_dmem_U5031 ( .A1(MEM_stage_inst_dmem_ram_344), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n4901) );
NAND2_X1 MEM_stage_inst_dmem_U5030 ( .A1(MEM_stage_inst_dmem_n4899), .A2(MEM_stage_inst_dmem_n4898), .ZN(MEM_stage_inst_dmem_n4903) );
NAND2_X1 MEM_stage_inst_dmem_U5029 ( .A1(MEM_stage_inst_dmem_ram_776), .A2(MEM_stage_inst_dmem_n37), .ZN(MEM_stage_inst_dmem_n4898) );
NAND2_X1 MEM_stage_inst_dmem_U5028 ( .A1(MEM_stage_inst_dmem_ram_440), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n4899) );
NAND2_X1 MEM_stage_inst_dmem_U5027 ( .A1(MEM_stage_inst_dmem_n4897), .A2(MEM_stage_inst_dmem_n4896), .ZN(MEM_stage_inst_dmem_n4913) );
NOR2_X1 MEM_stage_inst_dmem_U5026 ( .A1(MEM_stage_inst_dmem_n4895), .A2(MEM_stage_inst_dmem_n4894), .ZN(MEM_stage_inst_dmem_n4896) );
NAND2_X1 MEM_stage_inst_dmem_U5025 ( .A1(MEM_stage_inst_dmem_n4893), .A2(MEM_stage_inst_dmem_n4892), .ZN(MEM_stage_inst_dmem_n4894) );
NAND2_X1 MEM_stage_inst_dmem_U5024 ( .A1(MEM_stage_inst_dmem_ram_904), .A2(MEM_stage_inst_dmem_n72), .ZN(MEM_stage_inst_dmem_n4892) );
NAND2_X1 MEM_stage_inst_dmem_U5023 ( .A1(MEM_stage_inst_dmem_ram_808), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n4893) );
NAND2_X1 MEM_stage_inst_dmem_U5022 ( .A1(MEM_stage_inst_dmem_n4891), .A2(MEM_stage_inst_dmem_n4890), .ZN(MEM_stage_inst_dmem_n4895) );
NAND2_X1 MEM_stage_inst_dmem_U5021 ( .A1(MEM_stage_inst_dmem_ram_392), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n4890) );
NAND2_X1 MEM_stage_inst_dmem_U5020 ( .A1(MEM_stage_inst_dmem_ram_376), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n4891) );
NOR2_X1 MEM_stage_inst_dmem_U5019 ( .A1(MEM_stage_inst_dmem_n4889), .A2(MEM_stage_inst_dmem_n4888), .ZN(MEM_stage_inst_dmem_n4897) );
NAND2_X1 MEM_stage_inst_dmem_U5018 ( .A1(MEM_stage_inst_dmem_n4887), .A2(MEM_stage_inst_dmem_n4886), .ZN(MEM_stage_inst_dmem_n4888) );
NAND2_X1 MEM_stage_inst_dmem_U5017 ( .A1(MEM_stage_inst_dmem_ram_200), .A2(MEM_stage_inst_dmem_n36), .ZN(MEM_stage_inst_dmem_n4886) );
NAND2_X1 MEM_stage_inst_dmem_U5016 ( .A1(MEM_stage_inst_dmem_ram_552), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n4887) );
NAND2_X1 MEM_stage_inst_dmem_U5015 ( .A1(MEM_stage_inst_dmem_n4885), .A2(MEM_stage_inst_dmem_n4884), .ZN(MEM_stage_inst_dmem_n4889) );
NAND2_X1 MEM_stage_inst_dmem_U5014 ( .A1(MEM_stage_inst_dmem_ram_408), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n4884) );
NAND2_X1 MEM_stage_inst_dmem_U5013 ( .A1(MEM_stage_inst_dmem_ram_600), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n4885) );
NOR2_X1 MEM_stage_inst_dmem_U5012 ( .A1(MEM_stage_inst_dmem_n4883), .A2(MEM_stage_inst_dmem_n4882), .ZN(MEM_stage_inst_dmem_n4915) );
NAND2_X1 MEM_stage_inst_dmem_U5011 ( .A1(MEM_stage_inst_dmem_n4881), .A2(MEM_stage_inst_dmem_n4880), .ZN(MEM_stage_inst_dmem_n4882) );
NOR2_X1 MEM_stage_inst_dmem_U5010 ( .A1(MEM_stage_inst_dmem_n4879), .A2(MEM_stage_inst_dmem_n4878), .ZN(MEM_stage_inst_dmem_n4880) );
NAND2_X1 MEM_stage_inst_dmem_U5009 ( .A1(MEM_stage_inst_dmem_n4877), .A2(MEM_stage_inst_dmem_n4876), .ZN(MEM_stage_inst_dmem_n4878) );
NAND2_X1 MEM_stage_inst_dmem_U5008 ( .A1(MEM_stage_inst_dmem_ram_920), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n4876) );
NAND2_X1 MEM_stage_inst_dmem_U5007 ( .A1(MEM_stage_inst_dmem_ram_536), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n4877) );
NAND2_X1 MEM_stage_inst_dmem_U5006 ( .A1(MEM_stage_inst_dmem_n4875), .A2(MEM_stage_inst_dmem_n4874), .ZN(MEM_stage_inst_dmem_n4879) );
NAND2_X1 MEM_stage_inst_dmem_U5005 ( .A1(MEM_stage_inst_dmem_ram_488), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n4874) );
NAND2_X1 MEM_stage_inst_dmem_U5004 ( .A1(MEM_stage_inst_dmem_ram_168), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n4875) );
NOR2_X1 MEM_stage_inst_dmem_U5003 ( .A1(MEM_stage_inst_dmem_n4873), .A2(MEM_stage_inst_dmem_n4872), .ZN(MEM_stage_inst_dmem_n4881) );
NAND2_X1 MEM_stage_inst_dmem_U5002 ( .A1(MEM_stage_inst_dmem_n4871), .A2(MEM_stage_inst_dmem_n4870), .ZN(MEM_stage_inst_dmem_n4872) );
NAND2_X1 MEM_stage_inst_dmem_U5001 ( .A1(MEM_stage_inst_dmem_ram_232), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n4870) );
NAND2_X1 MEM_stage_inst_dmem_U5000 ( .A1(MEM_stage_inst_dmem_ram_88), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n4871) );
NAND2_X1 MEM_stage_inst_dmem_U4999 ( .A1(MEM_stage_inst_dmem_n4869), .A2(MEM_stage_inst_dmem_n4868), .ZN(MEM_stage_inst_dmem_n4873) );
NAND2_X1 MEM_stage_inst_dmem_U4998 ( .A1(MEM_stage_inst_dmem_ram_360), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n4868) );
NAND2_X1 MEM_stage_inst_dmem_U4997 ( .A1(MEM_stage_inst_dmem_ram_936), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n4869) );
NAND2_X1 MEM_stage_inst_dmem_U4996 ( .A1(MEM_stage_inst_dmem_n4867), .A2(MEM_stage_inst_dmem_n4866), .ZN(MEM_stage_inst_dmem_n4883) );
NOR2_X1 MEM_stage_inst_dmem_U4995 ( .A1(MEM_stage_inst_dmem_n4865), .A2(MEM_stage_inst_dmem_n4864), .ZN(MEM_stage_inst_dmem_n4866) );
NAND2_X1 MEM_stage_inst_dmem_U4994 ( .A1(MEM_stage_inst_dmem_n4863), .A2(MEM_stage_inst_dmem_n4862), .ZN(MEM_stage_inst_dmem_n4864) );
NAND2_X1 MEM_stage_inst_dmem_U4993 ( .A1(MEM_stage_inst_dmem_ram_888), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n4862) );
NAND2_X1 MEM_stage_inst_dmem_U4992 ( .A1(MEM_stage_inst_dmem_ram_616), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n4863) );
NAND2_X1 MEM_stage_inst_dmem_U4991 ( .A1(MEM_stage_inst_dmem_n4861), .A2(MEM_stage_inst_dmem_n4860), .ZN(MEM_stage_inst_dmem_n4865) );
NAND2_X1 MEM_stage_inst_dmem_U4990 ( .A1(MEM_stage_inst_dmem_ram_968), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n4860) );
NAND2_X1 MEM_stage_inst_dmem_U4989 ( .A1(MEM_stage_inst_dmem_ram_296), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n4861) );
NOR2_X1 MEM_stage_inst_dmem_U4988 ( .A1(MEM_stage_inst_dmem_n4859), .A2(MEM_stage_inst_dmem_n4858), .ZN(MEM_stage_inst_dmem_n4867) );
NAND2_X1 MEM_stage_inst_dmem_U4987 ( .A1(MEM_stage_inst_dmem_n4857), .A2(MEM_stage_inst_dmem_n4856), .ZN(MEM_stage_inst_dmem_n4858) );
NAND2_X1 MEM_stage_inst_dmem_U4986 ( .A1(MEM_stage_inst_dmem_ram_824), .A2(MEM_stage_inst_dmem_n46), .ZN(MEM_stage_inst_dmem_n4856) );
NAND2_X1 MEM_stage_inst_dmem_U4985 ( .A1(MEM_stage_inst_dmem_ram_456), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n4857) );
NAND2_X1 MEM_stage_inst_dmem_U4984 ( .A1(MEM_stage_inst_dmem_n4855), .A2(MEM_stage_inst_dmem_n4854), .ZN(MEM_stage_inst_dmem_n4859) );
NAND2_X1 MEM_stage_inst_dmem_U4983 ( .A1(MEM_stage_inst_dmem_ram_1000), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n4854) );
NAND2_X1 MEM_stage_inst_dmem_U4982 ( .A1(MEM_stage_inst_dmem_ram_120), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n4855) );
NAND2_X1 MEM_stage_inst_dmem_U4981 ( .A1(MEM_stage_inst_dmem_n4853), .A2(MEM_stage_inst_dmem_n4852), .ZN(MEM_stage_inst_dmem_n4917) );
NOR2_X1 MEM_stage_inst_dmem_U4980 ( .A1(MEM_stage_inst_dmem_n4851), .A2(MEM_stage_inst_dmem_n4850), .ZN(MEM_stage_inst_dmem_n4852) );
NAND2_X1 MEM_stage_inst_dmem_U4979 ( .A1(MEM_stage_inst_dmem_n4849), .A2(MEM_stage_inst_dmem_n4848), .ZN(MEM_stage_inst_dmem_n4850) );
NOR2_X1 MEM_stage_inst_dmem_U4978 ( .A1(MEM_stage_inst_dmem_n4847), .A2(MEM_stage_inst_dmem_n4846), .ZN(MEM_stage_inst_dmem_n4848) );
NAND2_X1 MEM_stage_inst_dmem_U4977 ( .A1(MEM_stage_inst_dmem_n4845), .A2(MEM_stage_inst_dmem_n4844), .ZN(MEM_stage_inst_dmem_n4846) );
NAND2_X1 MEM_stage_inst_dmem_U4976 ( .A1(MEM_stage_inst_dmem_ram_216), .A2(MEM_stage_inst_dmem_n51), .ZN(MEM_stage_inst_dmem_n4844) );
NAND2_X1 MEM_stage_inst_dmem_U4975 ( .A1(MEM_stage_inst_dmem_ram_584), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n4845) );
NAND2_X1 MEM_stage_inst_dmem_U4974 ( .A1(MEM_stage_inst_dmem_n4843), .A2(MEM_stage_inst_dmem_n4842), .ZN(MEM_stage_inst_dmem_n4847) );
NAND2_X1 MEM_stage_inst_dmem_U4973 ( .A1(MEM_stage_inst_dmem_ram_760), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n4842) );
NAND2_X1 MEM_stage_inst_dmem_U4972 ( .A1(MEM_stage_inst_dmem_ram_664), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n4843) );
NOR2_X1 MEM_stage_inst_dmem_U4971 ( .A1(MEM_stage_inst_dmem_n4841), .A2(MEM_stage_inst_dmem_n4840), .ZN(MEM_stage_inst_dmem_n4849) );
NAND2_X1 MEM_stage_inst_dmem_U4970 ( .A1(MEM_stage_inst_dmem_n4839), .A2(MEM_stage_inst_dmem_n4838), .ZN(MEM_stage_inst_dmem_n4840) );
NAND2_X1 MEM_stage_inst_dmem_U4969 ( .A1(MEM_stage_inst_dmem_ram_184), .A2(MEM_stage_inst_dmem_n55), .ZN(MEM_stage_inst_dmem_n4838) );
NAND2_X1 MEM_stage_inst_dmem_U4968 ( .A1(MEM_stage_inst_dmem_ram_104), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n4839) );
NAND2_X1 MEM_stage_inst_dmem_U4967 ( .A1(MEM_stage_inst_dmem_n4837), .A2(MEM_stage_inst_dmem_n4836), .ZN(MEM_stage_inst_dmem_n4841) );
NAND2_X1 MEM_stage_inst_dmem_U4966 ( .A1(MEM_stage_inst_dmem_ram_872), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n4836) );
NAND2_X1 MEM_stage_inst_dmem_U4965 ( .A1(MEM_stage_inst_dmem_ram_568), .A2(MEM_stage_inst_dmem_n41), .ZN(MEM_stage_inst_dmem_n4837) );
NAND2_X1 MEM_stage_inst_dmem_U4964 ( .A1(MEM_stage_inst_dmem_n4835), .A2(MEM_stage_inst_dmem_n4834), .ZN(MEM_stage_inst_dmem_n4851) );
NOR2_X1 MEM_stage_inst_dmem_U4963 ( .A1(MEM_stage_inst_dmem_n4833), .A2(MEM_stage_inst_dmem_n4832), .ZN(MEM_stage_inst_dmem_n4834) );
NAND2_X1 MEM_stage_inst_dmem_U4962 ( .A1(MEM_stage_inst_dmem_n4831), .A2(MEM_stage_inst_dmem_n4830), .ZN(MEM_stage_inst_dmem_n4832) );
NAND2_X1 MEM_stage_inst_dmem_U4961 ( .A1(MEM_stage_inst_dmem_ram_696), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n4830) );
NAND2_X1 MEM_stage_inst_dmem_U4960 ( .A1(MEM_stage_inst_dmem_ram_520), .A2(MEM_stage_inst_dmem_n71), .ZN(MEM_stage_inst_dmem_n4831) );
NAND2_X1 MEM_stage_inst_dmem_U4959 ( .A1(MEM_stage_inst_dmem_n4829), .A2(MEM_stage_inst_dmem_n4828), .ZN(MEM_stage_inst_dmem_n4833) );
NAND2_X1 MEM_stage_inst_dmem_U4958 ( .A1(MEM_stage_inst_dmem_ram_56), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n4828) );
NAND2_X1 MEM_stage_inst_dmem_U4957 ( .A1(MEM_stage_inst_dmem_ram_680), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n4829) );
NOR2_X1 MEM_stage_inst_dmem_U4956 ( .A1(MEM_stage_inst_dmem_n4827), .A2(MEM_stage_inst_dmem_n4826), .ZN(MEM_stage_inst_dmem_n4835) );
NAND2_X1 MEM_stage_inst_dmem_U4955 ( .A1(MEM_stage_inst_dmem_n4825), .A2(MEM_stage_inst_dmem_n4824), .ZN(MEM_stage_inst_dmem_n4826) );
NAND2_X1 MEM_stage_inst_dmem_U4954 ( .A1(MEM_stage_inst_dmem_ram_504), .A2(MEM_stage_inst_dmem_n64), .ZN(MEM_stage_inst_dmem_n4824) );
NAND2_X1 MEM_stage_inst_dmem_U4953 ( .A1(MEM_stage_inst_dmem_ram_952), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n4825) );
NAND2_X1 MEM_stage_inst_dmem_U4952 ( .A1(MEM_stage_inst_dmem_n4823), .A2(MEM_stage_inst_dmem_n4822), .ZN(MEM_stage_inst_dmem_n4827) );
NAND2_X1 MEM_stage_inst_dmem_U4951 ( .A1(MEM_stage_inst_dmem_ram_472), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n4822) );
NAND2_X1 MEM_stage_inst_dmem_U4950 ( .A1(MEM_stage_inst_dmem_ram_632), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n4823) );
NOR2_X1 MEM_stage_inst_dmem_U4949 ( .A1(MEM_stage_inst_dmem_n4821), .A2(MEM_stage_inst_dmem_n4820), .ZN(MEM_stage_inst_dmem_n4853) );
NAND2_X1 MEM_stage_inst_dmem_U4948 ( .A1(MEM_stage_inst_dmem_n4819), .A2(MEM_stage_inst_dmem_n4818), .ZN(MEM_stage_inst_dmem_n4820) );
NOR2_X1 MEM_stage_inst_dmem_U4947 ( .A1(MEM_stage_inst_dmem_n4817), .A2(MEM_stage_inst_dmem_n4816), .ZN(MEM_stage_inst_dmem_n4818) );
NAND2_X1 MEM_stage_inst_dmem_U4946 ( .A1(MEM_stage_inst_dmem_n4815), .A2(MEM_stage_inst_dmem_n4814), .ZN(MEM_stage_inst_dmem_n4816) );
NAND2_X1 MEM_stage_inst_dmem_U4945 ( .A1(MEM_stage_inst_dmem_ram_312), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n4814) );
NAND2_X1 MEM_stage_inst_dmem_U4944 ( .A1(MEM_stage_inst_dmem_ram_984), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n4815) );
NAND2_X1 MEM_stage_inst_dmem_U4943 ( .A1(MEM_stage_inst_dmem_n4813), .A2(MEM_stage_inst_dmem_n4812), .ZN(MEM_stage_inst_dmem_n4817) );
NAND2_X1 MEM_stage_inst_dmem_U4942 ( .A1(MEM_stage_inst_dmem_ram_792), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n4812) );
NAND2_X1 MEM_stage_inst_dmem_U4941 ( .A1(MEM_stage_inst_dmem_ram_728), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n4813) );
NOR2_X1 MEM_stage_inst_dmem_U4940 ( .A1(MEM_stage_inst_dmem_n4811), .A2(MEM_stage_inst_dmem_n4810), .ZN(MEM_stage_inst_dmem_n4819) );
NAND2_X1 MEM_stage_inst_dmem_U4939 ( .A1(MEM_stage_inst_dmem_n4809), .A2(MEM_stage_inst_dmem_n4808), .ZN(MEM_stage_inst_dmem_n4810) );
NAND2_X1 MEM_stage_inst_dmem_U4938 ( .A1(MEM_stage_inst_dmem_ram_136), .A2(MEM_stage_inst_dmem_n61), .ZN(MEM_stage_inst_dmem_n4808) );
NAND2_X1 MEM_stage_inst_dmem_U4937 ( .A1(MEM_stage_inst_dmem_ram_40), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n4809) );
NAND2_X1 MEM_stage_inst_dmem_U4936 ( .A1(MEM_stage_inst_dmem_n4807), .A2(MEM_stage_inst_dmem_n4806), .ZN(MEM_stage_inst_dmem_n4811) );
NAND2_X1 MEM_stage_inst_dmem_U4935 ( .A1(MEM_stage_inst_dmem_ram_328), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n4806) );
NAND2_X1 MEM_stage_inst_dmem_U4934 ( .A1(MEM_stage_inst_dmem_ram_648), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n4807) );
NAND2_X1 MEM_stage_inst_dmem_U4933 ( .A1(MEM_stage_inst_dmem_n4805), .A2(MEM_stage_inst_dmem_n4804), .ZN(MEM_stage_inst_dmem_n4821) );
NOR2_X1 MEM_stage_inst_dmem_U4932 ( .A1(MEM_stage_inst_dmem_n4803), .A2(MEM_stage_inst_dmem_n4802), .ZN(MEM_stage_inst_dmem_n4804) );
NAND2_X1 MEM_stage_inst_dmem_U4931 ( .A1(MEM_stage_inst_dmem_n4801), .A2(MEM_stage_inst_dmem_n4800), .ZN(MEM_stage_inst_dmem_n4802) );
NAND2_X1 MEM_stage_inst_dmem_U4930 ( .A1(MEM_stage_inst_dmem_ram_152), .A2(MEM_stage_inst_dmem_n5807), .ZN(MEM_stage_inst_dmem_n4800) );
NAND2_X1 MEM_stage_inst_dmem_U4929 ( .A1(MEM_stage_inst_dmem_ram_264), .A2(MEM_stage_inst_dmem_n7898), .ZN(MEM_stage_inst_dmem_n4801) );
NAND2_X1 MEM_stage_inst_dmem_U4928 ( .A1(MEM_stage_inst_dmem_n4799), .A2(MEM_stage_inst_dmem_n4798), .ZN(MEM_stage_inst_dmem_n4803) );
NAND2_X1 MEM_stage_inst_dmem_U4927 ( .A1(MEM_stage_inst_dmem_ram_424), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n4798) );
NAND2_X1 MEM_stage_inst_dmem_U4926 ( .A1(MEM_stage_inst_dmem_ram_280), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n4799) );
NOR2_X1 MEM_stage_inst_dmem_U4925 ( .A1(MEM_stage_inst_dmem_n4797), .A2(MEM_stage_inst_dmem_n4796), .ZN(MEM_stage_inst_dmem_n4805) );
NAND2_X1 MEM_stage_inst_dmem_U4924 ( .A1(MEM_stage_inst_dmem_n4795), .A2(MEM_stage_inst_dmem_n4794), .ZN(MEM_stage_inst_dmem_n4796) );
NAND2_X1 MEM_stage_inst_dmem_U4923 ( .A1(MEM_stage_inst_dmem_ram_248), .A2(MEM_stage_inst_dmem_n39), .ZN(MEM_stage_inst_dmem_n4794) );
NAND2_X1 MEM_stage_inst_dmem_U4922 ( .A1(MEM_stage_inst_dmem_ram_8), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n4795) );
NAND2_X1 MEM_stage_inst_dmem_U4921 ( .A1(MEM_stage_inst_dmem_n4793), .A2(MEM_stage_inst_dmem_n4792), .ZN(MEM_stage_inst_dmem_n4797) );
NAND2_X1 MEM_stage_inst_dmem_U4920 ( .A1(MEM_stage_inst_dmem_ram_712), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n4792) );
NAND2_X1 MEM_stage_inst_dmem_U4919 ( .A1(MEM_stage_inst_dmem_ram_72), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n4793) );
NOR2_X1 MEM_stage_inst_dmem_U4918 ( .A1(MEM_stage_inst_dmem_n4791), .A2(MEM_stage_inst_dmem_n8152), .ZN(MEM_stage_inst_dmem_n4920) );
NOR2_X1 MEM_stage_inst_dmem_U4917 ( .A1(MEM_stage_inst_dmem_n4790), .A2(MEM_stage_inst_dmem_n4789), .ZN(MEM_stage_inst_dmem_n4791) );
NAND2_X1 MEM_stage_inst_dmem_U4916 ( .A1(MEM_stage_inst_dmem_n4788), .A2(MEM_stage_inst_dmem_n4787), .ZN(MEM_stage_inst_dmem_n4789) );
NOR2_X1 MEM_stage_inst_dmem_U4915 ( .A1(MEM_stage_inst_dmem_n4786), .A2(MEM_stage_inst_dmem_n4785), .ZN(MEM_stage_inst_dmem_n4787) );
NAND2_X1 MEM_stage_inst_dmem_U4914 ( .A1(MEM_stage_inst_dmem_n4784), .A2(MEM_stage_inst_dmem_n4783), .ZN(MEM_stage_inst_dmem_n4785) );
NOR2_X1 MEM_stage_inst_dmem_U4913 ( .A1(MEM_stage_inst_dmem_n4782), .A2(MEM_stage_inst_dmem_n4781), .ZN(MEM_stage_inst_dmem_n4783) );
NAND2_X1 MEM_stage_inst_dmem_U4912 ( .A1(MEM_stage_inst_dmem_n4780), .A2(MEM_stage_inst_dmem_n4779), .ZN(MEM_stage_inst_dmem_n4781) );
NAND2_X1 MEM_stage_inst_dmem_U4911 ( .A1(MEM_stage_inst_dmem_ram_1176), .A2(MEM_stage_inst_dmem_n5807), .ZN(MEM_stage_inst_dmem_n4779) );
NAND2_X1 MEM_stage_inst_dmem_U4910 ( .A1(MEM_stage_inst_dmem_ram_1752), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n4780) );
NAND2_X1 MEM_stage_inst_dmem_U4909 ( .A1(MEM_stage_inst_dmem_n4778), .A2(MEM_stage_inst_dmem_n4777), .ZN(MEM_stage_inst_dmem_n4782) );
NAND2_X1 MEM_stage_inst_dmem_U4908 ( .A1(MEM_stage_inst_dmem_ram_1224), .A2(MEM_stage_inst_dmem_n36), .ZN(MEM_stage_inst_dmem_n4777) );
NAND2_X1 MEM_stage_inst_dmem_U4907 ( .A1(MEM_stage_inst_dmem_ram_1592), .A2(MEM_stage_inst_dmem_n41), .ZN(MEM_stage_inst_dmem_n4778) );
NOR2_X1 MEM_stage_inst_dmem_U4906 ( .A1(MEM_stage_inst_dmem_n4776), .A2(MEM_stage_inst_dmem_n4775), .ZN(MEM_stage_inst_dmem_n4784) );
NAND2_X1 MEM_stage_inst_dmem_U4905 ( .A1(MEM_stage_inst_dmem_n4774), .A2(MEM_stage_inst_dmem_n4773), .ZN(MEM_stage_inst_dmem_n4775) );
NAND2_X1 MEM_stage_inst_dmem_U4904 ( .A1(MEM_stage_inst_dmem_ram_1448), .A2(MEM_stage_inst_dmem_n4772), .ZN(MEM_stage_inst_dmem_n4773) );
NAND2_X1 MEM_stage_inst_dmem_U4903 ( .A1(MEM_stage_inst_dmem_ram_1192), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n4774) );
NAND2_X1 MEM_stage_inst_dmem_U4902 ( .A1(MEM_stage_inst_dmem_n4771), .A2(MEM_stage_inst_dmem_n4770), .ZN(MEM_stage_inst_dmem_n4776) );
NAND2_X1 MEM_stage_inst_dmem_U4901 ( .A1(MEM_stage_inst_dmem_ram_1976), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n4770) );
NAND2_X1 MEM_stage_inst_dmem_U4900 ( .A1(MEM_stage_inst_dmem_ram_1768), .A2(MEM_stage_inst_dmem_n4769), .ZN(MEM_stage_inst_dmem_n4771) );
NAND2_X1 MEM_stage_inst_dmem_U4899 ( .A1(MEM_stage_inst_dmem_n4768), .A2(MEM_stage_inst_dmem_n4767), .ZN(MEM_stage_inst_dmem_n4786) );
NOR2_X1 MEM_stage_inst_dmem_U4898 ( .A1(MEM_stage_inst_dmem_n4766), .A2(MEM_stage_inst_dmem_n4765), .ZN(MEM_stage_inst_dmem_n4767) );
NAND2_X1 MEM_stage_inst_dmem_U4897 ( .A1(MEM_stage_inst_dmem_n4764), .A2(MEM_stage_inst_dmem_n4763), .ZN(MEM_stage_inst_dmem_n4765) );
NAND2_X1 MEM_stage_inst_dmem_U4896 ( .A1(MEM_stage_inst_dmem_ram_2008), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n4763) );
NAND2_X1 MEM_stage_inst_dmem_U4895 ( .A1(MEM_stage_inst_dmem_ram_1544), .A2(MEM_stage_inst_dmem_n71), .ZN(MEM_stage_inst_dmem_n4764) );
NAND2_X1 MEM_stage_inst_dmem_U4894 ( .A1(MEM_stage_inst_dmem_n4762), .A2(MEM_stage_inst_dmem_n4761), .ZN(MEM_stage_inst_dmem_n4766) );
NAND2_X1 MEM_stage_inst_dmem_U4893 ( .A1(MEM_stage_inst_dmem_ram_1432), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n4761) );
NAND2_X1 MEM_stage_inst_dmem_U4892 ( .A1(MEM_stage_inst_dmem_ram_1064), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n4762) );
NOR2_X1 MEM_stage_inst_dmem_U4891 ( .A1(MEM_stage_inst_dmem_n4760), .A2(MEM_stage_inst_dmem_n4759), .ZN(MEM_stage_inst_dmem_n4768) );
NAND2_X1 MEM_stage_inst_dmem_U4890 ( .A1(MEM_stage_inst_dmem_n4758), .A2(MEM_stage_inst_dmem_n4757), .ZN(MEM_stage_inst_dmem_n4759) );
NAND2_X1 MEM_stage_inst_dmem_U4889 ( .A1(MEM_stage_inst_dmem_ram_1464), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n4757) );
NAND2_X1 MEM_stage_inst_dmem_U4888 ( .A1(MEM_stage_inst_dmem_ram_1256), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n4758) );
NAND2_X1 MEM_stage_inst_dmem_U4887 ( .A1(MEM_stage_inst_dmem_n4756), .A2(MEM_stage_inst_dmem_n4755), .ZN(MEM_stage_inst_dmem_n4760) );
NAND2_X1 MEM_stage_inst_dmem_U4886 ( .A1(MEM_stage_inst_dmem_ram_1944), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n4755) );
NAND2_X1 MEM_stage_inst_dmem_U4885 ( .A1(MEM_stage_inst_dmem_ram_1032), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n4756) );
NOR2_X1 MEM_stage_inst_dmem_U4884 ( .A1(MEM_stage_inst_dmem_n4754), .A2(MEM_stage_inst_dmem_n4753), .ZN(MEM_stage_inst_dmem_n4788) );
NAND2_X1 MEM_stage_inst_dmem_U4883 ( .A1(MEM_stage_inst_dmem_n4752), .A2(MEM_stage_inst_dmem_n4751), .ZN(MEM_stage_inst_dmem_n4753) );
NOR2_X1 MEM_stage_inst_dmem_U4882 ( .A1(MEM_stage_inst_dmem_n4750), .A2(MEM_stage_inst_dmem_n4749), .ZN(MEM_stage_inst_dmem_n4751) );
NAND2_X1 MEM_stage_inst_dmem_U4881 ( .A1(MEM_stage_inst_dmem_n4748), .A2(MEM_stage_inst_dmem_n4747), .ZN(MEM_stage_inst_dmem_n4749) );
NAND2_X1 MEM_stage_inst_dmem_U4880 ( .A1(MEM_stage_inst_dmem_ram_1784), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n4747) );
NAND2_X1 MEM_stage_inst_dmem_U4879 ( .A1(MEM_stage_inst_dmem_ram_1416), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n4748) );
NAND2_X1 MEM_stage_inst_dmem_U4878 ( .A1(MEM_stage_inst_dmem_n4746), .A2(MEM_stage_inst_dmem_n4745), .ZN(MEM_stage_inst_dmem_n4750) );
NAND2_X1 MEM_stage_inst_dmem_U4877 ( .A1(MEM_stage_inst_dmem_ram_1288), .A2(MEM_stage_inst_dmem_n7898), .ZN(MEM_stage_inst_dmem_n4745) );
NAND2_X1 MEM_stage_inst_dmem_U4876 ( .A1(MEM_stage_inst_dmem_ram_1688), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n4746) );
NOR2_X1 MEM_stage_inst_dmem_U4875 ( .A1(MEM_stage_inst_dmem_n4744), .A2(MEM_stage_inst_dmem_n4743), .ZN(MEM_stage_inst_dmem_n4752) );
NAND2_X1 MEM_stage_inst_dmem_U4874 ( .A1(MEM_stage_inst_dmem_n4742), .A2(MEM_stage_inst_dmem_n4741), .ZN(MEM_stage_inst_dmem_n4743) );
NAND2_X1 MEM_stage_inst_dmem_U4873 ( .A1(MEM_stage_inst_dmem_ram_1896), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n4741) );
NAND2_X1 MEM_stage_inst_dmem_U4872 ( .A1(MEM_stage_inst_dmem_ram_1848), .A2(MEM_stage_inst_dmem_n4740), .ZN(MEM_stage_inst_dmem_n4742) );
NAND2_X1 MEM_stage_inst_dmem_U4871 ( .A1(MEM_stage_inst_dmem_n4739), .A2(MEM_stage_inst_dmem_n4738), .ZN(MEM_stage_inst_dmem_n4744) );
NAND2_X1 MEM_stage_inst_dmem_U4870 ( .A1(MEM_stage_inst_dmem_ram_1800), .A2(MEM_stage_inst_dmem_n37), .ZN(MEM_stage_inst_dmem_n4738) );
NAND2_X1 MEM_stage_inst_dmem_U4869 ( .A1(MEM_stage_inst_dmem_ram_1096), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n4739) );
NAND2_X1 MEM_stage_inst_dmem_U4868 ( .A1(MEM_stage_inst_dmem_n4737), .A2(MEM_stage_inst_dmem_n4736), .ZN(MEM_stage_inst_dmem_n4754) );
NOR2_X1 MEM_stage_inst_dmem_U4867 ( .A1(MEM_stage_inst_dmem_n4735), .A2(MEM_stage_inst_dmem_n4734), .ZN(MEM_stage_inst_dmem_n4736) );
NAND2_X1 MEM_stage_inst_dmem_U4866 ( .A1(MEM_stage_inst_dmem_n4733), .A2(MEM_stage_inst_dmem_n4732), .ZN(MEM_stage_inst_dmem_n4734) );
NAND2_X1 MEM_stage_inst_dmem_U4865 ( .A1(MEM_stage_inst_dmem_ram_1336), .A2(MEM_stage_inst_dmem_n4731), .ZN(MEM_stage_inst_dmem_n4732) );
NAND2_X1 MEM_stage_inst_dmem_U4864 ( .A1(MEM_stage_inst_dmem_ram_1480), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n4733) );
NAND2_X1 MEM_stage_inst_dmem_U4863 ( .A1(MEM_stage_inst_dmem_n4730), .A2(MEM_stage_inst_dmem_n4729), .ZN(MEM_stage_inst_dmem_n4735) );
NAND2_X1 MEM_stage_inst_dmem_U4862 ( .A1(MEM_stage_inst_dmem_ram_1992), .A2(MEM_stage_inst_dmem_n4728), .ZN(MEM_stage_inst_dmem_n4729) );
NAND2_X1 MEM_stage_inst_dmem_U4861 ( .A1(MEM_stage_inst_dmem_ram_1320), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n4730) );
NOR2_X1 MEM_stage_inst_dmem_U4860 ( .A1(MEM_stage_inst_dmem_n4727), .A2(MEM_stage_inst_dmem_n4726), .ZN(MEM_stage_inst_dmem_n4737) );
NAND2_X1 MEM_stage_inst_dmem_U4859 ( .A1(MEM_stage_inst_dmem_n4725), .A2(MEM_stage_inst_dmem_n4724), .ZN(MEM_stage_inst_dmem_n4726) );
NAND2_X1 MEM_stage_inst_dmem_U4858 ( .A1(MEM_stage_inst_dmem_ram_1624), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n4724) );
NAND2_X1 MEM_stage_inst_dmem_U4857 ( .A1(MEM_stage_inst_dmem_ram_1608), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n4725) );
NAND2_X1 MEM_stage_inst_dmem_U4856 ( .A1(MEM_stage_inst_dmem_n4723), .A2(MEM_stage_inst_dmem_n4722), .ZN(MEM_stage_inst_dmem_n4727) );
NAND2_X1 MEM_stage_inst_dmem_U4855 ( .A1(MEM_stage_inst_dmem_ram_1368), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n4722) );
NAND2_X1 MEM_stage_inst_dmem_U4854 ( .A1(MEM_stage_inst_dmem_ram_1400), .A2(MEM_stage_inst_dmem_n4721), .ZN(MEM_stage_inst_dmem_n4723) );
NAND2_X1 MEM_stage_inst_dmem_U4853 ( .A1(MEM_stage_inst_dmem_n4720), .A2(MEM_stage_inst_dmem_n4719), .ZN(MEM_stage_inst_dmem_n4790) );
NOR2_X1 MEM_stage_inst_dmem_U4852 ( .A1(MEM_stage_inst_dmem_n4718), .A2(MEM_stage_inst_dmem_n4717), .ZN(MEM_stage_inst_dmem_n4719) );
NAND2_X1 MEM_stage_inst_dmem_U4851 ( .A1(MEM_stage_inst_dmem_n4716), .A2(MEM_stage_inst_dmem_n4715), .ZN(MEM_stage_inst_dmem_n4717) );
NOR2_X1 MEM_stage_inst_dmem_U4850 ( .A1(MEM_stage_inst_dmem_n4714), .A2(MEM_stage_inst_dmem_n4713), .ZN(MEM_stage_inst_dmem_n4715) );
NAND2_X1 MEM_stage_inst_dmem_U4849 ( .A1(MEM_stage_inst_dmem_n4712), .A2(MEM_stage_inst_dmem_n4711), .ZN(MEM_stage_inst_dmem_n4713) );
NAND2_X1 MEM_stage_inst_dmem_U4848 ( .A1(MEM_stage_inst_dmem_ram_1144), .A2(MEM_stage_inst_dmem_n4710), .ZN(MEM_stage_inst_dmem_n4711) );
NAND2_X1 MEM_stage_inst_dmem_U4847 ( .A1(MEM_stage_inst_dmem_ram_1720), .A2(MEM_stage_inst_dmem_n4709), .ZN(MEM_stage_inst_dmem_n4712) );
NAND2_X1 MEM_stage_inst_dmem_U4846 ( .A1(MEM_stage_inst_dmem_n4708), .A2(MEM_stage_inst_dmem_n4707), .ZN(MEM_stage_inst_dmem_n4714) );
NAND2_X1 MEM_stage_inst_dmem_U4845 ( .A1(MEM_stage_inst_dmem_ram_1352), .A2(MEM_stage_inst_dmem_n4706), .ZN(MEM_stage_inst_dmem_n4707) );
NAND2_X1 MEM_stage_inst_dmem_U4844 ( .A1(MEM_stage_inst_dmem_ram_1880), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n4708) );
NOR2_X1 MEM_stage_inst_dmem_U4843 ( .A1(MEM_stage_inst_dmem_n4705), .A2(MEM_stage_inst_dmem_n4704), .ZN(MEM_stage_inst_dmem_n4716) );
NAND2_X1 MEM_stage_inst_dmem_U4842 ( .A1(MEM_stage_inst_dmem_n4703), .A2(MEM_stage_inst_dmem_n4702), .ZN(MEM_stage_inst_dmem_n4704) );
NAND2_X1 MEM_stage_inst_dmem_U4841 ( .A1(MEM_stage_inst_dmem_ram_1528), .A2(MEM_stage_inst_dmem_n64), .ZN(MEM_stage_inst_dmem_n4702) );
NAND2_X1 MEM_stage_inst_dmem_U4840 ( .A1(MEM_stage_inst_dmem_ram_1640), .A2(MEM_stage_inst_dmem_n4701), .ZN(MEM_stage_inst_dmem_n4703) );
NAND2_X1 MEM_stage_inst_dmem_U4839 ( .A1(MEM_stage_inst_dmem_n4700), .A2(MEM_stage_inst_dmem_n4699), .ZN(MEM_stage_inst_dmem_n4705) );
NAND2_X1 MEM_stage_inst_dmem_U4838 ( .A1(MEM_stage_inst_dmem_ram_1384), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n4699) );
NAND2_X1 MEM_stage_inst_dmem_U4837 ( .A1(MEM_stage_inst_dmem_ram_1112), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n4700) );
NAND2_X1 MEM_stage_inst_dmem_U4836 ( .A1(MEM_stage_inst_dmem_n4698), .A2(MEM_stage_inst_dmem_n4697), .ZN(MEM_stage_inst_dmem_n4718) );
NOR2_X1 MEM_stage_inst_dmem_U4835 ( .A1(MEM_stage_inst_dmem_n4696), .A2(MEM_stage_inst_dmem_n4695), .ZN(MEM_stage_inst_dmem_n4697) );
NAND2_X1 MEM_stage_inst_dmem_U4834 ( .A1(MEM_stage_inst_dmem_n4694), .A2(MEM_stage_inst_dmem_n4693), .ZN(MEM_stage_inst_dmem_n4695) );
NAND2_X1 MEM_stage_inst_dmem_U4833 ( .A1(MEM_stage_inst_dmem_ram_1928), .A2(MEM_stage_inst_dmem_n72), .ZN(MEM_stage_inst_dmem_n4693) );
NAND2_X1 MEM_stage_inst_dmem_U4832 ( .A1(MEM_stage_inst_dmem_ram_1576), .A2(MEM_stage_inst_dmem_n4692), .ZN(MEM_stage_inst_dmem_n4694) );
NAND2_X1 MEM_stage_inst_dmem_U4831 ( .A1(MEM_stage_inst_dmem_n4691), .A2(MEM_stage_inst_dmem_n4690), .ZN(MEM_stage_inst_dmem_n4696) );
NAND2_X1 MEM_stage_inst_dmem_U4830 ( .A1(MEM_stage_inst_dmem_ram_1704), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n4690) );
NAND2_X1 MEM_stage_inst_dmem_U4829 ( .A1(MEM_stage_inst_dmem_ram_1128), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n4691) );
NOR2_X1 MEM_stage_inst_dmem_U4828 ( .A1(MEM_stage_inst_dmem_n4689), .A2(MEM_stage_inst_dmem_n4688), .ZN(MEM_stage_inst_dmem_n4698) );
NAND2_X1 MEM_stage_inst_dmem_U4827 ( .A1(MEM_stage_inst_dmem_n4687), .A2(MEM_stage_inst_dmem_n4686), .ZN(MEM_stage_inst_dmem_n4688) );
NAND2_X1 MEM_stage_inst_dmem_U4826 ( .A1(MEM_stage_inst_dmem_ram_1912), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n4686) );
NAND2_X1 MEM_stage_inst_dmem_U4825 ( .A1(MEM_stage_inst_dmem_ram_1864), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n4687) );
NAND2_X1 MEM_stage_inst_dmem_U4824 ( .A1(MEM_stage_inst_dmem_n4685), .A2(MEM_stage_inst_dmem_n4684), .ZN(MEM_stage_inst_dmem_n4689) );
NAND2_X1 MEM_stage_inst_dmem_U4823 ( .A1(MEM_stage_inst_dmem_ram_1240), .A2(MEM_stage_inst_dmem_n51), .ZN(MEM_stage_inst_dmem_n4684) );
NAND2_X1 MEM_stage_inst_dmem_U4822 ( .A1(MEM_stage_inst_dmem_ram_1560), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n4685) );
NOR2_X1 MEM_stage_inst_dmem_U4821 ( .A1(MEM_stage_inst_dmem_n4683), .A2(MEM_stage_inst_dmem_n4682), .ZN(MEM_stage_inst_dmem_n4720) );
NAND2_X1 MEM_stage_inst_dmem_U4820 ( .A1(MEM_stage_inst_dmem_n4681), .A2(MEM_stage_inst_dmem_n4680), .ZN(MEM_stage_inst_dmem_n4682) );
NOR2_X1 MEM_stage_inst_dmem_U4819 ( .A1(MEM_stage_inst_dmem_n4679), .A2(MEM_stage_inst_dmem_n4678), .ZN(MEM_stage_inst_dmem_n4680) );
NAND2_X1 MEM_stage_inst_dmem_U4818 ( .A1(MEM_stage_inst_dmem_n4677), .A2(MEM_stage_inst_dmem_n4676), .ZN(MEM_stage_inst_dmem_n4678) );
NAND2_X1 MEM_stage_inst_dmem_U4817 ( .A1(MEM_stage_inst_dmem_ram_1960), .A2(MEM_stage_inst_dmem_n4675), .ZN(MEM_stage_inst_dmem_n4676) );
NAND2_X1 MEM_stage_inst_dmem_U4816 ( .A1(MEM_stage_inst_dmem_ram_1816), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n4677) );
NAND2_X1 MEM_stage_inst_dmem_U4815 ( .A1(MEM_stage_inst_dmem_n4674), .A2(MEM_stage_inst_dmem_n4673), .ZN(MEM_stage_inst_dmem_n4679) );
NAND2_X1 MEM_stage_inst_dmem_U4814 ( .A1(MEM_stage_inst_dmem_ram_1080), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n4673) );
NAND2_X1 MEM_stage_inst_dmem_U4813 ( .A1(MEM_stage_inst_dmem_ram_1304), .A2(MEM_stage_inst_dmem_n4672), .ZN(MEM_stage_inst_dmem_n4674) );
NOR2_X1 MEM_stage_inst_dmem_U4812 ( .A1(MEM_stage_inst_dmem_n4671), .A2(MEM_stage_inst_dmem_n4670), .ZN(MEM_stage_inst_dmem_n4681) );
NAND2_X1 MEM_stage_inst_dmem_U4811 ( .A1(MEM_stage_inst_dmem_n4669), .A2(MEM_stage_inst_dmem_n4668), .ZN(MEM_stage_inst_dmem_n4670) );
NAND2_X1 MEM_stage_inst_dmem_U4810 ( .A1(MEM_stage_inst_dmem_ram_1512), .A2(MEM_stage_inst_dmem_n4667), .ZN(MEM_stage_inst_dmem_n4668) );
NAND2_X1 MEM_stage_inst_dmem_U4809 ( .A1(MEM_stage_inst_dmem_ram_1208), .A2(MEM_stage_inst_dmem_n55), .ZN(MEM_stage_inst_dmem_n4669) );
NAND2_X1 MEM_stage_inst_dmem_U4808 ( .A1(MEM_stage_inst_dmem_n4666), .A2(MEM_stage_inst_dmem_n4665), .ZN(MEM_stage_inst_dmem_n4671) );
NAND2_X1 MEM_stage_inst_dmem_U4807 ( .A1(MEM_stage_inst_dmem_ram_2024), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n4665) );
NAND2_X1 MEM_stage_inst_dmem_U4806 ( .A1(MEM_stage_inst_dmem_ram_1160), .A2(MEM_stage_inst_dmem_n61), .ZN(MEM_stage_inst_dmem_n4666) );
NAND2_X1 MEM_stage_inst_dmem_U4805 ( .A1(MEM_stage_inst_dmem_n4664), .A2(MEM_stage_inst_dmem_n4663), .ZN(MEM_stage_inst_dmem_n4683) );
NOR2_X1 MEM_stage_inst_dmem_U4804 ( .A1(MEM_stage_inst_dmem_n4662), .A2(MEM_stage_inst_dmem_n4661), .ZN(MEM_stage_inst_dmem_n4663) );
NAND2_X1 MEM_stage_inst_dmem_U4803 ( .A1(MEM_stage_inst_dmem_n4660), .A2(MEM_stage_inst_dmem_n4659), .ZN(MEM_stage_inst_dmem_n4661) );
NAND2_X1 MEM_stage_inst_dmem_U4802 ( .A1(MEM_stage_inst_dmem_ram_1672), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n4659) );
NAND2_X1 MEM_stage_inst_dmem_U4801 ( .A1(MEM_stage_inst_dmem_ram_1496), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n4660) );
NAND2_X1 MEM_stage_inst_dmem_U4800 ( .A1(MEM_stage_inst_dmem_n4658), .A2(MEM_stage_inst_dmem_n4657), .ZN(MEM_stage_inst_dmem_n4662) );
NAND2_X1 MEM_stage_inst_dmem_U4799 ( .A1(MEM_stage_inst_dmem_ram_1832), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n4657) );
NAND2_X1 MEM_stage_inst_dmem_U4798 ( .A1(MEM_stage_inst_dmem_ram_2040), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n4658) );
NOR2_X1 MEM_stage_inst_dmem_U4797 ( .A1(MEM_stage_inst_dmem_n4656), .A2(MEM_stage_inst_dmem_n4655), .ZN(MEM_stage_inst_dmem_n4664) );
NAND2_X1 MEM_stage_inst_dmem_U4796 ( .A1(MEM_stage_inst_dmem_n4654), .A2(MEM_stage_inst_dmem_n4653), .ZN(MEM_stage_inst_dmem_n4655) );
NAND2_X1 MEM_stage_inst_dmem_U4795 ( .A1(MEM_stage_inst_dmem_ram_1048), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n4653) );
NAND2_X1 MEM_stage_inst_dmem_U4794 ( .A1(MEM_stage_inst_dmem_ram_1656), .A2(MEM_stage_inst_dmem_n4652), .ZN(MEM_stage_inst_dmem_n4654) );
NAND2_X1 MEM_stage_inst_dmem_U4793 ( .A1(MEM_stage_inst_dmem_n4651), .A2(MEM_stage_inst_dmem_n4650), .ZN(MEM_stage_inst_dmem_n4656) );
NAND2_X1 MEM_stage_inst_dmem_U4792 ( .A1(MEM_stage_inst_dmem_ram_1736), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n4650) );
NAND2_X1 MEM_stage_inst_dmem_U4791 ( .A1(MEM_stage_inst_dmem_ram_1272), .A2(MEM_stage_inst_dmem_n4649), .ZN(MEM_stage_inst_dmem_n4651) );
NOR2_X1 MEM_stage_inst_dmem_U4790 ( .A1(MEM_stage_inst_dmem_n4648), .A2(MEM_stage_inst_dmem_n4647), .ZN(MEM_stage_inst_dmem_n4922) );
NOR2_X1 MEM_stage_inst_dmem_U4789 ( .A1(MEM_stage_inst_dmem_n4646), .A2(MEM_stage_inst_dmem_n8417), .ZN(MEM_stage_inst_dmem_n4647) );
NOR2_X1 MEM_stage_inst_dmem_U4788 ( .A1(MEM_stage_inst_dmem_n4645), .A2(MEM_stage_inst_dmem_n4644), .ZN(MEM_stage_inst_dmem_n4646) );
NAND2_X1 MEM_stage_inst_dmem_U4787 ( .A1(MEM_stage_inst_dmem_n4643), .A2(MEM_stage_inst_dmem_n4642), .ZN(MEM_stage_inst_dmem_n4644) );
NOR2_X1 MEM_stage_inst_dmem_U4786 ( .A1(MEM_stage_inst_dmem_n4641), .A2(MEM_stage_inst_dmem_n4640), .ZN(MEM_stage_inst_dmem_n4642) );
NAND2_X1 MEM_stage_inst_dmem_U4785 ( .A1(MEM_stage_inst_dmem_n4639), .A2(MEM_stage_inst_dmem_n4638), .ZN(MEM_stage_inst_dmem_n4640) );
NOR2_X1 MEM_stage_inst_dmem_U4784 ( .A1(MEM_stage_inst_dmem_n4637), .A2(MEM_stage_inst_dmem_n4636), .ZN(MEM_stage_inst_dmem_n4638) );
NAND2_X1 MEM_stage_inst_dmem_U4783 ( .A1(MEM_stage_inst_dmem_n4635), .A2(MEM_stage_inst_dmem_n4634), .ZN(MEM_stage_inst_dmem_n4636) );
NAND2_X1 MEM_stage_inst_dmem_U4782 ( .A1(MEM_stage_inst_dmem_ram_3432), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n4634) );
NAND2_X1 MEM_stage_inst_dmem_U4781 ( .A1(MEM_stage_inst_dmem_ram_3080), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n4635) );
NAND2_X1 MEM_stage_inst_dmem_U4780 ( .A1(MEM_stage_inst_dmem_n4633), .A2(MEM_stage_inst_dmem_n4632), .ZN(MEM_stage_inst_dmem_n4637) );
NAND2_X1 MEM_stage_inst_dmem_U4779 ( .A1(MEM_stage_inst_dmem_ram_3576), .A2(MEM_stage_inst_dmem_n64), .ZN(MEM_stage_inst_dmem_n4632) );
NAND2_X1 MEM_stage_inst_dmem_U4778 ( .A1(MEM_stage_inst_dmem_ram_3880), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n4633) );
NOR2_X1 MEM_stage_inst_dmem_U4777 ( .A1(MEM_stage_inst_dmem_n4631), .A2(MEM_stage_inst_dmem_n4630), .ZN(MEM_stage_inst_dmem_n4639) );
NAND2_X1 MEM_stage_inst_dmem_U4776 ( .A1(MEM_stage_inst_dmem_n4629), .A2(MEM_stage_inst_dmem_n4628), .ZN(MEM_stage_inst_dmem_n4630) );
NAND2_X1 MEM_stage_inst_dmem_U4775 ( .A1(MEM_stage_inst_dmem_ram_3848), .A2(MEM_stage_inst_dmem_n37), .ZN(MEM_stage_inst_dmem_n4628) );
NAND2_X1 MEM_stage_inst_dmem_U4774 ( .A1(MEM_stage_inst_dmem_ram_3608), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n4629) );
NAND2_X1 MEM_stage_inst_dmem_U4773 ( .A1(MEM_stage_inst_dmem_n4627), .A2(MEM_stage_inst_dmem_n4626), .ZN(MEM_stage_inst_dmem_n4631) );
NAND2_X1 MEM_stage_inst_dmem_U4772 ( .A1(MEM_stage_inst_dmem_ram_4072), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n4626) );
NAND2_X1 MEM_stage_inst_dmem_U4771 ( .A1(MEM_stage_inst_dmem_ram_3768), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n4627) );
NAND2_X1 MEM_stage_inst_dmem_U4770 ( .A1(MEM_stage_inst_dmem_n4625), .A2(MEM_stage_inst_dmem_n4624), .ZN(MEM_stage_inst_dmem_n4641) );
NOR2_X1 MEM_stage_inst_dmem_U4769 ( .A1(MEM_stage_inst_dmem_n4623), .A2(MEM_stage_inst_dmem_n4622), .ZN(MEM_stage_inst_dmem_n4624) );
NAND2_X1 MEM_stage_inst_dmem_U4768 ( .A1(MEM_stage_inst_dmem_n4621), .A2(MEM_stage_inst_dmem_n4620), .ZN(MEM_stage_inst_dmem_n4622) );
NAND2_X1 MEM_stage_inst_dmem_U4767 ( .A1(MEM_stage_inst_dmem_ram_3720), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n4620) );
NAND2_X1 MEM_stage_inst_dmem_U4766 ( .A1(MEM_stage_inst_dmem_ram_3224), .A2(MEM_stage_inst_dmem_n5807), .ZN(MEM_stage_inst_dmem_n4621) );
NAND2_X1 MEM_stage_inst_dmem_U4765 ( .A1(MEM_stage_inst_dmem_n4619), .A2(MEM_stage_inst_dmem_n4618), .ZN(MEM_stage_inst_dmem_n4623) );
NAND2_X1 MEM_stage_inst_dmem_U4764 ( .A1(MEM_stage_inst_dmem_ram_3736), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n4618) );
NAND2_X1 MEM_stage_inst_dmem_U4763 ( .A1(MEM_stage_inst_dmem_ram_3816), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n4619) );
NOR2_X1 MEM_stage_inst_dmem_U4762 ( .A1(MEM_stage_inst_dmem_n4617), .A2(MEM_stage_inst_dmem_n4616), .ZN(MEM_stage_inst_dmem_n4625) );
NAND2_X1 MEM_stage_inst_dmem_U4761 ( .A1(MEM_stage_inst_dmem_n4615), .A2(MEM_stage_inst_dmem_n4614), .ZN(MEM_stage_inst_dmem_n4616) );
NAND2_X1 MEM_stage_inst_dmem_U4760 ( .A1(MEM_stage_inst_dmem_ram_3752), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n4614) );
NAND2_X1 MEM_stage_inst_dmem_U4759 ( .A1(MEM_stage_inst_dmem_ram_3704), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n4615) );
NAND2_X1 MEM_stage_inst_dmem_U4758 ( .A1(MEM_stage_inst_dmem_n4613), .A2(MEM_stage_inst_dmem_n4612), .ZN(MEM_stage_inst_dmem_n4617) );
NAND2_X1 MEM_stage_inst_dmem_U4757 ( .A1(MEM_stage_inst_dmem_ram_3480), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n4612) );
NAND2_X1 MEM_stage_inst_dmem_U4756 ( .A1(MEM_stage_inst_dmem_ram_4008), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n4613) );
NOR2_X1 MEM_stage_inst_dmem_U4755 ( .A1(MEM_stage_inst_dmem_n4611), .A2(MEM_stage_inst_dmem_n4610), .ZN(MEM_stage_inst_dmem_n4643) );
NAND2_X1 MEM_stage_inst_dmem_U4754 ( .A1(MEM_stage_inst_dmem_n4609), .A2(MEM_stage_inst_dmem_n4608), .ZN(MEM_stage_inst_dmem_n4610) );
NOR2_X1 MEM_stage_inst_dmem_U4753 ( .A1(MEM_stage_inst_dmem_n4607), .A2(MEM_stage_inst_dmem_n4606), .ZN(MEM_stage_inst_dmem_n4608) );
NAND2_X1 MEM_stage_inst_dmem_U4752 ( .A1(MEM_stage_inst_dmem_n4605), .A2(MEM_stage_inst_dmem_n4604), .ZN(MEM_stage_inst_dmem_n4606) );
NAND2_X1 MEM_stage_inst_dmem_U4751 ( .A1(MEM_stage_inst_dmem_ram_3256), .A2(MEM_stage_inst_dmem_n55), .ZN(MEM_stage_inst_dmem_n4604) );
NAND2_X1 MEM_stage_inst_dmem_U4750 ( .A1(MEM_stage_inst_dmem_ram_3800), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n4605) );
NAND2_X1 MEM_stage_inst_dmem_U4749 ( .A1(MEM_stage_inst_dmem_n4603), .A2(MEM_stage_inst_dmem_n4602), .ZN(MEM_stage_inst_dmem_n4607) );
NAND2_X1 MEM_stage_inst_dmem_U4748 ( .A1(MEM_stage_inst_dmem_ram_3624), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n4602) );
NAND2_X1 MEM_stage_inst_dmem_U4747 ( .A1(MEM_stage_inst_dmem_ram_3192), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n4603) );
NOR2_X1 MEM_stage_inst_dmem_U4746 ( .A1(MEM_stage_inst_dmem_n4601), .A2(MEM_stage_inst_dmem_n4600), .ZN(MEM_stage_inst_dmem_n4609) );
NAND2_X1 MEM_stage_inst_dmem_U4745 ( .A1(MEM_stage_inst_dmem_n4599), .A2(MEM_stage_inst_dmem_n4598), .ZN(MEM_stage_inst_dmem_n4600) );
NAND2_X1 MEM_stage_inst_dmem_U4744 ( .A1(MEM_stage_inst_dmem_ram_3496), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n4598) );
NAND2_X1 MEM_stage_inst_dmem_U4743 ( .A1(MEM_stage_inst_dmem_ram_3352), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n4599) );
NAND2_X1 MEM_stage_inst_dmem_U4742 ( .A1(MEM_stage_inst_dmem_n4597), .A2(MEM_stage_inst_dmem_n4596), .ZN(MEM_stage_inst_dmem_n4601) );
NAND2_X1 MEM_stage_inst_dmem_U4741 ( .A1(MEM_stage_inst_dmem_ram_4040), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n4596) );
NAND2_X1 MEM_stage_inst_dmem_U4740 ( .A1(MEM_stage_inst_dmem_ram_3864), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n4597) );
NAND2_X1 MEM_stage_inst_dmem_U4739 ( .A1(MEM_stage_inst_dmem_n4595), .A2(MEM_stage_inst_dmem_n4594), .ZN(MEM_stage_inst_dmem_n4611) );
NOR2_X1 MEM_stage_inst_dmem_U4738 ( .A1(MEM_stage_inst_dmem_n4593), .A2(MEM_stage_inst_dmem_n4592), .ZN(MEM_stage_inst_dmem_n4594) );
NAND2_X1 MEM_stage_inst_dmem_U4737 ( .A1(MEM_stage_inst_dmem_n4591), .A2(MEM_stage_inst_dmem_n4590), .ZN(MEM_stage_inst_dmem_n4592) );
NAND2_X1 MEM_stage_inst_dmem_U4736 ( .A1(MEM_stage_inst_dmem_ram_3688), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n4590) );
NAND2_X1 MEM_stage_inst_dmem_U4735 ( .A1(MEM_stage_inst_dmem_ram_3672), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n4591) );
NAND2_X1 MEM_stage_inst_dmem_U4734 ( .A1(MEM_stage_inst_dmem_n4589), .A2(MEM_stage_inst_dmem_n4588), .ZN(MEM_stage_inst_dmem_n4593) );
NAND2_X1 MEM_stage_inst_dmem_U4733 ( .A1(MEM_stage_inst_dmem_ram_3304), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n4588) );
NAND2_X1 MEM_stage_inst_dmem_U4732 ( .A1(MEM_stage_inst_dmem_ram_3416), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n4589) );
NOR2_X1 MEM_stage_inst_dmem_U4731 ( .A1(MEM_stage_inst_dmem_n4587), .A2(MEM_stage_inst_dmem_n4586), .ZN(MEM_stage_inst_dmem_n4595) );
NAND2_X1 MEM_stage_inst_dmem_U4730 ( .A1(MEM_stage_inst_dmem_n4585), .A2(MEM_stage_inst_dmem_n4584), .ZN(MEM_stage_inst_dmem_n4586) );
NAND2_X1 MEM_stage_inst_dmem_U4729 ( .A1(MEM_stage_inst_dmem_ram_3128), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n4584) );
NAND2_X1 MEM_stage_inst_dmem_U4728 ( .A1(MEM_stage_inst_dmem_ram_3368), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n4585) );
NAND2_X1 MEM_stage_inst_dmem_U4727 ( .A1(MEM_stage_inst_dmem_n4583), .A2(MEM_stage_inst_dmem_n4582), .ZN(MEM_stage_inst_dmem_n4587) );
NAND2_X1 MEM_stage_inst_dmem_U4726 ( .A1(MEM_stage_inst_dmem_ram_3464), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n4582) );
NAND2_X1 MEM_stage_inst_dmem_U4725 ( .A1(MEM_stage_inst_dmem_ram_3240), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n4583) );
NAND2_X1 MEM_stage_inst_dmem_U4724 ( .A1(MEM_stage_inst_dmem_n4581), .A2(MEM_stage_inst_dmem_n4580), .ZN(MEM_stage_inst_dmem_n4645) );
NOR2_X1 MEM_stage_inst_dmem_U4723 ( .A1(MEM_stage_inst_dmem_n4579), .A2(MEM_stage_inst_dmem_n4578), .ZN(MEM_stage_inst_dmem_n4580) );
NAND2_X1 MEM_stage_inst_dmem_U4722 ( .A1(MEM_stage_inst_dmem_n4577), .A2(MEM_stage_inst_dmem_n4576), .ZN(MEM_stage_inst_dmem_n4578) );
NOR2_X1 MEM_stage_inst_dmem_U4721 ( .A1(MEM_stage_inst_dmem_n4575), .A2(MEM_stage_inst_dmem_n4574), .ZN(MEM_stage_inst_dmem_n4576) );
NAND2_X1 MEM_stage_inst_dmem_U4720 ( .A1(MEM_stage_inst_dmem_n4573), .A2(MEM_stage_inst_dmem_n4572), .ZN(MEM_stage_inst_dmem_n4574) );
NAND2_X1 MEM_stage_inst_dmem_U4719 ( .A1(MEM_stage_inst_dmem_ram_3912), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n4572) );
NAND2_X1 MEM_stage_inst_dmem_U4718 ( .A1(MEM_stage_inst_dmem_ram_3208), .A2(MEM_stage_inst_dmem_n61), .ZN(MEM_stage_inst_dmem_n4573) );
NAND2_X1 MEM_stage_inst_dmem_U4717 ( .A1(MEM_stage_inst_dmem_n4571), .A2(MEM_stage_inst_dmem_n4570), .ZN(MEM_stage_inst_dmem_n4575) );
NAND2_X1 MEM_stage_inst_dmem_U4716 ( .A1(MEM_stage_inst_dmem_ram_3144), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n4570) );
NAND2_X1 MEM_stage_inst_dmem_U4715 ( .A1(MEM_stage_inst_dmem_ram_3320), .A2(MEM_stage_inst_dmem_n39), .ZN(MEM_stage_inst_dmem_n4571) );
NOR2_X1 MEM_stage_inst_dmem_U4714 ( .A1(MEM_stage_inst_dmem_n4569), .A2(MEM_stage_inst_dmem_n4568), .ZN(MEM_stage_inst_dmem_n4577) );
NAND2_X1 MEM_stage_inst_dmem_U4713 ( .A1(MEM_stage_inst_dmem_n4567), .A2(MEM_stage_inst_dmem_n4566), .ZN(MEM_stage_inst_dmem_n4568) );
NAND2_X1 MEM_stage_inst_dmem_U4712 ( .A1(MEM_stage_inst_dmem_ram_3160), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n4566) );
NAND2_X1 MEM_stage_inst_dmem_U4711 ( .A1(MEM_stage_inst_dmem_ram_3592), .A2(MEM_stage_inst_dmem_n71), .ZN(MEM_stage_inst_dmem_n4567) );
NAND2_X1 MEM_stage_inst_dmem_U4710 ( .A1(MEM_stage_inst_dmem_n4565), .A2(MEM_stage_inst_dmem_n4564), .ZN(MEM_stage_inst_dmem_n4569) );
NAND2_X1 MEM_stage_inst_dmem_U4709 ( .A1(MEM_stage_inst_dmem_ram_4024), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n4564) );
NAND2_X1 MEM_stage_inst_dmem_U4708 ( .A1(MEM_stage_inst_dmem_ram_3544), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n4565) );
NAND2_X1 MEM_stage_inst_dmem_U4707 ( .A1(MEM_stage_inst_dmem_n4563), .A2(MEM_stage_inst_dmem_n4562), .ZN(MEM_stage_inst_dmem_n4579) );
NOR2_X1 MEM_stage_inst_dmem_U4706 ( .A1(MEM_stage_inst_dmem_n4561), .A2(MEM_stage_inst_dmem_n4560), .ZN(MEM_stage_inst_dmem_n4562) );
NAND2_X1 MEM_stage_inst_dmem_U4705 ( .A1(MEM_stage_inst_dmem_n4559), .A2(MEM_stage_inst_dmem_n4558), .ZN(MEM_stage_inst_dmem_n4560) );
NAND2_X1 MEM_stage_inst_dmem_U4704 ( .A1(MEM_stage_inst_dmem_ram_3928), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n4558) );
NAND2_X1 MEM_stage_inst_dmem_U4703 ( .A1(MEM_stage_inst_dmem_ram_3992), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n4559) );
NAND2_X1 MEM_stage_inst_dmem_U4702 ( .A1(MEM_stage_inst_dmem_n4557), .A2(MEM_stage_inst_dmem_n4556), .ZN(MEM_stage_inst_dmem_n4561) );
NAND2_X1 MEM_stage_inst_dmem_U4701 ( .A1(MEM_stage_inst_dmem_ram_3944), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n4556) );
NAND2_X1 MEM_stage_inst_dmem_U4700 ( .A1(MEM_stage_inst_dmem_ram_3096), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n4557) );
NOR2_X1 MEM_stage_inst_dmem_U4699 ( .A1(MEM_stage_inst_dmem_n4555), .A2(MEM_stage_inst_dmem_n4554), .ZN(MEM_stage_inst_dmem_n4563) );
NAND2_X1 MEM_stage_inst_dmem_U4698 ( .A1(MEM_stage_inst_dmem_n4553), .A2(MEM_stage_inst_dmem_n4552), .ZN(MEM_stage_inst_dmem_n4554) );
NAND2_X1 MEM_stage_inst_dmem_U4697 ( .A1(MEM_stage_inst_dmem_ram_3784), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n4552) );
NAND2_X1 MEM_stage_inst_dmem_U4696 ( .A1(MEM_stage_inst_dmem_ram_3832), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n4553) );
NAND2_X1 MEM_stage_inst_dmem_U4695 ( .A1(MEM_stage_inst_dmem_n4551), .A2(MEM_stage_inst_dmem_n4550), .ZN(MEM_stage_inst_dmem_n4555) );
NAND2_X1 MEM_stage_inst_dmem_U4694 ( .A1(MEM_stage_inst_dmem_ram_3960), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n4550) );
NAND2_X1 MEM_stage_inst_dmem_U4693 ( .A1(MEM_stage_inst_dmem_ram_3976), .A2(MEM_stage_inst_dmem_n72), .ZN(MEM_stage_inst_dmem_n4551) );
NOR2_X1 MEM_stage_inst_dmem_U4692 ( .A1(MEM_stage_inst_dmem_n4549), .A2(MEM_stage_inst_dmem_n4548), .ZN(MEM_stage_inst_dmem_n4581) );
NAND2_X1 MEM_stage_inst_dmem_U4691 ( .A1(MEM_stage_inst_dmem_n4547), .A2(MEM_stage_inst_dmem_n4546), .ZN(MEM_stage_inst_dmem_n4548) );
NOR2_X1 MEM_stage_inst_dmem_U4690 ( .A1(MEM_stage_inst_dmem_n4545), .A2(MEM_stage_inst_dmem_n4544), .ZN(MEM_stage_inst_dmem_n4546) );
NAND2_X1 MEM_stage_inst_dmem_U4689 ( .A1(MEM_stage_inst_dmem_n4543), .A2(MEM_stage_inst_dmem_n4542), .ZN(MEM_stage_inst_dmem_n4544) );
NAND2_X1 MEM_stage_inst_dmem_U4688 ( .A1(MEM_stage_inst_dmem_ram_3512), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n4542) );
NAND2_X1 MEM_stage_inst_dmem_U4687 ( .A1(MEM_stage_inst_dmem_ram_3336), .A2(MEM_stage_inst_dmem_n7898), .ZN(MEM_stage_inst_dmem_n4543) );
NAND2_X1 MEM_stage_inst_dmem_U4686 ( .A1(MEM_stage_inst_dmem_n4541), .A2(MEM_stage_inst_dmem_n4540), .ZN(MEM_stage_inst_dmem_n4545) );
NAND2_X1 MEM_stage_inst_dmem_U4685 ( .A1(MEM_stage_inst_dmem_ram_3400), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n4540) );
NAND2_X1 MEM_stage_inst_dmem_U4684 ( .A1(MEM_stage_inst_dmem_ram_3384), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n4541) );
NOR2_X1 MEM_stage_inst_dmem_U4683 ( .A1(MEM_stage_inst_dmem_n4539), .A2(MEM_stage_inst_dmem_n4538), .ZN(MEM_stage_inst_dmem_n4547) );
NAND2_X1 MEM_stage_inst_dmem_U4682 ( .A1(MEM_stage_inst_dmem_n4537), .A2(MEM_stage_inst_dmem_n4536), .ZN(MEM_stage_inst_dmem_n4538) );
NAND2_X1 MEM_stage_inst_dmem_U4681 ( .A1(MEM_stage_inst_dmem_ram_4056), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n4536) );
NAND2_X1 MEM_stage_inst_dmem_U4680 ( .A1(MEM_stage_inst_dmem_ram_3448), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n4537) );
NAND2_X1 MEM_stage_inst_dmem_U4679 ( .A1(MEM_stage_inst_dmem_n4535), .A2(MEM_stage_inst_dmem_n4534), .ZN(MEM_stage_inst_dmem_n4539) );
NAND2_X1 MEM_stage_inst_dmem_U4678 ( .A1(MEM_stage_inst_dmem_ram_3896), .A2(MEM_stage_inst_dmem_n46), .ZN(MEM_stage_inst_dmem_n4534) );
NAND2_X1 MEM_stage_inst_dmem_U4677 ( .A1(MEM_stage_inst_dmem_ram_4088), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n4535) );
NAND2_X1 MEM_stage_inst_dmem_U4676 ( .A1(MEM_stage_inst_dmem_n4533), .A2(MEM_stage_inst_dmem_n4532), .ZN(MEM_stage_inst_dmem_n4549) );
NOR2_X1 MEM_stage_inst_dmem_U4675 ( .A1(MEM_stage_inst_dmem_n4531), .A2(MEM_stage_inst_dmem_n4530), .ZN(MEM_stage_inst_dmem_n4532) );
NAND2_X1 MEM_stage_inst_dmem_U4674 ( .A1(MEM_stage_inst_dmem_n4529), .A2(MEM_stage_inst_dmem_n4528), .ZN(MEM_stage_inst_dmem_n4530) );
NAND2_X1 MEM_stage_inst_dmem_U4673 ( .A1(MEM_stage_inst_dmem_ram_3272), .A2(MEM_stage_inst_dmem_n36), .ZN(MEM_stage_inst_dmem_n4528) );
NAND2_X1 MEM_stage_inst_dmem_U4672 ( .A1(MEM_stage_inst_dmem_ram_3528), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n4529) );
NAND2_X1 MEM_stage_inst_dmem_U4671 ( .A1(MEM_stage_inst_dmem_n4527), .A2(MEM_stage_inst_dmem_n4526), .ZN(MEM_stage_inst_dmem_n4531) );
NAND2_X1 MEM_stage_inst_dmem_U4670 ( .A1(MEM_stage_inst_dmem_ram_3112), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n4526) );
NAND2_X1 MEM_stage_inst_dmem_U4669 ( .A1(MEM_stage_inst_dmem_ram_3656), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n4527) );
NOR2_X1 MEM_stage_inst_dmem_U4668 ( .A1(MEM_stage_inst_dmem_n4525), .A2(MEM_stage_inst_dmem_n4524), .ZN(MEM_stage_inst_dmem_n4533) );
NAND2_X1 MEM_stage_inst_dmem_U4667 ( .A1(MEM_stage_inst_dmem_n4523), .A2(MEM_stage_inst_dmem_n4522), .ZN(MEM_stage_inst_dmem_n4524) );
NAND2_X1 MEM_stage_inst_dmem_U4666 ( .A1(MEM_stage_inst_dmem_ram_3640), .A2(MEM_stage_inst_dmem_n41), .ZN(MEM_stage_inst_dmem_n4522) );
NAND2_X1 MEM_stage_inst_dmem_U4665 ( .A1(MEM_stage_inst_dmem_ram_3560), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n4523) );
NAND2_X1 MEM_stage_inst_dmem_U4664 ( .A1(MEM_stage_inst_dmem_n4521), .A2(MEM_stage_inst_dmem_n4520), .ZN(MEM_stage_inst_dmem_n4525) );
NAND2_X1 MEM_stage_inst_dmem_U4663 ( .A1(MEM_stage_inst_dmem_ram_3288), .A2(MEM_stage_inst_dmem_n51), .ZN(MEM_stage_inst_dmem_n4520) );
NAND2_X1 MEM_stage_inst_dmem_U4662 ( .A1(MEM_stage_inst_dmem_ram_3176), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n4521) );
NOR2_X1 MEM_stage_inst_dmem_U4661 ( .A1(MEM_stage_inst_dmem_n4519), .A2(MEM_stage_inst_dmem_n8286), .ZN(MEM_stage_inst_dmem_n4648) );
NOR2_X1 MEM_stage_inst_dmem_U4660 ( .A1(MEM_stage_inst_dmem_n4518), .A2(MEM_stage_inst_dmem_n4517), .ZN(MEM_stage_inst_dmem_n4519) );
NAND2_X1 MEM_stage_inst_dmem_U4659 ( .A1(MEM_stage_inst_dmem_n4516), .A2(MEM_stage_inst_dmem_n4515), .ZN(MEM_stage_inst_dmem_n4517) );
NOR2_X1 MEM_stage_inst_dmem_U4658 ( .A1(MEM_stage_inst_dmem_n4514), .A2(MEM_stage_inst_dmem_n4513), .ZN(MEM_stage_inst_dmem_n4515) );
NAND2_X1 MEM_stage_inst_dmem_U4657 ( .A1(MEM_stage_inst_dmem_n4512), .A2(MEM_stage_inst_dmem_n4511), .ZN(MEM_stage_inst_dmem_n4513) );
NOR2_X1 MEM_stage_inst_dmem_U4656 ( .A1(MEM_stage_inst_dmem_n4510), .A2(MEM_stage_inst_dmem_n4509), .ZN(MEM_stage_inst_dmem_n4511) );
NAND2_X1 MEM_stage_inst_dmem_U4655 ( .A1(MEM_stage_inst_dmem_n4508), .A2(MEM_stage_inst_dmem_n4507), .ZN(MEM_stage_inst_dmem_n4509) );
NAND2_X1 MEM_stage_inst_dmem_U4654 ( .A1(MEM_stage_inst_dmem_ram_2168), .A2(MEM_stage_inst_dmem_n4710), .ZN(MEM_stage_inst_dmem_n4507) );
NAND2_X1 MEM_stage_inst_dmem_U4653 ( .A1(MEM_stage_inst_dmem_ram_2216), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n4508) );
NAND2_X1 MEM_stage_inst_dmem_U4652 ( .A1(MEM_stage_inst_dmem_n4506), .A2(MEM_stage_inst_dmem_n4505), .ZN(MEM_stage_inst_dmem_n4510) );
NAND2_X1 MEM_stage_inst_dmem_U4651 ( .A1(MEM_stage_inst_dmem_ram_2104), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n4505) );
NAND2_X1 MEM_stage_inst_dmem_U4650 ( .A1(MEM_stage_inst_dmem_ram_2792), .A2(MEM_stage_inst_dmem_n4769), .ZN(MEM_stage_inst_dmem_n4506) );
NOR2_X1 MEM_stage_inst_dmem_U4649 ( .A1(MEM_stage_inst_dmem_n4504), .A2(MEM_stage_inst_dmem_n4503), .ZN(MEM_stage_inst_dmem_n4512) );
NAND2_X1 MEM_stage_inst_dmem_U4648 ( .A1(MEM_stage_inst_dmem_n4502), .A2(MEM_stage_inst_dmem_n4501), .ZN(MEM_stage_inst_dmem_n4503) );
NAND2_X1 MEM_stage_inst_dmem_U4647 ( .A1(MEM_stage_inst_dmem_ram_2296), .A2(MEM_stage_inst_dmem_n4649), .ZN(MEM_stage_inst_dmem_n4501) );
NAND2_X1 MEM_stage_inst_dmem_U4646 ( .A1(MEM_stage_inst_dmem_ram_2440), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n4502) );
NAND2_X1 MEM_stage_inst_dmem_U4645 ( .A1(MEM_stage_inst_dmem_n4500), .A2(MEM_stage_inst_dmem_n4499), .ZN(MEM_stage_inst_dmem_n4504) );
NAND2_X1 MEM_stage_inst_dmem_U4644 ( .A1(MEM_stage_inst_dmem_ram_2616), .A2(MEM_stage_inst_dmem_n41), .ZN(MEM_stage_inst_dmem_n4499) );
NAND2_X1 MEM_stage_inst_dmem_U4643 ( .A1(MEM_stage_inst_dmem_ram_2648), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n4500) );
NAND2_X1 MEM_stage_inst_dmem_U4642 ( .A1(MEM_stage_inst_dmem_n4498), .A2(MEM_stage_inst_dmem_n4497), .ZN(MEM_stage_inst_dmem_n4514) );
NOR2_X1 MEM_stage_inst_dmem_U4641 ( .A1(MEM_stage_inst_dmem_n4496), .A2(MEM_stage_inst_dmem_n4495), .ZN(MEM_stage_inst_dmem_n4497) );
NAND2_X1 MEM_stage_inst_dmem_U4640 ( .A1(MEM_stage_inst_dmem_n4494), .A2(MEM_stage_inst_dmem_n4493), .ZN(MEM_stage_inst_dmem_n4495) );
NAND2_X1 MEM_stage_inst_dmem_U4639 ( .A1(MEM_stage_inst_dmem_ram_2120), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n4493) );
NAND2_X1 MEM_stage_inst_dmem_U4638 ( .A1(MEM_stage_inst_dmem_ram_2712), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n4494) );
NAND2_X1 MEM_stage_inst_dmem_U4637 ( .A1(MEM_stage_inst_dmem_n4492), .A2(MEM_stage_inst_dmem_n4491), .ZN(MEM_stage_inst_dmem_n4496) );
NAND2_X1 MEM_stage_inst_dmem_U4636 ( .A1(MEM_stage_inst_dmem_ram_2952), .A2(MEM_stage_inst_dmem_n72), .ZN(MEM_stage_inst_dmem_n4491) );
NAND2_X1 MEM_stage_inst_dmem_U4635 ( .A1(MEM_stage_inst_dmem_ram_2200), .A2(MEM_stage_inst_dmem_n44), .ZN(MEM_stage_inst_dmem_n4492) );
NOR2_X1 MEM_stage_inst_dmem_U4634 ( .A1(MEM_stage_inst_dmem_n4490), .A2(MEM_stage_inst_dmem_n4489), .ZN(MEM_stage_inst_dmem_n4498) );
NAND2_X1 MEM_stage_inst_dmem_U4633 ( .A1(MEM_stage_inst_dmem_n4488), .A2(MEM_stage_inst_dmem_n4487), .ZN(MEM_stage_inst_dmem_n4489) );
NAND2_X1 MEM_stage_inst_dmem_U4632 ( .A1(MEM_stage_inst_dmem_ram_2072), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n4487) );
NAND2_X1 MEM_stage_inst_dmem_U4631 ( .A1(MEM_stage_inst_dmem_ram_2568), .A2(MEM_stage_inst_dmem_n71), .ZN(MEM_stage_inst_dmem_n4488) );
NAND2_X1 MEM_stage_inst_dmem_U4630 ( .A1(MEM_stage_inst_dmem_n4486), .A2(MEM_stage_inst_dmem_n4485), .ZN(MEM_stage_inst_dmem_n4490) );
NAND2_X1 MEM_stage_inst_dmem_U4629 ( .A1(MEM_stage_inst_dmem_ram_2872), .A2(MEM_stage_inst_dmem_n4740), .ZN(MEM_stage_inst_dmem_n4485) );
NAND2_X1 MEM_stage_inst_dmem_U4628 ( .A1(MEM_stage_inst_dmem_ram_2424), .A2(MEM_stage_inst_dmem_n4721), .ZN(MEM_stage_inst_dmem_n4486) );
NOR2_X1 MEM_stage_inst_dmem_U4627 ( .A1(MEM_stage_inst_dmem_n4484), .A2(MEM_stage_inst_dmem_n4483), .ZN(MEM_stage_inst_dmem_n4516) );
NAND2_X1 MEM_stage_inst_dmem_U4626 ( .A1(MEM_stage_inst_dmem_n4482), .A2(MEM_stage_inst_dmem_n4481), .ZN(MEM_stage_inst_dmem_n4483) );
NOR2_X1 MEM_stage_inst_dmem_U4625 ( .A1(MEM_stage_inst_dmem_n4480), .A2(MEM_stage_inst_dmem_n4479), .ZN(MEM_stage_inst_dmem_n4481) );
NAND2_X1 MEM_stage_inst_dmem_U4624 ( .A1(MEM_stage_inst_dmem_n4478), .A2(MEM_stage_inst_dmem_n4477), .ZN(MEM_stage_inst_dmem_n4479) );
NAND2_X1 MEM_stage_inst_dmem_U4623 ( .A1(MEM_stage_inst_dmem_ram_2088), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n4477) );
NAND2_X1 MEM_stage_inst_dmem_U4622 ( .A1(MEM_stage_inst_dmem_ram_2664), .A2(MEM_stage_inst_dmem_n4701), .ZN(MEM_stage_inst_dmem_n4478) );
NAND2_X1 MEM_stage_inst_dmem_U4621 ( .A1(MEM_stage_inst_dmem_n4476), .A2(MEM_stage_inst_dmem_n4475), .ZN(MEM_stage_inst_dmem_n4480) );
NAND2_X1 MEM_stage_inst_dmem_U4620 ( .A1(MEM_stage_inst_dmem_ram_2760), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n4475) );
NAND2_X1 MEM_stage_inst_dmem_U4619 ( .A1(MEM_stage_inst_dmem_ram_2520), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n4476) );
NOR2_X1 MEM_stage_inst_dmem_U4618 ( .A1(MEM_stage_inst_dmem_n4474), .A2(MEM_stage_inst_dmem_n4473), .ZN(MEM_stage_inst_dmem_n4482) );
NAND2_X1 MEM_stage_inst_dmem_U4617 ( .A1(MEM_stage_inst_dmem_n4472), .A2(MEM_stage_inst_dmem_n4471), .ZN(MEM_stage_inst_dmem_n4473) );
NAND2_X1 MEM_stage_inst_dmem_U4616 ( .A1(MEM_stage_inst_dmem_ram_2824), .A2(MEM_stage_inst_dmem_n8472), .ZN(MEM_stage_inst_dmem_n4471) );
NAND2_X1 MEM_stage_inst_dmem_U4615 ( .A1(MEM_stage_inst_dmem_ram_2056), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n4472) );
NAND2_X1 MEM_stage_inst_dmem_U4614 ( .A1(MEM_stage_inst_dmem_n4470), .A2(MEM_stage_inst_dmem_n4469), .ZN(MEM_stage_inst_dmem_n4474) );
NAND2_X1 MEM_stage_inst_dmem_U4613 ( .A1(MEM_stage_inst_dmem_ram_2408), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n4469) );
NAND2_X1 MEM_stage_inst_dmem_U4612 ( .A1(MEM_stage_inst_dmem_ram_2392), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n4470) );
NAND2_X1 MEM_stage_inst_dmem_U4611 ( .A1(MEM_stage_inst_dmem_n4468), .A2(MEM_stage_inst_dmem_n4467), .ZN(MEM_stage_inst_dmem_n4484) );
NOR2_X1 MEM_stage_inst_dmem_U4610 ( .A1(MEM_stage_inst_dmem_n4466), .A2(MEM_stage_inst_dmem_n4465), .ZN(MEM_stage_inst_dmem_n4467) );
NAND2_X1 MEM_stage_inst_dmem_U4609 ( .A1(MEM_stage_inst_dmem_n4464), .A2(MEM_stage_inst_dmem_n4463), .ZN(MEM_stage_inst_dmem_n4465) );
NAND2_X1 MEM_stage_inst_dmem_U4608 ( .A1(MEM_stage_inst_dmem_ram_3032), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n4463) );
NAND2_X1 MEM_stage_inst_dmem_U4607 ( .A1(MEM_stage_inst_dmem_ram_2264), .A2(MEM_stage_inst_dmem_n51), .ZN(MEM_stage_inst_dmem_n4464) );
NAND2_X1 MEM_stage_inst_dmem_U4606 ( .A1(MEM_stage_inst_dmem_n4462), .A2(MEM_stage_inst_dmem_n4461), .ZN(MEM_stage_inst_dmem_n4466) );
NAND2_X1 MEM_stage_inst_dmem_U4605 ( .A1(MEM_stage_inst_dmem_ram_3000), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n4461) );
NAND2_X1 MEM_stage_inst_dmem_U4604 ( .A1(MEM_stage_inst_dmem_ram_2136), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n4462) );
NOR2_X1 MEM_stage_inst_dmem_U4603 ( .A1(MEM_stage_inst_dmem_n4460), .A2(MEM_stage_inst_dmem_n4459), .ZN(MEM_stage_inst_dmem_n4468) );
NAND2_X1 MEM_stage_inst_dmem_U4602 ( .A1(MEM_stage_inst_dmem_n4458), .A2(MEM_stage_inst_dmem_n4457), .ZN(MEM_stage_inst_dmem_n4459) );
NAND2_X1 MEM_stage_inst_dmem_U4601 ( .A1(MEM_stage_inst_dmem_ram_2248), .A2(MEM_stage_inst_dmem_n36), .ZN(MEM_stage_inst_dmem_n4457) );
NAND2_X1 MEM_stage_inst_dmem_U4600 ( .A1(MEM_stage_inst_dmem_ram_2456), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n4458) );
NAND2_X1 MEM_stage_inst_dmem_U4599 ( .A1(MEM_stage_inst_dmem_n4456), .A2(MEM_stage_inst_dmem_n4455), .ZN(MEM_stage_inst_dmem_n4460) );
NAND2_X1 MEM_stage_inst_dmem_U4598 ( .A1(MEM_stage_inst_dmem_ram_3048), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n4455) );
NAND2_X1 MEM_stage_inst_dmem_U4597 ( .A1(MEM_stage_inst_dmem_ram_3064), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n4456) );
NAND2_X1 MEM_stage_inst_dmem_U4596 ( .A1(MEM_stage_inst_dmem_n4454), .A2(MEM_stage_inst_dmem_n4453), .ZN(MEM_stage_inst_dmem_n4518) );
NOR2_X1 MEM_stage_inst_dmem_U4595 ( .A1(MEM_stage_inst_dmem_n4452), .A2(MEM_stage_inst_dmem_n4451), .ZN(MEM_stage_inst_dmem_n4453) );
NAND2_X1 MEM_stage_inst_dmem_U4594 ( .A1(MEM_stage_inst_dmem_n4450), .A2(MEM_stage_inst_dmem_n4449), .ZN(MEM_stage_inst_dmem_n4451) );
NOR2_X1 MEM_stage_inst_dmem_U4593 ( .A1(MEM_stage_inst_dmem_n4448), .A2(MEM_stage_inst_dmem_n4447), .ZN(MEM_stage_inst_dmem_n4449) );
NAND2_X1 MEM_stage_inst_dmem_U4592 ( .A1(MEM_stage_inst_dmem_n4446), .A2(MEM_stage_inst_dmem_n4445), .ZN(MEM_stage_inst_dmem_n4447) );
NAND2_X1 MEM_stage_inst_dmem_U4591 ( .A1(MEM_stage_inst_dmem_ram_2920), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n4445) );
NAND2_X1 MEM_stage_inst_dmem_U4590 ( .A1(MEM_stage_inst_dmem_ram_2680), .A2(MEM_stage_inst_dmem_n4652), .ZN(MEM_stage_inst_dmem_n4446) );
NAND2_X1 MEM_stage_inst_dmem_U4589 ( .A1(MEM_stage_inst_dmem_n4444), .A2(MEM_stage_inst_dmem_n4443), .ZN(MEM_stage_inst_dmem_n4448) );
NAND2_X1 MEM_stage_inst_dmem_U4588 ( .A1(MEM_stage_inst_dmem_ram_2360), .A2(MEM_stage_inst_dmem_n4731), .ZN(MEM_stage_inst_dmem_n4443) );
NAND2_X1 MEM_stage_inst_dmem_U4587 ( .A1(MEM_stage_inst_dmem_ram_2808), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n4444) );
NOR2_X1 MEM_stage_inst_dmem_U4586 ( .A1(MEM_stage_inst_dmem_n4442), .A2(MEM_stage_inst_dmem_n4441), .ZN(MEM_stage_inst_dmem_n4450) );
NAND2_X1 MEM_stage_inst_dmem_U4585 ( .A1(MEM_stage_inst_dmem_n4440), .A2(MEM_stage_inst_dmem_n4439), .ZN(MEM_stage_inst_dmem_n4441) );
NAND2_X1 MEM_stage_inst_dmem_U4584 ( .A1(MEM_stage_inst_dmem_ram_2280), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n4439) );
NAND2_X1 MEM_stage_inst_dmem_U4583 ( .A1(MEM_stage_inst_dmem_ram_2984), .A2(MEM_stage_inst_dmem_n4675), .ZN(MEM_stage_inst_dmem_n4440) );
NAND2_X1 MEM_stage_inst_dmem_U4582 ( .A1(MEM_stage_inst_dmem_n4438), .A2(MEM_stage_inst_dmem_n4437), .ZN(MEM_stage_inst_dmem_n4442) );
NAND2_X1 MEM_stage_inst_dmem_U4581 ( .A1(MEM_stage_inst_dmem_ram_2728), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n4437) );
NAND2_X1 MEM_stage_inst_dmem_U4580 ( .A1(MEM_stage_inst_dmem_ram_2344), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n4438) );
NAND2_X1 MEM_stage_inst_dmem_U4579 ( .A1(MEM_stage_inst_dmem_n4436), .A2(MEM_stage_inst_dmem_n4435), .ZN(MEM_stage_inst_dmem_n4452) );
NOR2_X1 MEM_stage_inst_dmem_U4578 ( .A1(MEM_stage_inst_dmem_n4434), .A2(MEM_stage_inst_dmem_n4433), .ZN(MEM_stage_inst_dmem_n4435) );
NAND2_X1 MEM_stage_inst_dmem_U4577 ( .A1(MEM_stage_inst_dmem_n4432), .A2(MEM_stage_inst_dmem_n4431), .ZN(MEM_stage_inst_dmem_n4433) );
NAND2_X1 MEM_stage_inst_dmem_U4576 ( .A1(MEM_stage_inst_dmem_ram_2472), .A2(MEM_stage_inst_dmem_n4772), .ZN(MEM_stage_inst_dmem_n4431) );
NAND2_X1 MEM_stage_inst_dmem_U4575 ( .A1(MEM_stage_inst_dmem_ram_2600), .A2(MEM_stage_inst_dmem_n4692), .ZN(MEM_stage_inst_dmem_n4432) );
NAND2_X1 MEM_stage_inst_dmem_U4574 ( .A1(MEM_stage_inst_dmem_n4430), .A2(MEM_stage_inst_dmem_n4429), .ZN(MEM_stage_inst_dmem_n4434) );
NAND2_X1 MEM_stage_inst_dmem_U4573 ( .A1(MEM_stage_inst_dmem_ram_3016), .A2(MEM_stage_inst_dmem_n4728), .ZN(MEM_stage_inst_dmem_n4429) );
NAND2_X1 MEM_stage_inst_dmem_U4572 ( .A1(MEM_stage_inst_dmem_ram_2856), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n4430) );
NOR2_X1 MEM_stage_inst_dmem_U4571 ( .A1(MEM_stage_inst_dmem_n4428), .A2(MEM_stage_inst_dmem_n4427), .ZN(MEM_stage_inst_dmem_n4436) );
NAND2_X1 MEM_stage_inst_dmem_U4570 ( .A1(MEM_stage_inst_dmem_n4426), .A2(MEM_stage_inst_dmem_n4425), .ZN(MEM_stage_inst_dmem_n4427) );
NAND2_X1 MEM_stage_inst_dmem_U4569 ( .A1(MEM_stage_inst_dmem_ram_2232), .A2(MEM_stage_inst_dmem_n8434), .ZN(MEM_stage_inst_dmem_n4425) );
NAND2_X1 MEM_stage_inst_dmem_U4568 ( .A1(MEM_stage_inst_dmem_ram_2584), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n4426) );
NAND2_X1 MEM_stage_inst_dmem_U4567 ( .A1(MEM_stage_inst_dmem_n4424), .A2(MEM_stage_inst_dmem_n4423), .ZN(MEM_stage_inst_dmem_n4428) );
NAND2_X1 MEM_stage_inst_dmem_U4566 ( .A1(MEM_stage_inst_dmem_ram_2696), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n4423) );
NAND2_X1 MEM_stage_inst_dmem_U4565 ( .A1(MEM_stage_inst_dmem_ram_2744), .A2(MEM_stage_inst_dmem_n4709), .ZN(MEM_stage_inst_dmem_n4424) );
NOR2_X1 MEM_stage_inst_dmem_U4564 ( .A1(MEM_stage_inst_dmem_n4422), .A2(MEM_stage_inst_dmem_n4421), .ZN(MEM_stage_inst_dmem_n4454) );
NAND2_X1 MEM_stage_inst_dmem_U4563 ( .A1(MEM_stage_inst_dmem_n4420), .A2(MEM_stage_inst_dmem_n4419), .ZN(MEM_stage_inst_dmem_n4421) );
NOR2_X1 MEM_stage_inst_dmem_U4562 ( .A1(MEM_stage_inst_dmem_n4418), .A2(MEM_stage_inst_dmem_n4417), .ZN(MEM_stage_inst_dmem_n4419) );
NAND2_X1 MEM_stage_inst_dmem_U4561 ( .A1(MEM_stage_inst_dmem_n4416), .A2(MEM_stage_inst_dmem_n4415), .ZN(MEM_stage_inst_dmem_n4417) );
NAND2_X1 MEM_stage_inst_dmem_U4560 ( .A1(MEM_stage_inst_dmem_ram_2840), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n4415) );
NAND2_X1 MEM_stage_inst_dmem_U4559 ( .A1(MEM_stage_inst_dmem_ram_2776), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n4416) );
NAND2_X1 MEM_stage_inst_dmem_U4558 ( .A1(MEM_stage_inst_dmem_n4414), .A2(MEM_stage_inst_dmem_n4413), .ZN(MEM_stage_inst_dmem_n4418) );
NAND2_X1 MEM_stage_inst_dmem_U4557 ( .A1(MEM_stage_inst_dmem_ram_2184), .A2(MEM_stage_inst_dmem_n61), .ZN(MEM_stage_inst_dmem_n4413) );
NAND2_X1 MEM_stage_inst_dmem_U4556 ( .A1(MEM_stage_inst_dmem_ram_2504), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n4414) );
NOR2_X1 MEM_stage_inst_dmem_U4555 ( .A1(MEM_stage_inst_dmem_n4412), .A2(MEM_stage_inst_dmem_n4411), .ZN(MEM_stage_inst_dmem_n4420) );
NAND2_X1 MEM_stage_inst_dmem_U4554 ( .A1(MEM_stage_inst_dmem_n4410), .A2(MEM_stage_inst_dmem_n4409), .ZN(MEM_stage_inst_dmem_n4411) );
NAND2_X1 MEM_stage_inst_dmem_U4553 ( .A1(MEM_stage_inst_dmem_ram_2936), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n4409) );
NAND2_X1 MEM_stage_inst_dmem_U4552 ( .A1(MEM_stage_inst_dmem_ram_2904), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n4410) );
NAND2_X1 MEM_stage_inst_dmem_U4551 ( .A1(MEM_stage_inst_dmem_n4408), .A2(MEM_stage_inst_dmem_n4407), .ZN(MEM_stage_inst_dmem_n4412) );
NAND2_X1 MEM_stage_inst_dmem_U4550 ( .A1(MEM_stage_inst_dmem_ram_2552), .A2(MEM_stage_inst_dmem_n64), .ZN(MEM_stage_inst_dmem_n4407) );
NAND2_X1 MEM_stage_inst_dmem_U4549 ( .A1(MEM_stage_inst_dmem_ram_2888), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n4408) );
NAND2_X1 MEM_stage_inst_dmem_U4548 ( .A1(MEM_stage_inst_dmem_n4406), .A2(MEM_stage_inst_dmem_n4405), .ZN(MEM_stage_inst_dmem_n4422) );
NOR2_X1 MEM_stage_inst_dmem_U4547 ( .A1(MEM_stage_inst_dmem_n4404), .A2(MEM_stage_inst_dmem_n4403), .ZN(MEM_stage_inst_dmem_n4405) );
NAND2_X1 MEM_stage_inst_dmem_U4546 ( .A1(MEM_stage_inst_dmem_n4402), .A2(MEM_stage_inst_dmem_n4401), .ZN(MEM_stage_inst_dmem_n4403) );
NAND2_X1 MEM_stage_inst_dmem_U4545 ( .A1(MEM_stage_inst_dmem_ram_2152), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n4401) );
NAND2_X1 MEM_stage_inst_dmem_U4544 ( .A1(MEM_stage_inst_dmem_ram_2632), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n4402) );
NAND2_X1 MEM_stage_inst_dmem_U4543 ( .A1(MEM_stage_inst_dmem_n4400), .A2(MEM_stage_inst_dmem_n4399), .ZN(MEM_stage_inst_dmem_n4404) );
NAND2_X1 MEM_stage_inst_dmem_U4542 ( .A1(MEM_stage_inst_dmem_ram_2376), .A2(MEM_stage_inst_dmem_n4706), .ZN(MEM_stage_inst_dmem_n4399) );
NAND2_X1 MEM_stage_inst_dmem_U4541 ( .A1(MEM_stage_inst_dmem_ram_2328), .A2(MEM_stage_inst_dmem_n4672), .ZN(MEM_stage_inst_dmem_n4400) );
NOR2_X1 MEM_stage_inst_dmem_U4540 ( .A1(MEM_stage_inst_dmem_n4398), .A2(MEM_stage_inst_dmem_n4397), .ZN(MEM_stage_inst_dmem_n4406) );
NAND2_X1 MEM_stage_inst_dmem_U4539 ( .A1(MEM_stage_inst_dmem_n4396), .A2(MEM_stage_inst_dmem_n4395), .ZN(MEM_stage_inst_dmem_n4397) );
NAND2_X1 MEM_stage_inst_dmem_U4538 ( .A1(MEM_stage_inst_dmem_ram_2536), .A2(MEM_stage_inst_dmem_n4667), .ZN(MEM_stage_inst_dmem_n4395) );
NAND2_X1 MEM_stage_inst_dmem_U4537 ( .A1(MEM_stage_inst_dmem_ram_2968), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n4396) );
NAND2_X1 MEM_stage_inst_dmem_U4536 ( .A1(MEM_stage_inst_dmem_n4394), .A2(MEM_stage_inst_dmem_n4393), .ZN(MEM_stage_inst_dmem_n4398) );
NAND2_X1 MEM_stage_inst_dmem_U4535 ( .A1(MEM_stage_inst_dmem_ram_2488), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n4393) );
NAND2_X1 MEM_stage_inst_dmem_U4534 ( .A1(MEM_stage_inst_dmem_ram_2312), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n4394) );
NAND2_X1 MEM_stage_inst_dmem_U4533 ( .A1(MEM_stage_inst_dmem_n4392), .A2(MEM_stage_inst_dmem_n4391), .ZN(MEM_stage_inst_mem_read_data_7) );
NOR2_X1 MEM_stage_inst_dmem_U4532 ( .A1(MEM_stage_inst_dmem_n4390), .A2(MEM_stage_inst_dmem_n4389), .ZN(MEM_stage_inst_dmem_n4391) );
NOR2_X1 MEM_stage_inst_dmem_U4531 ( .A1(MEM_stage_inst_dmem_n4388), .A2(MEM_stage_inst_dmem_n8152), .ZN(MEM_stage_inst_dmem_n4389) );
NOR2_X1 MEM_stage_inst_dmem_U4530 ( .A1(MEM_stage_inst_dmem_n4387), .A2(MEM_stage_inst_dmem_n4386), .ZN(MEM_stage_inst_dmem_n4388) );
NAND2_X1 MEM_stage_inst_dmem_U4529 ( .A1(MEM_stage_inst_dmem_n4385), .A2(MEM_stage_inst_dmem_n4384), .ZN(MEM_stage_inst_dmem_n4386) );
NOR2_X1 MEM_stage_inst_dmem_U4528 ( .A1(MEM_stage_inst_dmem_n4383), .A2(MEM_stage_inst_dmem_n4382), .ZN(MEM_stage_inst_dmem_n4384) );
NAND2_X1 MEM_stage_inst_dmem_U4527 ( .A1(MEM_stage_inst_dmem_n4381), .A2(MEM_stage_inst_dmem_n4380), .ZN(MEM_stage_inst_dmem_n4382) );
NOR2_X1 MEM_stage_inst_dmem_U4526 ( .A1(MEM_stage_inst_dmem_n4379), .A2(MEM_stage_inst_dmem_n4378), .ZN(MEM_stage_inst_dmem_n4380) );
NAND2_X1 MEM_stage_inst_dmem_U4525 ( .A1(MEM_stage_inst_dmem_n4377), .A2(MEM_stage_inst_dmem_n4376), .ZN(MEM_stage_inst_dmem_n4378) );
NAND2_X1 MEM_stage_inst_dmem_U4524 ( .A1(MEM_stage_inst_dmem_ram_1511), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n4376) );
NAND2_X1 MEM_stage_inst_dmem_U4523 ( .A1(MEM_stage_inst_dmem_ram_1655), .A2(MEM_stage_inst_dmem_n4652), .ZN(MEM_stage_inst_dmem_n4377) );
NAND2_X1 MEM_stage_inst_dmem_U4522 ( .A1(MEM_stage_inst_dmem_n4375), .A2(MEM_stage_inst_dmem_n4374), .ZN(MEM_stage_inst_dmem_n4379) );
NAND2_X1 MEM_stage_inst_dmem_U4521 ( .A1(MEM_stage_inst_dmem_ram_1863), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n4374) );
NAND2_X1 MEM_stage_inst_dmem_U4520 ( .A1(MEM_stage_inst_dmem_ram_1175), .A2(MEM_stage_inst_dmem_n5807), .ZN(MEM_stage_inst_dmem_n4375) );
NOR2_X1 MEM_stage_inst_dmem_U4519 ( .A1(MEM_stage_inst_dmem_n4373), .A2(MEM_stage_inst_dmem_n4372), .ZN(MEM_stage_inst_dmem_n4381) );
NAND2_X1 MEM_stage_inst_dmem_U4518 ( .A1(MEM_stage_inst_dmem_n4371), .A2(MEM_stage_inst_dmem_n4370), .ZN(MEM_stage_inst_dmem_n4372) );
NAND2_X1 MEM_stage_inst_dmem_U4517 ( .A1(MEM_stage_inst_dmem_ram_1799), .A2(MEM_stage_inst_dmem_n37), .ZN(MEM_stage_inst_dmem_n4370) );
NAND2_X1 MEM_stage_inst_dmem_U4516 ( .A1(MEM_stage_inst_dmem_ram_2023), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n4371) );
NAND2_X1 MEM_stage_inst_dmem_U4515 ( .A1(MEM_stage_inst_dmem_n4369), .A2(MEM_stage_inst_dmem_n4368), .ZN(MEM_stage_inst_dmem_n4373) );
NAND2_X1 MEM_stage_inst_dmem_U4514 ( .A1(MEM_stage_inst_dmem_ram_1079), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n4368) );
NAND2_X1 MEM_stage_inst_dmem_U4513 ( .A1(MEM_stage_inst_dmem_ram_1783), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n4369) );
NAND2_X1 MEM_stage_inst_dmem_U4512 ( .A1(MEM_stage_inst_dmem_n4367), .A2(MEM_stage_inst_dmem_n4366), .ZN(MEM_stage_inst_dmem_n4383) );
NOR2_X1 MEM_stage_inst_dmem_U4511 ( .A1(MEM_stage_inst_dmem_n4365), .A2(MEM_stage_inst_dmem_n4364), .ZN(MEM_stage_inst_dmem_n4366) );
NAND2_X1 MEM_stage_inst_dmem_U4510 ( .A1(MEM_stage_inst_dmem_n4363), .A2(MEM_stage_inst_dmem_n4362), .ZN(MEM_stage_inst_dmem_n4364) );
NAND2_X1 MEM_stage_inst_dmem_U4509 ( .A1(MEM_stage_inst_dmem_ram_1575), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n4362) );
NAND2_X1 MEM_stage_inst_dmem_U4508 ( .A1(MEM_stage_inst_dmem_ram_1559), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n4363) );
NAND2_X1 MEM_stage_inst_dmem_U4507 ( .A1(MEM_stage_inst_dmem_n4361), .A2(MEM_stage_inst_dmem_n4360), .ZN(MEM_stage_inst_dmem_n4365) );
NAND2_X1 MEM_stage_inst_dmem_U4506 ( .A1(MEM_stage_inst_dmem_ram_2007), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n4360) );
NAND2_X1 MEM_stage_inst_dmem_U4505 ( .A1(MEM_stage_inst_dmem_ram_1719), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n4361) );
NOR2_X1 MEM_stage_inst_dmem_U4504 ( .A1(MEM_stage_inst_dmem_n4359), .A2(MEM_stage_inst_dmem_n4358), .ZN(MEM_stage_inst_dmem_n4367) );
NAND2_X1 MEM_stage_inst_dmem_U4503 ( .A1(MEM_stage_inst_dmem_n4357), .A2(MEM_stage_inst_dmem_n4356), .ZN(MEM_stage_inst_dmem_n4358) );
NAND2_X1 MEM_stage_inst_dmem_U4502 ( .A1(MEM_stage_inst_dmem_ram_1831), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n4356) );
NAND2_X1 MEM_stage_inst_dmem_U4501 ( .A1(MEM_stage_inst_dmem_ram_1687), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n4357) );
NAND2_X1 MEM_stage_inst_dmem_U4500 ( .A1(MEM_stage_inst_dmem_n4355), .A2(MEM_stage_inst_dmem_n4354), .ZN(MEM_stage_inst_dmem_n4359) );
NAND2_X1 MEM_stage_inst_dmem_U4499 ( .A1(MEM_stage_inst_dmem_ram_1527), .A2(MEM_stage_inst_dmem_n64), .ZN(MEM_stage_inst_dmem_n4354) );
NAND2_X1 MEM_stage_inst_dmem_U4498 ( .A1(MEM_stage_inst_dmem_ram_2039), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n4355) );
NOR2_X1 MEM_stage_inst_dmem_U4497 ( .A1(MEM_stage_inst_dmem_n4353), .A2(MEM_stage_inst_dmem_n4352), .ZN(MEM_stage_inst_dmem_n4385) );
NAND2_X1 MEM_stage_inst_dmem_U4496 ( .A1(MEM_stage_inst_dmem_n4351), .A2(MEM_stage_inst_dmem_n4350), .ZN(MEM_stage_inst_dmem_n4352) );
NOR2_X1 MEM_stage_inst_dmem_U4495 ( .A1(MEM_stage_inst_dmem_n4349), .A2(MEM_stage_inst_dmem_n4348), .ZN(MEM_stage_inst_dmem_n4350) );
NAND2_X1 MEM_stage_inst_dmem_U4494 ( .A1(MEM_stage_inst_dmem_n4347), .A2(MEM_stage_inst_dmem_n4346), .ZN(MEM_stage_inst_dmem_n4348) );
NAND2_X1 MEM_stage_inst_dmem_U4493 ( .A1(MEM_stage_inst_dmem_ram_1927), .A2(MEM_stage_inst_dmem_n72), .ZN(MEM_stage_inst_dmem_n4346) );
NAND2_X1 MEM_stage_inst_dmem_U4492 ( .A1(MEM_stage_inst_dmem_ram_1815), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n4347) );
NAND2_X1 MEM_stage_inst_dmem_U4491 ( .A1(MEM_stage_inst_dmem_n4345), .A2(MEM_stage_inst_dmem_n4344), .ZN(MEM_stage_inst_dmem_n4349) );
NAND2_X1 MEM_stage_inst_dmem_U4490 ( .A1(MEM_stage_inst_dmem_ram_1351), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n4344) );
NAND2_X1 MEM_stage_inst_dmem_U4489 ( .A1(MEM_stage_inst_dmem_ram_1063), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n4345) );
NOR2_X1 MEM_stage_inst_dmem_U4488 ( .A1(MEM_stage_inst_dmem_n4343), .A2(MEM_stage_inst_dmem_n4342), .ZN(MEM_stage_inst_dmem_n4351) );
NAND2_X1 MEM_stage_inst_dmem_U4487 ( .A1(MEM_stage_inst_dmem_n4341), .A2(MEM_stage_inst_dmem_n4340), .ZN(MEM_stage_inst_dmem_n4342) );
NAND2_X1 MEM_stage_inst_dmem_U4486 ( .A1(MEM_stage_inst_dmem_ram_1991), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n4340) );
NAND2_X1 MEM_stage_inst_dmem_U4485 ( .A1(MEM_stage_inst_dmem_ram_1271), .A2(MEM_stage_inst_dmem_n39), .ZN(MEM_stage_inst_dmem_n4341) );
NAND2_X1 MEM_stage_inst_dmem_U4484 ( .A1(MEM_stage_inst_dmem_n4339), .A2(MEM_stage_inst_dmem_n4338), .ZN(MEM_stage_inst_dmem_n4343) );
NAND2_X1 MEM_stage_inst_dmem_U4483 ( .A1(MEM_stage_inst_dmem_ram_1207), .A2(MEM_stage_inst_dmem_n55), .ZN(MEM_stage_inst_dmem_n4338) );
NAND2_X1 MEM_stage_inst_dmem_U4482 ( .A1(MEM_stage_inst_dmem_ram_1607), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n4339) );
NAND2_X1 MEM_stage_inst_dmem_U4481 ( .A1(MEM_stage_inst_dmem_n4337), .A2(MEM_stage_inst_dmem_n4336), .ZN(MEM_stage_inst_dmem_n4353) );
NOR2_X1 MEM_stage_inst_dmem_U4480 ( .A1(MEM_stage_inst_dmem_n4335), .A2(MEM_stage_inst_dmem_n4334), .ZN(MEM_stage_inst_dmem_n4336) );
NAND2_X1 MEM_stage_inst_dmem_U4479 ( .A1(MEM_stage_inst_dmem_n4333), .A2(MEM_stage_inst_dmem_n4332), .ZN(MEM_stage_inst_dmem_n4334) );
NAND2_X1 MEM_stage_inst_dmem_U4478 ( .A1(MEM_stage_inst_dmem_ram_1735), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n4332) );
NAND2_X1 MEM_stage_inst_dmem_U4477 ( .A1(MEM_stage_inst_dmem_ram_1767), .A2(MEM_stage_inst_dmem_n4769), .ZN(MEM_stage_inst_dmem_n4333) );
NAND2_X1 MEM_stage_inst_dmem_U4476 ( .A1(MEM_stage_inst_dmem_n4331), .A2(MEM_stage_inst_dmem_n4330), .ZN(MEM_stage_inst_dmem_n4335) );
NAND2_X1 MEM_stage_inst_dmem_U4475 ( .A1(MEM_stage_inst_dmem_ram_1447), .A2(MEM_stage_inst_dmem_n4772), .ZN(MEM_stage_inst_dmem_n4330) );
NAND2_X1 MEM_stage_inst_dmem_U4474 ( .A1(MEM_stage_inst_dmem_ram_1623), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n4331) );
NOR2_X1 MEM_stage_inst_dmem_U4473 ( .A1(MEM_stage_inst_dmem_n4329), .A2(MEM_stage_inst_dmem_n4328), .ZN(MEM_stage_inst_dmem_n4337) );
NAND2_X1 MEM_stage_inst_dmem_U4472 ( .A1(MEM_stage_inst_dmem_n4327), .A2(MEM_stage_inst_dmem_n4326), .ZN(MEM_stage_inst_dmem_n4328) );
NAND2_X1 MEM_stage_inst_dmem_U4471 ( .A1(MEM_stage_inst_dmem_ram_1703), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n4326) );
NAND2_X1 MEM_stage_inst_dmem_U4470 ( .A1(MEM_stage_inst_dmem_ram_1479), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n4327) );
NAND2_X1 MEM_stage_inst_dmem_U4469 ( .A1(MEM_stage_inst_dmem_n4325), .A2(MEM_stage_inst_dmem_n4324), .ZN(MEM_stage_inst_dmem_n4329) );
NAND2_X1 MEM_stage_inst_dmem_U4468 ( .A1(MEM_stage_inst_dmem_ram_1383), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n4324) );
NAND2_X1 MEM_stage_inst_dmem_U4467 ( .A1(MEM_stage_inst_dmem_ram_1191), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n4325) );
NAND2_X1 MEM_stage_inst_dmem_U4466 ( .A1(MEM_stage_inst_dmem_n4323), .A2(MEM_stage_inst_dmem_n4322), .ZN(MEM_stage_inst_dmem_n4387) );
NOR2_X1 MEM_stage_inst_dmem_U4465 ( .A1(MEM_stage_inst_dmem_n4321), .A2(MEM_stage_inst_dmem_n4320), .ZN(MEM_stage_inst_dmem_n4322) );
NAND2_X1 MEM_stage_inst_dmem_U4464 ( .A1(MEM_stage_inst_dmem_n4319), .A2(MEM_stage_inst_dmem_n4318), .ZN(MEM_stage_inst_dmem_n4320) );
NOR2_X1 MEM_stage_inst_dmem_U4463 ( .A1(MEM_stage_inst_dmem_n4317), .A2(MEM_stage_inst_dmem_n4316), .ZN(MEM_stage_inst_dmem_n4318) );
NAND2_X1 MEM_stage_inst_dmem_U4462 ( .A1(MEM_stage_inst_dmem_n4315), .A2(MEM_stage_inst_dmem_n4314), .ZN(MEM_stage_inst_dmem_n4316) );
NAND2_X1 MEM_stage_inst_dmem_U4461 ( .A1(MEM_stage_inst_dmem_ram_1671), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n4314) );
NAND2_X1 MEM_stage_inst_dmem_U4460 ( .A1(MEM_stage_inst_dmem_ram_1639), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n4315) );
NAND2_X1 MEM_stage_inst_dmem_U4459 ( .A1(MEM_stage_inst_dmem_n4313), .A2(MEM_stage_inst_dmem_n4312), .ZN(MEM_stage_inst_dmem_n4317) );
NAND2_X1 MEM_stage_inst_dmem_U4458 ( .A1(MEM_stage_inst_dmem_ram_1095), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n4312) );
NAND2_X1 MEM_stage_inst_dmem_U4457 ( .A1(MEM_stage_inst_dmem_ram_1111), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n4313) );
NOR2_X1 MEM_stage_inst_dmem_U4456 ( .A1(MEM_stage_inst_dmem_n4311), .A2(MEM_stage_inst_dmem_n4310), .ZN(MEM_stage_inst_dmem_n4319) );
NAND2_X1 MEM_stage_inst_dmem_U4455 ( .A1(MEM_stage_inst_dmem_n4309), .A2(MEM_stage_inst_dmem_n4308), .ZN(MEM_stage_inst_dmem_n4310) );
NAND2_X1 MEM_stage_inst_dmem_U4454 ( .A1(MEM_stage_inst_dmem_ram_1223), .A2(MEM_stage_inst_dmem_n36), .ZN(MEM_stage_inst_dmem_n4308) );
NAND2_X1 MEM_stage_inst_dmem_U4453 ( .A1(MEM_stage_inst_dmem_ram_1159), .A2(MEM_stage_inst_dmem_n61), .ZN(MEM_stage_inst_dmem_n4309) );
NAND2_X1 MEM_stage_inst_dmem_U4452 ( .A1(MEM_stage_inst_dmem_n4307), .A2(MEM_stage_inst_dmem_n4306), .ZN(MEM_stage_inst_dmem_n4311) );
NAND2_X1 MEM_stage_inst_dmem_U4451 ( .A1(MEM_stage_inst_dmem_ram_1335), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n4306) );
NAND2_X1 MEM_stage_inst_dmem_U4450 ( .A1(MEM_stage_inst_dmem_ram_1543), .A2(MEM_stage_inst_dmem_n71), .ZN(MEM_stage_inst_dmem_n4307) );
NAND2_X1 MEM_stage_inst_dmem_U4449 ( .A1(MEM_stage_inst_dmem_n4305), .A2(MEM_stage_inst_dmem_n4304), .ZN(MEM_stage_inst_dmem_n4321) );
NOR2_X1 MEM_stage_inst_dmem_U4448 ( .A1(MEM_stage_inst_dmem_n4303), .A2(MEM_stage_inst_dmem_n4302), .ZN(MEM_stage_inst_dmem_n4304) );
NAND2_X1 MEM_stage_inst_dmem_U4447 ( .A1(MEM_stage_inst_dmem_n4301), .A2(MEM_stage_inst_dmem_n4300), .ZN(MEM_stage_inst_dmem_n4302) );
NAND2_X1 MEM_stage_inst_dmem_U4446 ( .A1(MEM_stage_inst_dmem_ram_1911), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n4300) );
NAND2_X1 MEM_stage_inst_dmem_U4445 ( .A1(MEM_stage_inst_dmem_ram_1143), .A2(MEM_stage_inst_dmem_n4710), .ZN(MEM_stage_inst_dmem_n4301) );
NAND2_X1 MEM_stage_inst_dmem_U4444 ( .A1(MEM_stage_inst_dmem_n4299), .A2(MEM_stage_inst_dmem_n4298), .ZN(MEM_stage_inst_dmem_n4303) );
NAND2_X1 MEM_stage_inst_dmem_U4443 ( .A1(MEM_stage_inst_dmem_ram_1031), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n4298) );
NAND2_X1 MEM_stage_inst_dmem_U4442 ( .A1(MEM_stage_inst_dmem_ram_1287), .A2(MEM_stage_inst_dmem_n7898), .ZN(MEM_stage_inst_dmem_n4299) );
NOR2_X1 MEM_stage_inst_dmem_U4441 ( .A1(MEM_stage_inst_dmem_n4297), .A2(MEM_stage_inst_dmem_n4296), .ZN(MEM_stage_inst_dmem_n4305) );
NAND2_X1 MEM_stage_inst_dmem_U4440 ( .A1(MEM_stage_inst_dmem_n4295), .A2(MEM_stage_inst_dmem_n4294), .ZN(MEM_stage_inst_dmem_n4296) );
NAND2_X1 MEM_stage_inst_dmem_U4439 ( .A1(MEM_stage_inst_dmem_ram_1895), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n4294) );
NAND2_X1 MEM_stage_inst_dmem_U4438 ( .A1(MEM_stage_inst_dmem_ram_1943), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n4295) );
NAND2_X1 MEM_stage_inst_dmem_U4437 ( .A1(MEM_stage_inst_dmem_n4293), .A2(MEM_stage_inst_dmem_n4292), .ZN(MEM_stage_inst_dmem_n4297) );
NAND2_X1 MEM_stage_inst_dmem_U4436 ( .A1(MEM_stage_inst_dmem_ram_1239), .A2(MEM_stage_inst_dmem_n51), .ZN(MEM_stage_inst_dmem_n4292) );
NAND2_X1 MEM_stage_inst_dmem_U4435 ( .A1(MEM_stage_inst_dmem_ram_1127), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n4293) );
NOR2_X1 MEM_stage_inst_dmem_U4434 ( .A1(MEM_stage_inst_dmem_n4291), .A2(MEM_stage_inst_dmem_n4290), .ZN(MEM_stage_inst_dmem_n4323) );
NAND2_X1 MEM_stage_inst_dmem_U4433 ( .A1(MEM_stage_inst_dmem_n4289), .A2(MEM_stage_inst_dmem_n4288), .ZN(MEM_stage_inst_dmem_n4290) );
NOR2_X1 MEM_stage_inst_dmem_U4432 ( .A1(MEM_stage_inst_dmem_n4287), .A2(MEM_stage_inst_dmem_n4286), .ZN(MEM_stage_inst_dmem_n4288) );
NAND2_X1 MEM_stage_inst_dmem_U4431 ( .A1(MEM_stage_inst_dmem_n4285), .A2(MEM_stage_inst_dmem_n4284), .ZN(MEM_stage_inst_dmem_n4286) );
NAND2_X1 MEM_stage_inst_dmem_U4430 ( .A1(MEM_stage_inst_dmem_ram_1959), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n4284) );
NAND2_X1 MEM_stage_inst_dmem_U4429 ( .A1(MEM_stage_inst_dmem_ram_1319), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n4285) );
NAND2_X1 MEM_stage_inst_dmem_U4428 ( .A1(MEM_stage_inst_dmem_n4283), .A2(MEM_stage_inst_dmem_n4282), .ZN(MEM_stage_inst_dmem_n4287) );
NAND2_X1 MEM_stage_inst_dmem_U4427 ( .A1(MEM_stage_inst_dmem_ram_1255), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n4282) );
NAND2_X1 MEM_stage_inst_dmem_U4426 ( .A1(MEM_stage_inst_dmem_ram_1431), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n4283) );
NOR2_X1 MEM_stage_inst_dmem_U4425 ( .A1(MEM_stage_inst_dmem_n4281), .A2(MEM_stage_inst_dmem_n4280), .ZN(MEM_stage_inst_dmem_n4289) );
NAND2_X1 MEM_stage_inst_dmem_U4424 ( .A1(MEM_stage_inst_dmem_n4279), .A2(MEM_stage_inst_dmem_n4278), .ZN(MEM_stage_inst_dmem_n4280) );
NAND2_X1 MEM_stage_inst_dmem_U4423 ( .A1(MEM_stage_inst_dmem_ram_1975), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n4278) );
NAND2_X1 MEM_stage_inst_dmem_U4422 ( .A1(MEM_stage_inst_dmem_ram_1303), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n4279) );
NAND2_X1 MEM_stage_inst_dmem_U4421 ( .A1(MEM_stage_inst_dmem_n4277), .A2(MEM_stage_inst_dmem_n4276), .ZN(MEM_stage_inst_dmem_n4281) );
NAND2_X1 MEM_stage_inst_dmem_U4420 ( .A1(MEM_stage_inst_dmem_ram_1879), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n4276) );
NAND2_X1 MEM_stage_inst_dmem_U4419 ( .A1(MEM_stage_inst_dmem_ram_1399), .A2(MEM_stage_inst_dmem_n4721), .ZN(MEM_stage_inst_dmem_n4277) );
NAND2_X1 MEM_stage_inst_dmem_U4418 ( .A1(MEM_stage_inst_dmem_n4275), .A2(MEM_stage_inst_dmem_n4274), .ZN(MEM_stage_inst_dmem_n4291) );
NOR2_X1 MEM_stage_inst_dmem_U4417 ( .A1(MEM_stage_inst_dmem_n4273), .A2(MEM_stage_inst_dmem_n4272), .ZN(MEM_stage_inst_dmem_n4274) );
NAND2_X1 MEM_stage_inst_dmem_U4416 ( .A1(MEM_stage_inst_dmem_n4271), .A2(MEM_stage_inst_dmem_n4270), .ZN(MEM_stage_inst_dmem_n4272) );
NAND2_X1 MEM_stage_inst_dmem_U4415 ( .A1(MEM_stage_inst_dmem_ram_1495), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n4270) );
NAND2_X1 MEM_stage_inst_dmem_U4414 ( .A1(MEM_stage_inst_dmem_ram_1415), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n4271) );
NAND2_X1 MEM_stage_inst_dmem_U4413 ( .A1(MEM_stage_inst_dmem_n4269), .A2(MEM_stage_inst_dmem_n4268), .ZN(MEM_stage_inst_dmem_n4273) );
NAND2_X1 MEM_stage_inst_dmem_U4412 ( .A1(MEM_stage_inst_dmem_ram_1847), .A2(MEM_stage_inst_dmem_n46), .ZN(MEM_stage_inst_dmem_n4268) );
NAND2_X1 MEM_stage_inst_dmem_U4411 ( .A1(MEM_stage_inst_dmem_ram_1751), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n4269) );
NOR2_X1 MEM_stage_inst_dmem_U4410 ( .A1(MEM_stage_inst_dmem_n4267), .A2(MEM_stage_inst_dmem_n4266), .ZN(MEM_stage_inst_dmem_n4275) );
NAND2_X1 MEM_stage_inst_dmem_U4409 ( .A1(MEM_stage_inst_dmem_n4265), .A2(MEM_stage_inst_dmem_n4264), .ZN(MEM_stage_inst_dmem_n4266) );
NAND2_X1 MEM_stage_inst_dmem_U4408 ( .A1(MEM_stage_inst_dmem_ram_1591), .A2(MEM_stage_inst_dmem_n41), .ZN(MEM_stage_inst_dmem_n4264) );
NAND2_X1 MEM_stage_inst_dmem_U4407 ( .A1(MEM_stage_inst_dmem_ram_1047), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n4265) );
NAND2_X1 MEM_stage_inst_dmem_U4406 ( .A1(MEM_stage_inst_dmem_n4263), .A2(MEM_stage_inst_dmem_n4262), .ZN(MEM_stage_inst_dmem_n4267) );
NAND2_X1 MEM_stage_inst_dmem_U4405 ( .A1(MEM_stage_inst_dmem_ram_1463), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n4262) );
NAND2_X1 MEM_stage_inst_dmem_U4404 ( .A1(MEM_stage_inst_dmem_ram_1367), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n4263) );
NOR2_X1 MEM_stage_inst_dmem_U4403 ( .A1(MEM_stage_inst_dmem_n4261), .A2(MEM_stage_inst_dmem_n8551), .ZN(MEM_stage_inst_dmem_n4390) );
NOR2_X1 MEM_stage_inst_dmem_U4402 ( .A1(MEM_stage_inst_dmem_n4260), .A2(MEM_stage_inst_dmem_n4259), .ZN(MEM_stage_inst_dmem_n4261) );
NAND2_X1 MEM_stage_inst_dmem_U4401 ( .A1(MEM_stage_inst_dmem_n4258), .A2(MEM_stage_inst_dmem_n4257), .ZN(MEM_stage_inst_dmem_n4259) );
NOR2_X1 MEM_stage_inst_dmem_U4400 ( .A1(MEM_stage_inst_dmem_n4256), .A2(MEM_stage_inst_dmem_n4255), .ZN(MEM_stage_inst_dmem_n4257) );
NAND2_X1 MEM_stage_inst_dmem_U4399 ( .A1(MEM_stage_inst_dmem_n4254), .A2(MEM_stage_inst_dmem_n4253), .ZN(MEM_stage_inst_dmem_n4255) );
NOR2_X1 MEM_stage_inst_dmem_U4398 ( .A1(MEM_stage_inst_dmem_n4252), .A2(MEM_stage_inst_dmem_n4251), .ZN(MEM_stage_inst_dmem_n4253) );
NAND2_X1 MEM_stage_inst_dmem_U4397 ( .A1(MEM_stage_inst_dmem_n4250), .A2(MEM_stage_inst_dmem_n4249), .ZN(MEM_stage_inst_dmem_n4251) );
NAND2_X1 MEM_stage_inst_dmem_U4396 ( .A1(MEM_stage_inst_dmem_ram_695), .A2(MEM_stage_inst_dmem_n4709), .ZN(MEM_stage_inst_dmem_n4249) );
NAND2_X1 MEM_stage_inst_dmem_U4395 ( .A1(MEM_stage_inst_dmem_ram_583), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n4250) );
NAND2_X1 MEM_stage_inst_dmem_U4394 ( .A1(MEM_stage_inst_dmem_n4248), .A2(MEM_stage_inst_dmem_n4247), .ZN(MEM_stage_inst_dmem_n4252) );
NAND2_X1 MEM_stage_inst_dmem_U4393 ( .A1(MEM_stage_inst_dmem_ram_231), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n4247) );
NAND2_X1 MEM_stage_inst_dmem_U4392 ( .A1(MEM_stage_inst_dmem_ram_647), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n4248) );
NOR2_X1 MEM_stage_inst_dmem_U4391 ( .A1(MEM_stage_inst_dmem_n4246), .A2(MEM_stage_inst_dmem_n4245), .ZN(MEM_stage_inst_dmem_n4254) );
NAND2_X1 MEM_stage_inst_dmem_U4390 ( .A1(MEM_stage_inst_dmem_n4244), .A2(MEM_stage_inst_dmem_n4243), .ZN(MEM_stage_inst_dmem_n4245) );
NAND2_X1 MEM_stage_inst_dmem_U4389 ( .A1(MEM_stage_inst_dmem_ram_599), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n4243) );
NAND2_X1 MEM_stage_inst_dmem_U4388 ( .A1(MEM_stage_inst_dmem_ram_743), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n4244) );
NAND2_X1 MEM_stage_inst_dmem_U4387 ( .A1(MEM_stage_inst_dmem_n4242), .A2(MEM_stage_inst_dmem_n4241), .ZN(MEM_stage_inst_dmem_n4246) );
NAND2_X1 MEM_stage_inst_dmem_U4386 ( .A1(MEM_stage_inst_dmem_ram_855), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n4241) );
NAND2_X1 MEM_stage_inst_dmem_U4385 ( .A1(MEM_stage_inst_dmem_ram_295), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n4242) );
NAND2_X1 MEM_stage_inst_dmem_U4384 ( .A1(MEM_stage_inst_dmem_n4240), .A2(MEM_stage_inst_dmem_n4239), .ZN(MEM_stage_inst_dmem_n4256) );
NOR2_X1 MEM_stage_inst_dmem_U4383 ( .A1(MEM_stage_inst_dmem_n4238), .A2(MEM_stage_inst_dmem_n4237), .ZN(MEM_stage_inst_dmem_n4239) );
NAND2_X1 MEM_stage_inst_dmem_U4382 ( .A1(MEM_stage_inst_dmem_n4236), .A2(MEM_stage_inst_dmem_n4235), .ZN(MEM_stage_inst_dmem_n4237) );
NAND2_X1 MEM_stage_inst_dmem_U4381 ( .A1(MEM_stage_inst_dmem_ram_71), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n4235) );
NAND2_X1 MEM_stage_inst_dmem_U4380 ( .A1(MEM_stage_inst_dmem_ram_727), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n4236) );
NAND2_X1 MEM_stage_inst_dmem_U4379 ( .A1(MEM_stage_inst_dmem_n4234), .A2(MEM_stage_inst_dmem_n4233), .ZN(MEM_stage_inst_dmem_n4238) );
NAND2_X1 MEM_stage_inst_dmem_U4378 ( .A1(MEM_stage_inst_dmem_ram_503), .A2(MEM_stage_inst_dmem_n64), .ZN(MEM_stage_inst_dmem_n4233) );
NAND2_X1 MEM_stage_inst_dmem_U4377 ( .A1(MEM_stage_inst_dmem_ram_247), .A2(MEM_stage_inst_dmem_n4649), .ZN(MEM_stage_inst_dmem_n4234) );
NOR2_X1 MEM_stage_inst_dmem_U4376 ( .A1(MEM_stage_inst_dmem_n4232), .A2(MEM_stage_inst_dmem_n4231), .ZN(MEM_stage_inst_dmem_n4240) );
NAND2_X1 MEM_stage_inst_dmem_U4375 ( .A1(MEM_stage_inst_dmem_n4230), .A2(MEM_stage_inst_dmem_n4229), .ZN(MEM_stage_inst_dmem_n4231) );
NAND2_X1 MEM_stage_inst_dmem_U4374 ( .A1(MEM_stage_inst_dmem_ram_439), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n4229) );
NAND2_X1 MEM_stage_inst_dmem_U4373 ( .A1(MEM_stage_inst_dmem_ram_679), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n4230) );
NAND2_X1 MEM_stage_inst_dmem_U4372 ( .A1(MEM_stage_inst_dmem_n4228), .A2(MEM_stage_inst_dmem_n4227), .ZN(MEM_stage_inst_dmem_n4232) );
NAND2_X1 MEM_stage_inst_dmem_U4371 ( .A1(MEM_stage_inst_dmem_ram_711), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n4227) );
NAND2_X1 MEM_stage_inst_dmem_U4370 ( .A1(MEM_stage_inst_dmem_ram_631), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n4228) );
NOR2_X1 MEM_stage_inst_dmem_U4369 ( .A1(MEM_stage_inst_dmem_n4226), .A2(MEM_stage_inst_dmem_n4225), .ZN(MEM_stage_inst_dmem_n4258) );
NAND2_X1 MEM_stage_inst_dmem_U4368 ( .A1(MEM_stage_inst_dmem_n4224), .A2(MEM_stage_inst_dmem_n4223), .ZN(MEM_stage_inst_dmem_n4225) );
NOR2_X1 MEM_stage_inst_dmem_U4367 ( .A1(MEM_stage_inst_dmem_n4222), .A2(MEM_stage_inst_dmem_n4221), .ZN(MEM_stage_inst_dmem_n4223) );
NAND2_X1 MEM_stage_inst_dmem_U4366 ( .A1(MEM_stage_inst_dmem_n4220), .A2(MEM_stage_inst_dmem_n4219), .ZN(MEM_stage_inst_dmem_n4221) );
NAND2_X1 MEM_stage_inst_dmem_U4365 ( .A1(MEM_stage_inst_dmem_ram_919), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n4219) );
NAND2_X1 MEM_stage_inst_dmem_U4364 ( .A1(MEM_stage_inst_dmem_ram_119), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n4220) );
NAND2_X1 MEM_stage_inst_dmem_U4363 ( .A1(MEM_stage_inst_dmem_n4218), .A2(MEM_stage_inst_dmem_n4217), .ZN(MEM_stage_inst_dmem_n4222) );
NAND2_X1 MEM_stage_inst_dmem_U4362 ( .A1(MEM_stage_inst_dmem_ram_759), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n4217) );
NAND2_X1 MEM_stage_inst_dmem_U4361 ( .A1(MEM_stage_inst_dmem_ram_983), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n4218) );
NOR2_X1 MEM_stage_inst_dmem_U4360 ( .A1(MEM_stage_inst_dmem_n4216), .A2(MEM_stage_inst_dmem_n4215), .ZN(MEM_stage_inst_dmem_n4224) );
NAND2_X1 MEM_stage_inst_dmem_U4359 ( .A1(MEM_stage_inst_dmem_n4214), .A2(MEM_stage_inst_dmem_n4213), .ZN(MEM_stage_inst_dmem_n4215) );
NAND2_X1 MEM_stage_inst_dmem_U4358 ( .A1(MEM_stage_inst_dmem_ram_135), .A2(MEM_stage_inst_dmem_n61), .ZN(MEM_stage_inst_dmem_n4213) );
NAND2_X1 MEM_stage_inst_dmem_U4357 ( .A1(MEM_stage_inst_dmem_ram_7), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n4214) );
NAND2_X1 MEM_stage_inst_dmem_U4356 ( .A1(MEM_stage_inst_dmem_n4212), .A2(MEM_stage_inst_dmem_n4211), .ZN(MEM_stage_inst_dmem_n4216) );
NAND2_X1 MEM_stage_inst_dmem_U4355 ( .A1(MEM_stage_inst_dmem_ram_199), .A2(MEM_stage_inst_dmem_n36), .ZN(MEM_stage_inst_dmem_n4211) );
NAND2_X1 MEM_stage_inst_dmem_U4354 ( .A1(MEM_stage_inst_dmem_ram_55), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n4212) );
NAND2_X1 MEM_stage_inst_dmem_U4353 ( .A1(MEM_stage_inst_dmem_n4210), .A2(MEM_stage_inst_dmem_n4209), .ZN(MEM_stage_inst_dmem_n4226) );
NOR2_X1 MEM_stage_inst_dmem_U4352 ( .A1(MEM_stage_inst_dmem_n4208), .A2(MEM_stage_inst_dmem_n4207), .ZN(MEM_stage_inst_dmem_n4209) );
NAND2_X1 MEM_stage_inst_dmem_U4351 ( .A1(MEM_stage_inst_dmem_n4206), .A2(MEM_stage_inst_dmem_n4205), .ZN(MEM_stage_inst_dmem_n4207) );
NAND2_X1 MEM_stage_inst_dmem_U4350 ( .A1(MEM_stage_inst_dmem_ram_823), .A2(MEM_stage_inst_dmem_n4740), .ZN(MEM_stage_inst_dmem_n4205) );
NAND2_X1 MEM_stage_inst_dmem_U4349 ( .A1(MEM_stage_inst_dmem_ram_791), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n4206) );
NAND2_X1 MEM_stage_inst_dmem_U4348 ( .A1(MEM_stage_inst_dmem_n4204), .A2(MEM_stage_inst_dmem_n4203), .ZN(MEM_stage_inst_dmem_n4208) );
NAND2_X1 MEM_stage_inst_dmem_U4347 ( .A1(MEM_stage_inst_dmem_ram_567), .A2(MEM_stage_inst_dmem_n41), .ZN(MEM_stage_inst_dmem_n4203) );
NAND2_X1 MEM_stage_inst_dmem_U4346 ( .A1(MEM_stage_inst_dmem_ram_615), .A2(MEM_stage_inst_dmem_n4701), .ZN(MEM_stage_inst_dmem_n4204) );
NOR2_X1 MEM_stage_inst_dmem_U4345 ( .A1(MEM_stage_inst_dmem_n4202), .A2(MEM_stage_inst_dmem_n4201), .ZN(MEM_stage_inst_dmem_n4210) );
NAND2_X1 MEM_stage_inst_dmem_U4344 ( .A1(MEM_stage_inst_dmem_n4200), .A2(MEM_stage_inst_dmem_n4199), .ZN(MEM_stage_inst_dmem_n4201) );
NAND2_X1 MEM_stage_inst_dmem_U4343 ( .A1(MEM_stage_inst_dmem_ram_871), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n4199) );
NAND2_X1 MEM_stage_inst_dmem_U4342 ( .A1(MEM_stage_inst_dmem_ram_167), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n4200) );
NAND2_X1 MEM_stage_inst_dmem_U4341 ( .A1(MEM_stage_inst_dmem_n4198), .A2(MEM_stage_inst_dmem_n4197), .ZN(MEM_stage_inst_dmem_n4202) );
NAND2_X1 MEM_stage_inst_dmem_U4340 ( .A1(MEM_stage_inst_dmem_ram_999), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n4197) );
NAND2_X1 MEM_stage_inst_dmem_U4339 ( .A1(MEM_stage_inst_dmem_ram_343), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n4198) );
NAND2_X1 MEM_stage_inst_dmem_U4338 ( .A1(MEM_stage_inst_dmem_n4196), .A2(MEM_stage_inst_dmem_n4195), .ZN(MEM_stage_inst_dmem_n4260) );
NOR2_X1 MEM_stage_inst_dmem_U4337 ( .A1(MEM_stage_inst_dmem_n4194), .A2(MEM_stage_inst_dmem_n4193), .ZN(MEM_stage_inst_dmem_n4195) );
NAND2_X1 MEM_stage_inst_dmem_U4336 ( .A1(MEM_stage_inst_dmem_n4192), .A2(MEM_stage_inst_dmem_n4191), .ZN(MEM_stage_inst_dmem_n4193) );
NOR2_X1 MEM_stage_inst_dmem_U4335 ( .A1(MEM_stage_inst_dmem_n4190), .A2(MEM_stage_inst_dmem_n4189), .ZN(MEM_stage_inst_dmem_n4191) );
NAND2_X1 MEM_stage_inst_dmem_U4334 ( .A1(MEM_stage_inst_dmem_n4188), .A2(MEM_stage_inst_dmem_n4187), .ZN(MEM_stage_inst_dmem_n4189) );
NAND2_X1 MEM_stage_inst_dmem_U4333 ( .A1(MEM_stage_inst_dmem_ram_151), .A2(MEM_stage_inst_dmem_n5807), .ZN(MEM_stage_inst_dmem_n4187) );
NAND2_X1 MEM_stage_inst_dmem_U4332 ( .A1(MEM_stage_inst_dmem_ram_375), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n4188) );
NAND2_X1 MEM_stage_inst_dmem_U4331 ( .A1(MEM_stage_inst_dmem_n4186), .A2(MEM_stage_inst_dmem_n4185), .ZN(MEM_stage_inst_dmem_n4190) );
NAND2_X1 MEM_stage_inst_dmem_U4330 ( .A1(MEM_stage_inst_dmem_ram_903), .A2(MEM_stage_inst_dmem_n72), .ZN(MEM_stage_inst_dmem_n4185) );
NAND2_X1 MEM_stage_inst_dmem_U4329 ( .A1(MEM_stage_inst_dmem_ram_279), .A2(MEM_stage_inst_dmem_n4672), .ZN(MEM_stage_inst_dmem_n4186) );
NOR2_X1 MEM_stage_inst_dmem_U4328 ( .A1(MEM_stage_inst_dmem_n4184), .A2(MEM_stage_inst_dmem_n4183), .ZN(MEM_stage_inst_dmem_n4192) );
NAND2_X1 MEM_stage_inst_dmem_U4327 ( .A1(MEM_stage_inst_dmem_n4182), .A2(MEM_stage_inst_dmem_n4181), .ZN(MEM_stage_inst_dmem_n4183) );
NAND2_X1 MEM_stage_inst_dmem_U4326 ( .A1(MEM_stage_inst_dmem_ram_535), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n4181) );
NAND2_X1 MEM_stage_inst_dmem_U4325 ( .A1(MEM_stage_inst_dmem_ram_103), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n4182) );
NAND2_X1 MEM_stage_inst_dmem_U4324 ( .A1(MEM_stage_inst_dmem_n4180), .A2(MEM_stage_inst_dmem_n4179), .ZN(MEM_stage_inst_dmem_n4184) );
NAND2_X1 MEM_stage_inst_dmem_U4323 ( .A1(MEM_stage_inst_dmem_ram_311), .A2(MEM_stage_inst_dmem_n4731), .ZN(MEM_stage_inst_dmem_n4179) );
NAND2_X1 MEM_stage_inst_dmem_U4322 ( .A1(MEM_stage_inst_dmem_ram_551), .A2(MEM_stage_inst_dmem_n4692), .ZN(MEM_stage_inst_dmem_n4180) );
NAND2_X1 MEM_stage_inst_dmem_U4321 ( .A1(MEM_stage_inst_dmem_n4178), .A2(MEM_stage_inst_dmem_n4177), .ZN(MEM_stage_inst_dmem_n4194) );
NOR2_X1 MEM_stage_inst_dmem_U4320 ( .A1(MEM_stage_inst_dmem_n4176), .A2(MEM_stage_inst_dmem_n4175), .ZN(MEM_stage_inst_dmem_n4177) );
NAND2_X1 MEM_stage_inst_dmem_U4319 ( .A1(MEM_stage_inst_dmem_n4174), .A2(MEM_stage_inst_dmem_n4173), .ZN(MEM_stage_inst_dmem_n4175) );
NAND2_X1 MEM_stage_inst_dmem_U4318 ( .A1(MEM_stage_inst_dmem_ram_519), .A2(MEM_stage_inst_dmem_n71), .ZN(MEM_stage_inst_dmem_n4173) );
NAND2_X1 MEM_stage_inst_dmem_U4317 ( .A1(MEM_stage_inst_dmem_ram_263), .A2(MEM_stage_inst_dmem_n7898), .ZN(MEM_stage_inst_dmem_n4174) );
NAND2_X1 MEM_stage_inst_dmem_U4316 ( .A1(MEM_stage_inst_dmem_n4172), .A2(MEM_stage_inst_dmem_n4171), .ZN(MEM_stage_inst_dmem_n4176) );
NAND2_X1 MEM_stage_inst_dmem_U4315 ( .A1(MEM_stage_inst_dmem_ram_951), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n4171) );
NAND2_X1 MEM_stage_inst_dmem_U4314 ( .A1(MEM_stage_inst_dmem_ram_1015), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n4172) );
NOR2_X1 MEM_stage_inst_dmem_U4313 ( .A1(MEM_stage_inst_dmem_n4170), .A2(MEM_stage_inst_dmem_n4169), .ZN(MEM_stage_inst_dmem_n4178) );
NAND2_X1 MEM_stage_inst_dmem_U4312 ( .A1(MEM_stage_inst_dmem_n4168), .A2(MEM_stage_inst_dmem_n4167), .ZN(MEM_stage_inst_dmem_n4169) );
NAND2_X1 MEM_stage_inst_dmem_U4311 ( .A1(MEM_stage_inst_dmem_ram_967), .A2(MEM_stage_inst_dmem_n4728), .ZN(MEM_stage_inst_dmem_n4167) );
NAND2_X1 MEM_stage_inst_dmem_U4310 ( .A1(MEM_stage_inst_dmem_ram_215), .A2(MEM_stage_inst_dmem_n51), .ZN(MEM_stage_inst_dmem_n4168) );
NAND2_X1 MEM_stage_inst_dmem_U4309 ( .A1(MEM_stage_inst_dmem_n4166), .A2(MEM_stage_inst_dmem_n4165), .ZN(MEM_stage_inst_dmem_n4170) );
NAND2_X1 MEM_stage_inst_dmem_U4308 ( .A1(MEM_stage_inst_dmem_ram_839), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n4165) );
NAND2_X1 MEM_stage_inst_dmem_U4307 ( .A1(MEM_stage_inst_dmem_ram_807), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n4166) );
NOR2_X1 MEM_stage_inst_dmem_U4306 ( .A1(MEM_stage_inst_dmem_n4164), .A2(MEM_stage_inst_dmem_n4163), .ZN(MEM_stage_inst_dmem_n4196) );
NAND2_X1 MEM_stage_inst_dmem_U4305 ( .A1(MEM_stage_inst_dmem_n4162), .A2(MEM_stage_inst_dmem_n4161), .ZN(MEM_stage_inst_dmem_n4163) );
NOR2_X1 MEM_stage_inst_dmem_U4304 ( .A1(MEM_stage_inst_dmem_n4160), .A2(MEM_stage_inst_dmem_n4159), .ZN(MEM_stage_inst_dmem_n4161) );
NAND2_X1 MEM_stage_inst_dmem_U4303 ( .A1(MEM_stage_inst_dmem_n4158), .A2(MEM_stage_inst_dmem_n4157), .ZN(MEM_stage_inst_dmem_n4159) );
NAND2_X1 MEM_stage_inst_dmem_U4302 ( .A1(MEM_stage_inst_dmem_ram_423), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n4157) );
NAND2_X1 MEM_stage_inst_dmem_U4301 ( .A1(MEM_stage_inst_dmem_ram_455), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n4158) );
NAND2_X1 MEM_stage_inst_dmem_U4300 ( .A1(MEM_stage_inst_dmem_n4156), .A2(MEM_stage_inst_dmem_n4155), .ZN(MEM_stage_inst_dmem_n4160) );
NAND2_X1 MEM_stage_inst_dmem_U4299 ( .A1(MEM_stage_inst_dmem_ram_87), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n4155) );
NAND2_X1 MEM_stage_inst_dmem_U4298 ( .A1(MEM_stage_inst_dmem_ram_663), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n4156) );
NOR2_X1 MEM_stage_inst_dmem_U4297 ( .A1(MEM_stage_inst_dmem_n4154), .A2(MEM_stage_inst_dmem_n4153), .ZN(MEM_stage_inst_dmem_n4162) );
NAND2_X1 MEM_stage_inst_dmem_U4296 ( .A1(MEM_stage_inst_dmem_n4152), .A2(MEM_stage_inst_dmem_n4151), .ZN(MEM_stage_inst_dmem_n4153) );
NAND2_X1 MEM_stage_inst_dmem_U4295 ( .A1(MEM_stage_inst_dmem_ram_487), .A2(MEM_stage_inst_dmem_n4667), .ZN(MEM_stage_inst_dmem_n4151) );
NAND2_X1 MEM_stage_inst_dmem_U4294 ( .A1(MEM_stage_inst_dmem_ram_23), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n4152) );
NAND2_X1 MEM_stage_inst_dmem_U4293 ( .A1(MEM_stage_inst_dmem_n4150), .A2(MEM_stage_inst_dmem_n4149), .ZN(MEM_stage_inst_dmem_n4154) );
NAND2_X1 MEM_stage_inst_dmem_U4292 ( .A1(MEM_stage_inst_dmem_ram_471), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n4149) );
NAND2_X1 MEM_stage_inst_dmem_U4291 ( .A1(MEM_stage_inst_dmem_ram_391), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n4150) );
NAND2_X1 MEM_stage_inst_dmem_U4290 ( .A1(MEM_stage_inst_dmem_n4148), .A2(MEM_stage_inst_dmem_n4147), .ZN(MEM_stage_inst_dmem_n4164) );
NOR2_X1 MEM_stage_inst_dmem_U4289 ( .A1(MEM_stage_inst_dmem_n4146), .A2(MEM_stage_inst_dmem_n4145), .ZN(MEM_stage_inst_dmem_n4147) );
NAND2_X1 MEM_stage_inst_dmem_U4288 ( .A1(MEM_stage_inst_dmem_n4144), .A2(MEM_stage_inst_dmem_n4143), .ZN(MEM_stage_inst_dmem_n4145) );
NAND2_X1 MEM_stage_inst_dmem_U4287 ( .A1(MEM_stage_inst_dmem_ram_39), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n4143) );
NAND2_X1 MEM_stage_inst_dmem_U4286 ( .A1(MEM_stage_inst_dmem_ram_935), .A2(MEM_stage_inst_dmem_n4675), .ZN(MEM_stage_inst_dmem_n4144) );
NAND2_X1 MEM_stage_inst_dmem_U4285 ( .A1(MEM_stage_inst_dmem_n4142), .A2(MEM_stage_inst_dmem_n4141), .ZN(MEM_stage_inst_dmem_n4146) );
NAND2_X1 MEM_stage_inst_dmem_U4284 ( .A1(MEM_stage_inst_dmem_ram_775), .A2(MEM_stage_inst_dmem_n37), .ZN(MEM_stage_inst_dmem_n4141) );
NAND2_X1 MEM_stage_inst_dmem_U4283 ( .A1(MEM_stage_inst_dmem_ram_359), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n4142) );
NOR2_X1 MEM_stage_inst_dmem_U4282 ( .A1(MEM_stage_inst_dmem_n4140), .A2(MEM_stage_inst_dmem_n4139), .ZN(MEM_stage_inst_dmem_n4148) );
NAND2_X1 MEM_stage_inst_dmem_U4281 ( .A1(MEM_stage_inst_dmem_n4138), .A2(MEM_stage_inst_dmem_n4137), .ZN(MEM_stage_inst_dmem_n4139) );
NAND2_X1 MEM_stage_inst_dmem_U4280 ( .A1(MEM_stage_inst_dmem_ram_887), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n4137) );
NAND2_X1 MEM_stage_inst_dmem_U4279 ( .A1(MEM_stage_inst_dmem_ram_327), .A2(MEM_stage_inst_dmem_n4706), .ZN(MEM_stage_inst_dmem_n4138) );
NAND2_X1 MEM_stage_inst_dmem_U4278 ( .A1(MEM_stage_inst_dmem_n4136), .A2(MEM_stage_inst_dmem_n4135), .ZN(MEM_stage_inst_dmem_n4140) );
NAND2_X1 MEM_stage_inst_dmem_U4277 ( .A1(MEM_stage_inst_dmem_ram_407), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n4135) );
NAND2_X1 MEM_stage_inst_dmem_U4276 ( .A1(MEM_stage_inst_dmem_ram_183), .A2(MEM_stage_inst_dmem_n55), .ZN(MEM_stage_inst_dmem_n4136) );
NOR2_X1 MEM_stage_inst_dmem_U4275 ( .A1(MEM_stage_inst_dmem_n4134), .A2(MEM_stage_inst_dmem_n4133), .ZN(MEM_stage_inst_dmem_n4392) );
NOR2_X1 MEM_stage_inst_dmem_U4274 ( .A1(MEM_stage_inst_dmem_n4132), .A2(MEM_stage_inst_dmem_n8286), .ZN(MEM_stage_inst_dmem_n4133) );
NOR2_X1 MEM_stage_inst_dmem_U4273 ( .A1(MEM_stage_inst_dmem_n4131), .A2(MEM_stage_inst_dmem_n4130), .ZN(MEM_stage_inst_dmem_n4132) );
NAND2_X1 MEM_stage_inst_dmem_U4272 ( .A1(MEM_stage_inst_dmem_n4129), .A2(MEM_stage_inst_dmem_n4128), .ZN(MEM_stage_inst_dmem_n4130) );
NOR2_X1 MEM_stage_inst_dmem_U4271 ( .A1(MEM_stage_inst_dmem_n4127), .A2(MEM_stage_inst_dmem_n4126), .ZN(MEM_stage_inst_dmem_n4128) );
NAND2_X1 MEM_stage_inst_dmem_U4270 ( .A1(MEM_stage_inst_dmem_n4125), .A2(MEM_stage_inst_dmem_n4124), .ZN(MEM_stage_inst_dmem_n4126) );
NOR2_X1 MEM_stage_inst_dmem_U4269 ( .A1(MEM_stage_inst_dmem_n4123), .A2(MEM_stage_inst_dmem_n4122), .ZN(MEM_stage_inst_dmem_n4124) );
NAND2_X1 MEM_stage_inst_dmem_U4268 ( .A1(MEM_stage_inst_dmem_n4121), .A2(MEM_stage_inst_dmem_n4120), .ZN(MEM_stage_inst_dmem_n4122) );
NAND2_X1 MEM_stage_inst_dmem_U4267 ( .A1(MEM_stage_inst_dmem_ram_2759), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n4120) );
NAND2_X1 MEM_stage_inst_dmem_U4266 ( .A1(MEM_stage_inst_dmem_ram_2343), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n4121) );
NAND2_X1 MEM_stage_inst_dmem_U4265 ( .A1(MEM_stage_inst_dmem_n4119), .A2(MEM_stage_inst_dmem_n4118), .ZN(MEM_stage_inst_dmem_n4123) );
NAND2_X1 MEM_stage_inst_dmem_U4264 ( .A1(MEM_stage_inst_dmem_ram_2295), .A2(MEM_stage_inst_dmem_n39), .ZN(MEM_stage_inst_dmem_n4118) );
NAND2_X1 MEM_stage_inst_dmem_U4263 ( .A1(MEM_stage_inst_dmem_ram_2839), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n4119) );
NOR2_X1 MEM_stage_inst_dmem_U4262 ( .A1(MEM_stage_inst_dmem_n4117), .A2(MEM_stage_inst_dmem_n4116), .ZN(MEM_stage_inst_dmem_n4125) );
NAND2_X1 MEM_stage_inst_dmem_U4261 ( .A1(MEM_stage_inst_dmem_n4115), .A2(MEM_stage_inst_dmem_n4114), .ZN(MEM_stage_inst_dmem_n4116) );
NAND2_X1 MEM_stage_inst_dmem_U4260 ( .A1(MEM_stage_inst_dmem_ram_2519), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n4114) );
NAND2_X1 MEM_stage_inst_dmem_U4259 ( .A1(MEM_stage_inst_dmem_ram_2055), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n4115) );
NAND2_X1 MEM_stage_inst_dmem_U4258 ( .A1(MEM_stage_inst_dmem_n4113), .A2(MEM_stage_inst_dmem_n4112), .ZN(MEM_stage_inst_dmem_n4117) );
NAND2_X1 MEM_stage_inst_dmem_U4257 ( .A1(MEM_stage_inst_dmem_ram_2263), .A2(MEM_stage_inst_dmem_n51), .ZN(MEM_stage_inst_dmem_n4112) );
NAND2_X1 MEM_stage_inst_dmem_U4256 ( .A1(MEM_stage_inst_dmem_ram_2391), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n4113) );
NAND2_X1 MEM_stage_inst_dmem_U4255 ( .A1(MEM_stage_inst_dmem_n4111), .A2(MEM_stage_inst_dmem_n4110), .ZN(MEM_stage_inst_dmem_n4127) );
NOR2_X1 MEM_stage_inst_dmem_U4254 ( .A1(MEM_stage_inst_dmem_n4109), .A2(MEM_stage_inst_dmem_n4108), .ZN(MEM_stage_inst_dmem_n4110) );
NAND2_X1 MEM_stage_inst_dmem_U4253 ( .A1(MEM_stage_inst_dmem_n4107), .A2(MEM_stage_inst_dmem_n4106), .ZN(MEM_stage_inst_dmem_n4108) );
NAND2_X1 MEM_stage_inst_dmem_U4252 ( .A1(MEM_stage_inst_dmem_ram_2455), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n4106) );
NAND2_X1 MEM_stage_inst_dmem_U4251 ( .A1(MEM_stage_inst_dmem_ram_2119), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n4107) );
NAND2_X1 MEM_stage_inst_dmem_U4250 ( .A1(MEM_stage_inst_dmem_n4105), .A2(MEM_stage_inst_dmem_n4104), .ZN(MEM_stage_inst_dmem_n4109) );
NAND2_X1 MEM_stage_inst_dmem_U4249 ( .A1(MEM_stage_inst_dmem_ram_2375), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n4104) );
NAND2_X1 MEM_stage_inst_dmem_U4248 ( .A1(MEM_stage_inst_dmem_ram_2487), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n4105) );
NOR2_X1 MEM_stage_inst_dmem_U4247 ( .A1(MEM_stage_inst_dmem_n4103), .A2(MEM_stage_inst_dmem_n4102), .ZN(MEM_stage_inst_dmem_n4111) );
NAND2_X1 MEM_stage_inst_dmem_U4246 ( .A1(MEM_stage_inst_dmem_n4101), .A2(MEM_stage_inst_dmem_n4100), .ZN(MEM_stage_inst_dmem_n4102) );
NAND2_X1 MEM_stage_inst_dmem_U4245 ( .A1(MEM_stage_inst_dmem_ram_3031), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n4100) );
NAND2_X1 MEM_stage_inst_dmem_U4244 ( .A1(MEM_stage_inst_dmem_ram_2791), .A2(MEM_stage_inst_dmem_n4769), .ZN(MEM_stage_inst_dmem_n4101) );
NAND2_X1 MEM_stage_inst_dmem_U4243 ( .A1(MEM_stage_inst_dmem_n4099), .A2(MEM_stage_inst_dmem_n4098), .ZN(MEM_stage_inst_dmem_n4103) );
NAND2_X1 MEM_stage_inst_dmem_U4242 ( .A1(MEM_stage_inst_dmem_ram_2935), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n4098) );
NAND2_X1 MEM_stage_inst_dmem_U4241 ( .A1(MEM_stage_inst_dmem_ram_2167), .A2(MEM_stage_inst_dmem_n4710), .ZN(MEM_stage_inst_dmem_n4099) );
NOR2_X1 MEM_stage_inst_dmem_U4240 ( .A1(MEM_stage_inst_dmem_n4097), .A2(MEM_stage_inst_dmem_n4096), .ZN(MEM_stage_inst_dmem_n4129) );
NAND2_X1 MEM_stage_inst_dmem_U4239 ( .A1(MEM_stage_inst_dmem_n4095), .A2(MEM_stage_inst_dmem_n4094), .ZN(MEM_stage_inst_dmem_n4096) );
NOR2_X1 MEM_stage_inst_dmem_U4238 ( .A1(MEM_stage_inst_dmem_n4093), .A2(MEM_stage_inst_dmem_n4092), .ZN(MEM_stage_inst_dmem_n4094) );
NAND2_X1 MEM_stage_inst_dmem_U4237 ( .A1(MEM_stage_inst_dmem_n4091), .A2(MEM_stage_inst_dmem_n4090), .ZN(MEM_stage_inst_dmem_n4092) );
NAND2_X1 MEM_stage_inst_dmem_U4236 ( .A1(MEM_stage_inst_dmem_ram_2615), .A2(MEM_stage_inst_dmem_n41), .ZN(MEM_stage_inst_dmem_n4090) );
NAND2_X1 MEM_stage_inst_dmem_U4235 ( .A1(MEM_stage_inst_dmem_ram_2439), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n4091) );
NAND2_X1 MEM_stage_inst_dmem_U4234 ( .A1(MEM_stage_inst_dmem_n4089), .A2(MEM_stage_inst_dmem_n4088), .ZN(MEM_stage_inst_dmem_n4093) );
NAND2_X1 MEM_stage_inst_dmem_U4233 ( .A1(MEM_stage_inst_dmem_ram_2423), .A2(MEM_stage_inst_dmem_n4721), .ZN(MEM_stage_inst_dmem_n4088) );
NAND2_X1 MEM_stage_inst_dmem_U4232 ( .A1(MEM_stage_inst_dmem_ram_2711), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n4089) );
NOR2_X1 MEM_stage_inst_dmem_U4231 ( .A1(MEM_stage_inst_dmem_n4087), .A2(MEM_stage_inst_dmem_n4086), .ZN(MEM_stage_inst_dmem_n4095) );
NAND2_X1 MEM_stage_inst_dmem_U4230 ( .A1(MEM_stage_inst_dmem_n4085), .A2(MEM_stage_inst_dmem_n4084), .ZN(MEM_stage_inst_dmem_n4086) );
NAND2_X1 MEM_stage_inst_dmem_U4229 ( .A1(MEM_stage_inst_dmem_ram_3015), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n4084) );
NAND2_X1 MEM_stage_inst_dmem_U4228 ( .A1(MEM_stage_inst_dmem_ram_2871), .A2(MEM_stage_inst_dmem_n46), .ZN(MEM_stage_inst_dmem_n4085) );
NAND2_X1 MEM_stage_inst_dmem_U4227 ( .A1(MEM_stage_inst_dmem_n4083), .A2(MEM_stage_inst_dmem_n4082), .ZN(MEM_stage_inst_dmem_n4087) );
NAND2_X1 MEM_stage_inst_dmem_U4226 ( .A1(MEM_stage_inst_dmem_ram_2983), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n4082) );
NAND2_X1 MEM_stage_inst_dmem_U4225 ( .A1(MEM_stage_inst_dmem_ram_2631), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n4083) );
NAND2_X1 MEM_stage_inst_dmem_U4224 ( .A1(MEM_stage_inst_dmem_n4081), .A2(MEM_stage_inst_dmem_n4080), .ZN(MEM_stage_inst_dmem_n4097) );
NOR2_X1 MEM_stage_inst_dmem_U4223 ( .A1(MEM_stage_inst_dmem_n4079), .A2(MEM_stage_inst_dmem_n4078), .ZN(MEM_stage_inst_dmem_n4080) );
NAND2_X1 MEM_stage_inst_dmem_U4222 ( .A1(MEM_stage_inst_dmem_n4077), .A2(MEM_stage_inst_dmem_n4076), .ZN(MEM_stage_inst_dmem_n4078) );
NAND2_X1 MEM_stage_inst_dmem_U4221 ( .A1(MEM_stage_inst_dmem_ram_2743), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n4076) );
NAND2_X1 MEM_stage_inst_dmem_U4220 ( .A1(MEM_stage_inst_dmem_ram_2199), .A2(MEM_stage_inst_dmem_n5807), .ZN(MEM_stage_inst_dmem_n4077) );
NAND2_X1 MEM_stage_inst_dmem_U4219 ( .A1(MEM_stage_inst_dmem_n4075), .A2(MEM_stage_inst_dmem_n4074), .ZN(MEM_stage_inst_dmem_n4079) );
NAND2_X1 MEM_stage_inst_dmem_U4218 ( .A1(MEM_stage_inst_dmem_ram_2919), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n4074) );
NAND2_X1 MEM_stage_inst_dmem_U4217 ( .A1(MEM_stage_inst_dmem_ram_2071), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n4075) );
NOR2_X1 MEM_stage_inst_dmem_U4216 ( .A1(MEM_stage_inst_dmem_n4073), .A2(MEM_stage_inst_dmem_n4072), .ZN(MEM_stage_inst_dmem_n4081) );
NAND2_X1 MEM_stage_inst_dmem_U4215 ( .A1(MEM_stage_inst_dmem_n4071), .A2(MEM_stage_inst_dmem_n4070), .ZN(MEM_stage_inst_dmem_n4072) );
NAND2_X1 MEM_stage_inst_dmem_U4214 ( .A1(MEM_stage_inst_dmem_ram_2855), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n4070) );
NAND2_X1 MEM_stage_inst_dmem_U4213 ( .A1(MEM_stage_inst_dmem_ram_2727), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n4071) );
NAND2_X1 MEM_stage_inst_dmem_U4212 ( .A1(MEM_stage_inst_dmem_n4069), .A2(MEM_stage_inst_dmem_n4068), .ZN(MEM_stage_inst_dmem_n4073) );
NAND2_X1 MEM_stage_inst_dmem_U4211 ( .A1(MEM_stage_inst_dmem_ram_2183), .A2(MEM_stage_inst_dmem_n61), .ZN(MEM_stage_inst_dmem_n4068) );
NAND2_X1 MEM_stage_inst_dmem_U4210 ( .A1(MEM_stage_inst_dmem_ram_2327), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n4069) );
NAND2_X1 MEM_stage_inst_dmem_U4209 ( .A1(MEM_stage_inst_dmem_n4067), .A2(MEM_stage_inst_dmem_n4066), .ZN(MEM_stage_inst_dmem_n4131) );
NOR2_X1 MEM_stage_inst_dmem_U4208 ( .A1(MEM_stage_inst_dmem_n4065), .A2(MEM_stage_inst_dmem_n4064), .ZN(MEM_stage_inst_dmem_n4066) );
NAND2_X1 MEM_stage_inst_dmem_U4207 ( .A1(MEM_stage_inst_dmem_n4063), .A2(MEM_stage_inst_dmem_n4062), .ZN(MEM_stage_inst_dmem_n4064) );
NOR2_X1 MEM_stage_inst_dmem_U4206 ( .A1(MEM_stage_inst_dmem_n4061), .A2(MEM_stage_inst_dmem_n4060), .ZN(MEM_stage_inst_dmem_n4062) );
NAND2_X1 MEM_stage_inst_dmem_U4205 ( .A1(MEM_stage_inst_dmem_n4059), .A2(MEM_stage_inst_dmem_n4058), .ZN(MEM_stage_inst_dmem_n4060) );
NAND2_X1 MEM_stage_inst_dmem_U4204 ( .A1(MEM_stage_inst_dmem_ram_2903), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n4058) );
NAND2_X1 MEM_stage_inst_dmem_U4203 ( .A1(MEM_stage_inst_dmem_ram_2471), .A2(MEM_stage_inst_dmem_n4772), .ZN(MEM_stage_inst_dmem_n4059) );
NAND2_X1 MEM_stage_inst_dmem_U4202 ( .A1(MEM_stage_inst_dmem_n4057), .A2(MEM_stage_inst_dmem_n4056), .ZN(MEM_stage_inst_dmem_n4061) );
NAND2_X1 MEM_stage_inst_dmem_U4201 ( .A1(MEM_stage_inst_dmem_ram_2679), .A2(MEM_stage_inst_dmem_n4652), .ZN(MEM_stage_inst_dmem_n4056) );
NAND2_X1 MEM_stage_inst_dmem_U4200 ( .A1(MEM_stage_inst_dmem_ram_2311), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n4057) );
NOR2_X1 MEM_stage_inst_dmem_U4199 ( .A1(MEM_stage_inst_dmem_n4055), .A2(MEM_stage_inst_dmem_n4054), .ZN(MEM_stage_inst_dmem_n4063) );
NAND2_X1 MEM_stage_inst_dmem_U4198 ( .A1(MEM_stage_inst_dmem_n4053), .A2(MEM_stage_inst_dmem_n4052), .ZN(MEM_stage_inst_dmem_n4054) );
NAND2_X1 MEM_stage_inst_dmem_U4197 ( .A1(MEM_stage_inst_dmem_ram_2967), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n4052) );
NAND2_X1 MEM_stage_inst_dmem_U4196 ( .A1(MEM_stage_inst_dmem_ram_2567), .A2(MEM_stage_inst_dmem_n71), .ZN(MEM_stage_inst_dmem_n4053) );
NAND2_X1 MEM_stage_inst_dmem_U4195 ( .A1(MEM_stage_inst_dmem_n4051), .A2(MEM_stage_inst_dmem_n4050), .ZN(MEM_stage_inst_dmem_n4055) );
NAND2_X1 MEM_stage_inst_dmem_U4194 ( .A1(MEM_stage_inst_dmem_ram_2951), .A2(MEM_stage_inst_dmem_n72), .ZN(MEM_stage_inst_dmem_n4050) );
NAND2_X1 MEM_stage_inst_dmem_U4193 ( .A1(MEM_stage_inst_dmem_ram_2135), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n4051) );
NAND2_X1 MEM_stage_inst_dmem_U4192 ( .A1(MEM_stage_inst_dmem_n4049), .A2(MEM_stage_inst_dmem_n4048), .ZN(MEM_stage_inst_dmem_n4065) );
NOR2_X1 MEM_stage_inst_dmem_U4191 ( .A1(MEM_stage_inst_dmem_n4047), .A2(MEM_stage_inst_dmem_n4046), .ZN(MEM_stage_inst_dmem_n4048) );
NAND2_X1 MEM_stage_inst_dmem_U4190 ( .A1(MEM_stage_inst_dmem_n4045), .A2(MEM_stage_inst_dmem_n4044), .ZN(MEM_stage_inst_dmem_n4046) );
NAND2_X1 MEM_stage_inst_dmem_U4189 ( .A1(MEM_stage_inst_dmem_ram_2279), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n4044) );
NAND2_X1 MEM_stage_inst_dmem_U4188 ( .A1(MEM_stage_inst_dmem_ram_2151), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n4045) );
NAND2_X1 MEM_stage_inst_dmem_U4187 ( .A1(MEM_stage_inst_dmem_n4043), .A2(MEM_stage_inst_dmem_n4042), .ZN(MEM_stage_inst_dmem_n4047) );
NAND2_X1 MEM_stage_inst_dmem_U4186 ( .A1(MEM_stage_inst_dmem_ram_2823), .A2(MEM_stage_inst_dmem_n37), .ZN(MEM_stage_inst_dmem_n4042) );
NAND2_X1 MEM_stage_inst_dmem_U4185 ( .A1(MEM_stage_inst_dmem_ram_2231), .A2(MEM_stage_inst_dmem_n55), .ZN(MEM_stage_inst_dmem_n4043) );
NOR2_X1 MEM_stage_inst_dmem_U4184 ( .A1(MEM_stage_inst_dmem_n4041), .A2(MEM_stage_inst_dmem_n4040), .ZN(MEM_stage_inst_dmem_n4049) );
NAND2_X1 MEM_stage_inst_dmem_U4183 ( .A1(MEM_stage_inst_dmem_n4039), .A2(MEM_stage_inst_dmem_n4038), .ZN(MEM_stage_inst_dmem_n4040) );
NAND2_X1 MEM_stage_inst_dmem_U4182 ( .A1(MEM_stage_inst_dmem_ram_2599), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n4038) );
NAND2_X1 MEM_stage_inst_dmem_U4181 ( .A1(MEM_stage_inst_dmem_ram_2663), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n4039) );
NAND2_X1 MEM_stage_inst_dmem_U4180 ( .A1(MEM_stage_inst_dmem_n4037), .A2(MEM_stage_inst_dmem_n4036), .ZN(MEM_stage_inst_dmem_n4041) );
NAND2_X1 MEM_stage_inst_dmem_U4179 ( .A1(MEM_stage_inst_dmem_ram_2359), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n4036) );
NAND2_X1 MEM_stage_inst_dmem_U4178 ( .A1(MEM_stage_inst_dmem_ram_2647), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n4037) );
NOR2_X1 MEM_stage_inst_dmem_U4177 ( .A1(MEM_stage_inst_dmem_n4035), .A2(MEM_stage_inst_dmem_n4034), .ZN(MEM_stage_inst_dmem_n4067) );
NAND2_X1 MEM_stage_inst_dmem_U4176 ( .A1(MEM_stage_inst_dmem_n4033), .A2(MEM_stage_inst_dmem_n4032), .ZN(MEM_stage_inst_dmem_n4034) );
NOR2_X1 MEM_stage_inst_dmem_U4175 ( .A1(MEM_stage_inst_dmem_n4031), .A2(MEM_stage_inst_dmem_n4030), .ZN(MEM_stage_inst_dmem_n4032) );
NAND2_X1 MEM_stage_inst_dmem_U4174 ( .A1(MEM_stage_inst_dmem_n4029), .A2(MEM_stage_inst_dmem_n4028), .ZN(MEM_stage_inst_dmem_n4030) );
NAND2_X1 MEM_stage_inst_dmem_U4173 ( .A1(MEM_stage_inst_dmem_ram_2551), .A2(MEM_stage_inst_dmem_n64), .ZN(MEM_stage_inst_dmem_n4028) );
NAND2_X1 MEM_stage_inst_dmem_U4172 ( .A1(MEM_stage_inst_dmem_ram_2583), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n4029) );
NAND2_X1 MEM_stage_inst_dmem_U4171 ( .A1(MEM_stage_inst_dmem_n4027), .A2(MEM_stage_inst_dmem_n4026), .ZN(MEM_stage_inst_dmem_n4031) );
NAND2_X1 MEM_stage_inst_dmem_U4170 ( .A1(MEM_stage_inst_dmem_ram_2407), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n4026) );
NAND2_X1 MEM_stage_inst_dmem_U4169 ( .A1(MEM_stage_inst_dmem_ram_3063), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n4027) );
NOR2_X1 MEM_stage_inst_dmem_U4168 ( .A1(MEM_stage_inst_dmem_n4025), .A2(MEM_stage_inst_dmem_n4024), .ZN(MEM_stage_inst_dmem_n4033) );
NAND2_X1 MEM_stage_inst_dmem_U4167 ( .A1(MEM_stage_inst_dmem_n4023), .A2(MEM_stage_inst_dmem_n4022), .ZN(MEM_stage_inst_dmem_n4024) );
NAND2_X1 MEM_stage_inst_dmem_U4166 ( .A1(MEM_stage_inst_dmem_ram_2535), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n4022) );
NAND2_X1 MEM_stage_inst_dmem_U4165 ( .A1(MEM_stage_inst_dmem_ram_3047), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n4023) );
NAND2_X1 MEM_stage_inst_dmem_U4164 ( .A1(MEM_stage_inst_dmem_n4021), .A2(MEM_stage_inst_dmem_n4020), .ZN(MEM_stage_inst_dmem_n4025) );
NAND2_X1 MEM_stage_inst_dmem_U4163 ( .A1(MEM_stage_inst_dmem_ram_2807), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n4020) );
NAND2_X1 MEM_stage_inst_dmem_U4162 ( .A1(MEM_stage_inst_dmem_ram_2215), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n4021) );
NAND2_X1 MEM_stage_inst_dmem_U4161 ( .A1(MEM_stage_inst_dmem_n4019), .A2(MEM_stage_inst_dmem_n4018), .ZN(MEM_stage_inst_dmem_n4035) );
NOR2_X1 MEM_stage_inst_dmem_U4160 ( .A1(MEM_stage_inst_dmem_n4017), .A2(MEM_stage_inst_dmem_n4016), .ZN(MEM_stage_inst_dmem_n4018) );
NAND2_X1 MEM_stage_inst_dmem_U4159 ( .A1(MEM_stage_inst_dmem_n4015), .A2(MEM_stage_inst_dmem_n4014), .ZN(MEM_stage_inst_dmem_n4016) );
NAND2_X1 MEM_stage_inst_dmem_U4158 ( .A1(MEM_stage_inst_dmem_ram_2247), .A2(MEM_stage_inst_dmem_n36), .ZN(MEM_stage_inst_dmem_n4014) );
NAND2_X1 MEM_stage_inst_dmem_U4157 ( .A1(MEM_stage_inst_dmem_ram_2503), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n4015) );
NAND2_X1 MEM_stage_inst_dmem_U4156 ( .A1(MEM_stage_inst_dmem_n4013), .A2(MEM_stage_inst_dmem_n4012), .ZN(MEM_stage_inst_dmem_n4017) );
NAND2_X1 MEM_stage_inst_dmem_U4155 ( .A1(MEM_stage_inst_dmem_ram_2887), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n4012) );
NAND2_X1 MEM_stage_inst_dmem_U4154 ( .A1(MEM_stage_inst_dmem_ram_2087), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n4013) );
NOR2_X1 MEM_stage_inst_dmem_U4153 ( .A1(MEM_stage_inst_dmem_n4011), .A2(MEM_stage_inst_dmem_n4010), .ZN(MEM_stage_inst_dmem_n4019) );
NAND2_X1 MEM_stage_inst_dmem_U4152 ( .A1(MEM_stage_inst_dmem_n4009), .A2(MEM_stage_inst_dmem_n4008), .ZN(MEM_stage_inst_dmem_n4010) );
NAND2_X1 MEM_stage_inst_dmem_U4151 ( .A1(MEM_stage_inst_dmem_ram_2103), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n4008) );
NAND2_X1 MEM_stage_inst_dmem_U4150 ( .A1(MEM_stage_inst_dmem_ram_2999), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n4009) );
NAND2_X1 MEM_stage_inst_dmem_U4149 ( .A1(MEM_stage_inst_dmem_n4007), .A2(MEM_stage_inst_dmem_n4006), .ZN(MEM_stage_inst_dmem_n4011) );
NAND2_X1 MEM_stage_inst_dmem_U4148 ( .A1(MEM_stage_inst_dmem_ram_2695), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n4006) );
NAND2_X1 MEM_stage_inst_dmem_U4147 ( .A1(MEM_stage_inst_dmem_ram_2775), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n4007) );
NOR2_X1 MEM_stage_inst_dmem_U4146 ( .A1(MEM_stage_inst_dmem_n4005), .A2(MEM_stage_inst_dmem_n8417), .ZN(MEM_stage_inst_dmem_n4134) );
NOR2_X1 MEM_stage_inst_dmem_U4145 ( .A1(MEM_stage_inst_dmem_n4004), .A2(MEM_stage_inst_dmem_n4003), .ZN(MEM_stage_inst_dmem_n4005) );
NAND2_X1 MEM_stage_inst_dmem_U4144 ( .A1(MEM_stage_inst_dmem_n4002), .A2(MEM_stage_inst_dmem_n4001), .ZN(MEM_stage_inst_dmem_n4003) );
NOR2_X1 MEM_stage_inst_dmem_U4143 ( .A1(MEM_stage_inst_dmem_n4000), .A2(MEM_stage_inst_dmem_n3999), .ZN(MEM_stage_inst_dmem_n4001) );
NAND2_X1 MEM_stage_inst_dmem_U4142 ( .A1(MEM_stage_inst_dmem_n3998), .A2(MEM_stage_inst_dmem_n3997), .ZN(MEM_stage_inst_dmem_n3999) );
NOR2_X1 MEM_stage_inst_dmem_U4141 ( .A1(MEM_stage_inst_dmem_n3996), .A2(MEM_stage_inst_dmem_n3995), .ZN(MEM_stage_inst_dmem_n3997) );
NAND2_X1 MEM_stage_inst_dmem_U4140 ( .A1(MEM_stage_inst_dmem_n3994), .A2(MEM_stage_inst_dmem_n3993), .ZN(MEM_stage_inst_dmem_n3995) );
NAND2_X1 MEM_stage_inst_dmem_U4139 ( .A1(MEM_stage_inst_dmem_ram_3351), .A2(MEM_stage_inst_dmem_n4672), .ZN(MEM_stage_inst_dmem_n3993) );
NAND2_X1 MEM_stage_inst_dmem_U4138 ( .A1(MEM_stage_inst_dmem_ram_3079), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n3994) );
NAND2_X1 MEM_stage_inst_dmem_U4137 ( .A1(MEM_stage_inst_dmem_n3992), .A2(MEM_stage_inst_dmem_n3991), .ZN(MEM_stage_inst_dmem_n3996) );
NAND2_X1 MEM_stage_inst_dmem_U4136 ( .A1(MEM_stage_inst_dmem_ram_3879), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n3991) );
NAND2_X1 MEM_stage_inst_dmem_U4135 ( .A1(MEM_stage_inst_dmem_ram_3159), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n3992) );
NOR2_X1 MEM_stage_inst_dmem_U4134 ( .A1(MEM_stage_inst_dmem_n3990), .A2(MEM_stage_inst_dmem_n3989), .ZN(MEM_stage_inst_dmem_n3998) );
NAND2_X1 MEM_stage_inst_dmem_U4133 ( .A1(MEM_stage_inst_dmem_n3988), .A2(MEM_stage_inst_dmem_n3987), .ZN(MEM_stage_inst_dmem_n3989) );
NAND2_X1 MEM_stage_inst_dmem_U4132 ( .A1(MEM_stage_inst_dmem_ram_4071), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n3987) );
NAND2_X1 MEM_stage_inst_dmem_U4131 ( .A1(MEM_stage_inst_dmem_ram_3367), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n3988) );
NAND2_X1 MEM_stage_inst_dmem_U4130 ( .A1(MEM_stage_inst_dmem_n3986), .A2(MEM_stage_inst_dmem_n3985), .ZN(MEM_stage_inst_dmem_n3990) );
NAND2_X1 MEM_stage_inst_dmem_U4129 ( .A1(MEM_stage_inst_dmem_ram_3543), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n3985) );
NAND2_X1 MEM_stage_inst_dmem_U4128 ( .A1(MEM_stage_inst_dmem_ram_3463), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n3986) );
NAND2_X1 MEM_stage_inst_dmem_U4127 ( .A1(MEM_stage_inst_dmem_n3984), .A2(MEM_stage_inst_dmem_n3983), .ZN(MEM_stage_inst_dmem_n4000) );
NOR2_X1 MEM_stage_inst_dmem_U4126 ( .A1(MEM_stage_inst_dmem_n3982), .A2(MEM_stage_inst_dmem_n3981), .ZN(MEM_stage_inst_dmem_n3983) );
NAND2_X1 MEM_stage_inst_dmem_U4125 ( .A1(MEM_stage_inst_dmem_n3980), .A2(MEM_stage_inst_dmem_n3979), .ZN(MEM_stage_inst_dmem_n3981) );
NAND2_X1 MEM_stage_inst_dmem_U4124 ( .A1(MEM_stage_inst_dmem_ram_3127), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n3979) );
NAND2_X1 MEM_stage_inst_dmem_U4123 ( .A1(MEM_stage_inst_dmem_ram_3767), .A2(MEM_stage_inst_dmem_n4709), .ZN(MEM_stage_inst_dmem_n3980) );
NAND2_X1 MEM_stage_inst_dmem_U4122 ( .A1(MEM_stage_inst_dmem_n3978), .A2(MEM_stage_inst_dmem_n3977), .ZN(MEM_stage_inst_dmem_n3982) );
NAND2_X1 MEM_stage_inst_dmem_U4121 ( .A1(MEM_stage_inst_dmem_ram_3959), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n3977) );
NAND2_X1 MEM_stage_inst_dmem_U4120 ( .A1(MEM_stage_inst_dmem_ram_4055), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n3978) );
NOR2_X1 MEM_stage_inst_dmem_U4119 ( .A1(MEM_stage_inst_dmem_n3976), .A2(MEM_stage_inst_dmem_n3975), .ZN(MEM_stage_inst_dmem_n3984) );
NAND2_X1 MEM_stage_inst_dmem_U4118 ( .A1(MEM_stage_inst_dmem_n3974), .A2(MEM_stage_inst_dmem_n3973), .ZN(MEM_stage_inst_dmem_n3975) );
NAND2_X1 MEM_stage_inst_dmem_U4117 ( .A1(MEM_stage_inst_dmem_ram_3479), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n3973) );
NAND2_X1 MEM_stage_inst_dmem_U4116 ( .A1(MEM_stage_inst_dmem_ram_3335), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n3974) );
NAND2_X1 MEM_stage_inst_dmem_U4115 ( .A1(MEM_stage_inst_dmem_n3972), .A2(MEM_stage_inst_dmem_n3971), .ZN(MEM_stage_inst_dmem_n3976) );
NAND2_X1 MEM_stage_inst_dmem_U4114 ( .A1(MEM_stage_inst_dmem_ram_3303), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n3971) );
NAND2_X1 MEM_stage_inst_dmem_U4113 ( .A1(MEM_stage_inst_dmem_ram_3559), .A2(MEM_stage_inst_dmem_n4667), .ZN(MEM_stage_inst_dmem_n3972) );
NOR2_X1 MEM_stage_inst_dmem_U4112 ( .A1(MEM_stage_inst_dmem_n3970), .A2(MEM_stage_inst_dmem_n3969), .ZN(MEM_stage_inst_dmem_n4002) );
NAND2_X1 MEM_stage_inst_dmem_U4111 ( .A1(MEM_stage_inst_dmem_n3968), .A2(MEM_stage_inst_dmem_n3967), .ZN(MEM_stage_inst_dmem_n3969) );
NOR2_X1 MEM_stage_inst_dmem_U4110 ( .A1(MEM_stage_inst_dmem_n3966), .A2(MEM_stage_inst_dmem_n3965), .ZN(MEM_stage_inst_dmem_n3967) );
NAND2_X1 MEM_stage_inst_dmem_U4109 ( .A1(MEM_stage_inst_dmem_n3964), .A2(MEM_stage_inst_dmem_n3963), .ZN(MEM_stage_inst_dmem_n3965) );
NAND2_X1 MEM_stage_inst_dmem_U4108 ( .A1(MEM_stage_inst_dmem_ram_3895), .A2(MEM_stage_inst_dmem_n4740), .ZN(MEM_stage_inst_dmem_n3963) );
NAND2_X1 MEM_stage_inst_dmem_U4107 ( .A1(MEM_stage_inst_dmem_ram_3223), .A2(MEM_stage_inst_dmem_n5807), .ZN(MEM_stage_inst_dmem_n3964) );
NAND2_X1 MEM_stage_inst_dmem_U4106 ( .A1(MEM_stage_inst_dmem_n3962), .A2(MEM_stage_inst_dmem_n3961), .ZN(MEM_stage_inst_dmem_n3966) );
NAND2_X1 MEM_stage_inst_dmem_U4105 ( .A1(MEM_stage_inst_dmem_ram_3927), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n3961) );
NAND2_X1 MEM_stage_inst_dmem_U4104 ( .A1(MEM_stage_inst_dmem_ram_3911), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n3962) );
NOR2_X1 MEM_stage_inst_dmem_U4103 ( .A1(MEM_stage_inst_dmem_n3960), .A2(MEM_stage_inst_dmem_n3959), .ZN(MEM_stage_inst_dmem_n3968) );
NAND2_X1 MEM_stage_inst_dmem_U4102 ( .A1(MEM_stage_inst_dmem_n3958), .A2(MEM_stage_inst_dmem_n3957), .ZN(MEM_stage_inst_dmem_n3959) );
NAND2_X1 MEM_stage_inst_dmem_U4101 ( .A1(MEM_stage_inst_dmem_ram_3991), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n3957) );
NAND2_X1 MEM_stage_inst_dmem_U4100 ( .A1(MEM_stage_inst_dmem_ram_3751), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n3958) );
NAND2_X1 MEM_stage_inst_dmem_U4099 ( .A1(MEM_stage_inst_dmem_n3956), .A2(MEM_stage_inst_dmem_n3955), .ZN(MEM_stage_inst_dmem_n3960) );
NAND2_X1 MEM_stage_inst_dmem_U4098 ( .A1(MEM_stage_inst_dmem_ram_4087), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n3955) );
NAND2_X1 MEM_stage_inst_dmem_U4097 ( .A1(MEM_stage_inst_dmem_ram_3735), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n3956) );
NAND2_X1 MEM_stage_inst_dmem_U4096 ( .A1(MEM_stage_inst_dmem_n3954), .A2(MEM_stage_inst_dmem_n3953), .ZN(MEM_stage_inst_dmem_n3970) );
NOR2_X1 MEM_stage_inst_dmem_U4095 ( .A1(MEM_stage_inst_dmem_n3952), .A2(MEM_stage_inst_dmem_n3951), .ZN(MEM_stage_inst_dmem_n3953) );
NAND2_X1 MEM_stage_inst_dmem_U4094 ( .A1(MEM_stage_inst_dmem_n3950), .A2(MEM_stage_inst_dmem_n3949), .ZN(MEM_stage_inst_dmem_n3951) );
NAND2_X1 MEM_stage_inst_dmem_U4093 ( .A1(MEM_stage_inst_dmem_ram_3399), .A2(MEM_stage_inst_dmem_n4706), .ZN(MEM_stage_inst_dmem_n3949) );
NAND2_X1 MEM_stage_inst_dmem_U4092 ( .A1(MEM_stage_inst_dmem_ram_3975), .A2(MEM_stage_inst_dmem_n72), .ZN(MEM_stage_inst_dmem_n3950) );
NAND2_X1 MEM_stage_inst_dmem_U4091 ( .A1(MEM_stage_inst_dmem_n3948), .A2(MEM_stage_inst_dmem_n3947), .ZN(MEM_stage_inst_dmem_n3952) );
NAND2_X1 MEM_stage_inst_dmem_U4090 ( .A1(MEM_stage_inst_dmem_ram_3575), .A2(MEM_stage_inst_dmem_n64), .ZN(MEM_stage_inst_dmem_n3947) );
NAND2_X1 MEM_stage_inst_dmem_U4089 ( .A1(MEM_stage_inst_dmem_ram_3591), .A2(MEM_stage_inst_dmem_n71), .ZN(MEM_stage_inst_dmem_n3948) );
NOR2_X1 MEM_stage_inst_dmem_U4088 ( .A1(MEM_stage_inst_dmem_n3946), .A2(MEM_stage_inst_dmem_n3945), .ZN(MEM_stage_inst_dmem_n3954) );
NAND2_X1 MEM_stage_inst_dmem_U4087 ( .A1(MEM_stage_inst_dmem_n3944), .A2(MEM_stage_inst_dmem_n3943), .ZN(MEM_stage_inst_dmem_n3945) );
NAND2_X1 MEM_stage_inst_dmem_U4086 ( .A1(MEM_stage_inst_dmem_ram_3639), .A2(MEM_stage_inst_dmem_n41), .ZN(MEM_stage_inst_dmem_n3943) );
NAND2_X1 MEM_stage_inst_dmem_U4085 ( .A1(MEM_stage_inst_dmem_ram_3527), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n3944) );
NAND2_X1 MEM_stage_inst_dmem_U4084 ( .A1(MEM_stage_inst_dmem_n3942), .A2(MEM_stage_inst_dmem_n3941), .ZN(MEM_stage_inst_dmem_n3946) );
NAND2_X1 MEM_stage_inst_dmem_U4083 ( .A1(MEM_stage_inst_dmem_ram_3943), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n3941) );
NAND2_X1 MEM_stage_inst_dmem_U4082 ( .A1(MEM_stage_inst_dmem_ram_3671), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n3942) );
NAND2_X1 MEM_stage_inst_dmem_U4081 ( .A1(MEM_stage_inst_dmem_n3940), .A2(MEM_stage_inst_dmem_n3939), .ZN(MEM_stage_inst_dmem_n4004) );
NOR2_X1 MEM_stage_inst_dmem_U4080 ( .A1(MEM_stage_inst_dmem_n3938), .A2(MEM_stage_inst_dmem_n3937), .ZN(MEM_stage_inst_dmem_n3939) );
NAND2_X1 MEM_stage_inst_dmem_U4079 ( .A1(MEM_stage_inst_dmem_n3936), .A2(MEM_stage_inst_dmem_n3935), .ZN(MEM_stage_inst_dmem_n3937) );
NOR2_X1 MEM_stage_inst_dmem_U4078 ( .A1(MEM_stage_inst_dmem_n3934), .A2(MEM_stage_inst_dmem_n3933), .ZN(MEM_stage_inst_dmem_n3935) );
NAND2_X1 MEM_stage_inst_dmem_U4077 ( .A1(MEM_stage_inst_dmem_n3932), .A2(MEM_stage_inst_dmem_n3931), .ZN(MEM_stage_inst_dmem_n3933) );
NAND2_X1 MEM_stage_inst_dmem_U4076 ( .A1(MEM_stage_inst_dmem_ram_3191), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n3931) );
NAND2_X1 MEM_stage_inst_dmem_U4075 ( .A1(MEM_stage_inst_dmem_ram_3687), .A2(MEM_stage_inst_dmem_n4701), .ZN(MEM_stage_inst_dmem_n3932) );
NAND2_X1 MEM_stage_inst_dmem_U4074 ( .A1(MEM_stage_inst_dmem_n3930), .A2(MEM_stage_inst_dmem_n3929), .ZN(MEM_stage_inst_dmem_n3934) );
NAND2_X1 MEM_stage_inst_dmem_U4073 ( .A1(MEM_stage_inst_dmem_ram_3511), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n3929) );
NAND2_X1 MEM_stage_inst_dmem_U4072 ( .A1(MEM_stage_inst_dmem_ram_3319), .A2(MEM_stage_inst_dmem_n4649), .ZN(MEM_stage_inst_dmem_n3930) );
NOR2_X1 MEM_stage_inst_dmem_U4071 ( .A1(MEM_stage_inst_dmem_n3928), .A2(MEM_stage_inst_dmem_n3927), .ZN(MEM_stage_inst_dmem_n3936) );
NAND2_X1 MEM_stage_inst_dmem_U4070 ( .A1(MEM_stage_inst_dmem_n3926), .A2(MEM_stage_inst_dmem_n3925), .ZN(MEM_stage_inst_dmem_n3927) );
NAND2_X1 MEM_stage_inst_dmem_U4069 ( .A1(MEM_stage_inst_dmem_ram_3095), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n3925) );
NAND2_X1 MEM_stage_inst_dmem_U4068 ( .A1(MEM_stage_inst_dmem_ram_3287), .A2(MEM_stage_inst_dmem_n51), .ZN(MEM_stage_inst_dmem_n3926) );
NAND2_X1 MEM_stage_inst_dmem_U4067 ( .A1(MEM_stage_inst_dmem_n3924), .A2(MEM_stage_inst_dmem_n3923), .ZN(MEM_stage_inst_dmem_n3928) );
NAND2_X1 MEM_stage_inst_dmem_U4066 ( .A1(MEM_stage_inst_dmem_ram_3623), .A2(MEM_stage_inst_dmem_n4692), .ZN(MEM_stage_inst_dmem_n3923) );
NAND2_X1 MEM_stage_inst_dmem_U4065 ( .A1(MEM_stage_inst_dmem_ram_4007), .A2(MEM_stage_inst_dmem_n4675), .ZN(MEM_stage_inst_dmem_n3924) );
NAND2_X1 MEM_stage_inst_dmem_U4064 ( .A1(MEM_stage_inst_dmem_n3922), .A2(MEM_stage_inst_dmem_n3921), .ZN(MEM_stage_inst_dmem_n3938) );
NOR2_X1 MEM_stage_inst_dmem_U4063 ( .A1(MEM_stage_inst_dmem_n3920), .A2(MEM_stage_inst_dmem_n3919), .ZN(MEM_stage_inst_dmem_n3921) );
NAND2_X1 MEM_stage_inst_dmem_U4062 ( .A1(MEM_stage_inst_dmem_n3918), .A2(MEM_stage_inst_dmem_n3917), .ZN(MEM_stage_inst_dmem_n3919) );
NAND2_X1 MEM_stage_inst_dmem_U4061 ( .A1(MEM_stage_inst_dmem_ram_3431), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n3917) );
NAND2_X1 MEM_stage_inst_dmem_U4060 ( .A1(MEM_stage_inst_dmem_ram_3655), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n3918) );
NAND2_X1 MEM_stage_inst_dmem_U4059 ( .A1(MEM_stage_inst_dmem_n3916), .A2(MEM_stage_inst_dmem_n3915), .ZN(MEM_stage_inst_dmem_n3920) );
NAND2_X1 MEM_stage_inst_dmem_U4058 ( .A1(MEM_stage_inst_dmem_ram_3719), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n3915) );
NAND2_X1 MEM_stage_inst_dmem_U4057 ( .A1(MEM_stage_inst_dmem_ram_3255), .A2(MEM_stage_inst_dmem_n55), .ZN(MEM_stage_inst_dmem_n3916) );
NOR2_X1 MEM_stage_inst_dmem_U4056 ( .A1(MEM_stage_inst_dmem_n3914), .A2(MEM_stage_inst_dmem_n3913), .ZN(MEM_stage_inst_dmem_n3922) );
NAND2_X1 MEM_stage_inst_dmem_U4055 ( .A1(MEM_stage_inst_dmem_n3912), .A2(MEM_stage_inst_dmem_n3911), .ZN(MEM_stage_inst_dmem_n3913) );
NAND2_X1 MEM_stage_inst_dmem_U4054 ( .A1(MEM_stage_inst_dmem_ram_3271), .A2(MEM_stage_inst_dmem_n36), .ZN(MEM_stage_inst_dmem_n3911) );
NAND2_X1 MEM_stage_inst_dmem_U4053 ( .A1(MEM_stage_inst_dmem_ram_3703), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n3912) );
NAND2_X1 MEM_stage_inst_dmem_U4052 ( .A1(MEM_stage_inst_dmem_n3910), .A2(MEM_stage_inst_dmem_n3909), .ZN(MEM_stage_inst_dmem_n3914) );
NAND2_X1 MEM_stage_inst_dmem_U4051 ( .A1(MEM_stage_inst_dmem_ram_3143), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n3909) );
NAND2_X1 MEM_stage_inst_dmem_U4050 ( .A1(MEM_stage_inst_dmem_ram_3175), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n3910) );
NOR2_X1 MEM_stage_inst_dmem_U4049 ( .A1(MEM_stage_inst_dmem_n3908), .A2(MEM_stage_inst_dmem_n3907), .ZN(MEM_stage_inst_dmem_n3940) );
NAND2_X1 MEM_stage_inst_dmem_U4048 ( .A1(MEM_stage_inst_dmem_n3906), .A2(MEM_stage_inst_dmem_n3905), .ZN(MEM_stage_inst_dmem_n3907) );
NOR2_X1 MEM_stage_inst_dmem_U4047 ( .A1(MEM_stage_inst_dmem_n3904), .A2(MEM_stage_inst_dmem_n3903), .ZN(MEM_stage_inst_dmem_n3905) );
NAND2_X1 MEM_stage_inst_dmem_U4046 ( .A1(MEM_stage_inst_dmem_n3902), .A2(MEM_stage_inst_dmem_n3901), .ZN(MEM_stage_inst_dmem_n3903) );
NAND2_X1 MEM_stage_inst_dmem_U4045 ( .A1(MEM_stage_inst_dmem_ram_3847), .A2(MEM_stage_inst_dmem_n37), .ZN(MEM_stage_inst_dmem_n3901) );
NAND2_X1 MEM_stage_inst_dmem_U4044 ( .A1(MEM_stage_inst_dmem_ram_3415), .A2(MEM_stage_inst_dmem_n3216), .ZN(MEM_stage_inst_dmem_n3902) );
NAND2_X1 MEM_stage_inst_dmem_U4043 ( .A1(MEM_stage_inst_dmem_n3900), .A2(MEM_stage_inst_dmem_n3899), .ZN(MEM_stage_inst_dmem_n3904) );
NAND2_X1 MEM_stage_inst_dmem_U4042 ( .A1(MEM_stage_inst_dmem_ram_3239), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n3899) );
NAND2_X1 MEM_stage_inst_dmem_U4041 ( .A1(MEM_stage_inst_dmem_ram_3815), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n3900) );
NOR2_X1 MEM_stage_inst_dmem_U4040 ( .A1(MEM_stage_inst_dmem_n3898), .A2(MEM_stage_inst_dmem_n3897), .ZN(MEM_stage_inst_dmem_n3906) );
NAND2_X1 MEM_stage_inst_dmem_U4039 ( .A1(MEM_stage_inst_dmem_n3896), .A2(MEM_stage_inst_dmem_n3895), .ZN(MEM_stage_inst_dmem_n3897) );
NAND2_X1 MEM_stage_inst_dmem_U4038 ( .A1(MEM_stage_inst_dmem_ram_3831), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n3895) );
NAND2_X1 MEM_stage_inst_dmem_U4037 ( .A1(MEM_stage_inst_dmem_ram_3863), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n3896) );
NAND2_X1 MEM_stage_inst_dmem_U4036 ( .A1(MEM_stage_inst_dmem_n3894), .A2(MEM_stage_inst_dmem_n3893), .ZN(MEM_stage_inst_dmem_n3898) );
NAND2_X1 MEM_stage_inst_dmem_U4035 ( .A1(MEM_stage_inst_dmem_ram_3495), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n3893) );
NAND2_X1 MEM_stage_inst_dmem_U4034 ( .A1(MEM_stage_inst_dmem_ram_3111), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n3894) );
NAND2_X1 MEM_stage_inst_dmem_U4033 ( .A1(MEM_stage_inst_dmem_n3892), .A2(MEM_stage_inst_dmem_n3891), .ZN(MEM_stage_inst_dmem_n3908) );
NOR2_X1 MEM_stage_inst_dmem_U4032 ( .A1(MEM_stage_inst_dmem_n3890), .A2(MEM_stage_inst_dmem_n3889), .ZN(MEM_stage_inst_dmem_n3891) );
NAND2_X1 MEM_stage_inst_dmem_U4031 ( .A1(MEM_stage_inst_dmem_n3888), .A2(MEM_stage_inst_dmem_n3887), .ZN(MEM_stage_inst_dmem_n3889) );
NAND2_X1 MEM_stage_inst_dmem_U4030 ( .A1(MEM_stage_inst_dmem_ram_4023), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n3887) );
NAND2_X1 MEM_stage_inst_dmem_U4029 ( .A1(MEM_stage_inst_dmem_ram_3207), .A2(MEM_stage_inst_dmem_n61), .ZN(MEM_stage_inst_dmem_n3888) );
NAND2_X1 MEM_stage_inst_dmem_U4028 ( .A1(MEM_stage_inst_dmem_n3886), .A2(MEM_stage_inst_dmem_n3885), .ZN(MEM_stage_inst_dmem_n3890) );
NAND2_X1 MEM_stage_inst_dmem_U4027 ( .A1(MEM_stage_inst_dmem_ram_3383), .A2(MEM_stage_inst_dmem_n4731), .ZN(MEM_stage_inst_dmem_n3885) );
NAND2_X1 MEM_stage_inst_dmem_U4026 ( .A1(MEM_stage_inst_dmem_ram_3607), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n3886) );
NOR2_X1 MEM_stage_inst_dmem_U4025 ( .A1(MEM_stage_inst_dmem_n3884), .A2(MEM_stage_inst_dmem_n3883), .ZN(MEM_stage_inst_dmem_n3892) );
NAND2_X1 MEM_stage_inst_dmem_U4024 ( .A1(MEM_stage_inst_dmem_n3882), .A2(MEM_stage_inst_dmem_n3881), .ZN(MEM_stage_inst_dmem_n3883) );
NAND2_X1 MEM_stage_inst_dmem_U4023 ( .A1(MEM_stage_inst_dmem_ram_4039), .A2(MEM_stage_inst_dmem_n4728), .ZN(MEM_stage_inst_dmem_n3881) );
NAND2_X1 MEM_stage_inst_dmem_U4022 ( .A1(MEM_stage_inst_dmem_ram_3799), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n3882) );
NAND2_X1 MEM_stage_inst_dmem_U4021 ( .A1(MEM_stage_inst_dmem_n3880), .A2(MEM_stage_inst_dmem_n3879), .ZN(MEM_stage_inst_dmem_n3884) );
NAND2_X1 MEM_stage_inst_dmem_U4020 ( .A1(MEM_stage_inst_dmem_ram_3783), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n3879) );
NAND2_X1 MEM_stage_inst_dmem_U4019 ( .A1(MEM_stage_inst_dmem_ram_3447), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n3880) );
NAND2_X1 MEM_stage_inst_dmem_U4018 ( .A1(MEM_stage_inst_dmem_n3878), .A2(MEM_stage_inst_dmem_n3877), .ZN(MEM_stage_inst_mem_read_data_6) );
NOR2_X1 MEM_stage_inst_dmem_U4017 ( .A1(MEM_stage_inst_dmem_n3876), .A2(MEM_stage_inst_dmem_n3875), .ZN(MEM_stage_inst_dmem_n3877) );
NOR2_X1 MEM_stage_inst_dmem_U4016 ( .A1(MEM_stage_inst_dmem_n3874), .A2(MEM_stage_inst_dmem_n8551), .ZN(MEM_stage_inst_dmem_n3875) );
NOR2_X1 MEM_stage_inst_dmem_U4015 ( .A1(MEM_stage_inst_dmem_n3873), .A2(MEM_stage_inst_dmem_n3872), .ZN(MEM_stage_inst_dmem_n3874) );
NAND2_X1 MEM_stage_inst_dmem_U4014 ( .A1(MEM_stage_inst_dmem_n3871), .A2(MEM_stage_inst_dmem_n3870), .ZN(MEM_stage_inst_dmem_n3872) );
NOR2_X1 MEM_stage_inst_dmem_U4013 ( .A1(MEM_stage_inst_dmem_n3869), .A2(MEM_stage_inst_dmem_n3868), .ZN(MEM_stage_inst_dmem_n3870) );
NAND2_X1 MEM_stage_inst_dmem_U4012 ( .A1(MEM_stage_inst_dmem_n3867), .A2(MEM_stage_inst_dmem_n3866), .ZN(MEM_stage_inst_dmem_n3868) );
NOR2_X1 MEM_stage_inst_dmem_U4011 ( .A1(MEM_stage_inst_dmem_n3865), .A2(MEM_stage_inst_dmem_n3864), .ZN(MEM_stage_inst_dmem_n3866) );
NAND2_X1 MEM_stage_inst_dmem_U4010 ( .A1(MEM_stage_inst_dmem_n3863), .A2(MEM_stage_inst_dmem_n3862), .ZN(MEM_stage_inst_dmem_n3864) );
NAND2_X1 MEM_stage_inst_dmem_U4009 ( .A1(MEM_stage_inst_dmem_ram_566), .A2(MEM_stage_inst_dmem_n41), .ZN(MEM_stage_inst_dmem_n3862) );
NAND2_X1 MEM_stage_inst_dmem_U4008 ( .A1(MEM_stage_inst_dmem_ram_486), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n3863) );
NAND2_X1 MEM_stage_inst_dmem_U4007 ( .A1(MEM_stage_inst_dmem_n3861), .A2(MEM_stage_inst_dmem_n3860), .ZN(MEM_stage_inst_dmem_n3865) );
NAND2_X1 MEM_stage_inst_dmem_U4006 ( .A1(MEM_stage_inst_dmem_ram_918), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n3860) );
NAND2_X1 MEM_stage_inst_dmem_U4005 ( .A1(MEM_stage_inst_dmem_ram_614), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n3861) );
NOR2_X1 MEM_stage_inst_dmem_U4004 ( .A1(MEM_stage_inst_dmem_n3859), .A2(MEM_stage_inst_dmem_n3858), .ZN(MEM_stage_inst_dmem_n3867) );
NAND2_X1 MEM_stage_inst_dmem_U4003 ( .A1(MEM_stage_inst_dmem_n3857), .A2(MEM_stage_inst_dmem_n3856), .ZN(MEM_stage_inst_dmem_n3858) );
NAND2_X1 MEM_stage_inst_dmem_U4002 ( .A1(MEM_stage_inst_dmem_ram_726), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n3856) );
NAND2_X1 MEM_stage_inst_dmem_U4001 ( .A1(MEM_stage_inst_dmem_ram_742), .A2(MEM_stage_inst_dmem_n4769), .ZN(MEM_stage_inst_dmem_n3857) );
NAND2_X1 MEM_stage_inst_dmem_U4000 ( .A1(MEM_stage_inst_dmem_n3855), .A2(MEM_stage_inst_dmem_n3854), .ZN(MEM_stage_inst_dmem_n3859) );
NAND2_X1 MEM_stage_inst_dmem_U3999 ( .A1(MEM_stage_inst_dmem_ram_822), .A2(MEM_stage_inst_dmem_n46), .ZN(MEM_stage_inst_dmem_n3854) );
NAND2_X1 MEM_stage_inst_dmem_U3998 ( .A1(MEM_stage_inst_dmem_ram_790), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n3855) );
NAND2_X1 MEM_stage_inst_dmem_U3997 ( .A1(MEM_stage_inst_dmem_n3853), .A2(MEM_stage_inst_dmem_n3852), .ZN(MEM_stage_inst_dmem_n3869) );
NOR2_X1 MEM_stage_inst_dmem_U3996 ( .A1(MEM_stage_inst_dmem_n3851), .A2(MEM_stage_inst_dmem_n3850), .ZN(MEM_stage_inst_dmem_n3852) );
NAND2_X1 MEM_stage_inst_dmem_U3995 ( .A1(MEM_stage_inst_dmem_n3849), .A2(MEM_stage_inst_dmem_n3848), .ZN(MEM_stage_inst_dmem_n3850) );
NAND2_X1 MEM_stage_inst_dmem_U3994 ( .A1(MEM_stage_inst_dmem_ram_246), .A2(MEM_stage_inst_dmem_n39), .ZN(MEM_stage_inst_dmem_n3848) );
NAND2_X1 MEM_stage_inst_dmem_U3993 ( .A1(MEM_stage_inst_dmem_ram_982), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n3849) );
NAND2_X1 MEM_stage_inst_dmem_U3992 ( .A1(MEM_stage_inst_dmem_n3847), .A2(MEM_stage_inst_dmem_n3846), .ZN(MEM_stage_inst_dmem_n3851) );
NAND2_X1 MEM_stage_inst_dmem_U3991 ( .A1(MEM_stage_inst_dmem_ram_950), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n3846) );
NAND2_X1 MEM_stage_inst_dmem_U3990 ( .A1(MEM_stage_inst_dmem_ram_454), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n3847) );
NOR2_X1 MEM_stage_inst_dmem_U3989 ( .A1(MEM_stage_inst_dmem_n3845), .A2(MEM_stage_inst_dmem_n3844), .ZN(MEM_stage_inst_dmem_n3853) );
NAND2_X1 MEM_stage_inst_dmem_U3988 ( .A1(MEM_stage_inst_dmem_n3843), .A2(MEM_stage_inst_dmem_n3842), .ZN(MEM_stage_inst_dmem_n3844) );
NAND2_X1 MEM_stage_inst_dmem_U3987 ( .A1(MEM_stage_inst_dmem_ram_310), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n3842) );
NAND2_X1 MEM_stage_inst_dmem_U3986 ( .A1(MEM_stage_inst_dmem_ram_678), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n3843) );
NAND2_X1 MEM_stage_inst_dmem_U3985 ( .A1(MEM_stage_inst_dmem_n3841), .A2(MEM_stage_inst_dmem_n3840), .ZN(MEM_stage_inst_dmem_n3845) );
NAND2_X1 MEM_stage_inst_dmem_U3984 ( .A1(MEM_stage_inst_dmem_ram_326), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n3840) );
NAND2_X1 MEM_stage_inst_dmem_U3983 ( .A1(MEM_stage_inst_dmem_ram_934), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n3841) );
NOR2_X1 MEM_stage_inst_dmem_U3982 ( .A1(MEM_stage_inst_dmem_n3839), .A2(MEM_stage_inst_dmem_n3838), .ZN(MEM_stage_inst_dmem_n3871) );
NAND2_X1 MEM_stage_inst_dmem_U3981 ( .A1(MEM_stage_inst_dmem_n3837), .A2(MEM_stage_inst_dmem_n3836), .ZN(MEM_stage_inst_dmem_n3838) );
NOR2_X1 MEM_stage_inst_dmem_U3980 ( .A1(MEM_stage_inst_dmem_n3835), .A2(MEM_stage_inst_dmem_n3834), .ZN(MEM_stage_inst_dmem_n3836) );
NAND2_X1 MEM_stage_inst_dmem_U3979 ( .A1(MEM_stage_inst_dmem_n3833), .A2(MEM_stage_inst_dmem_n3832), .ZN(MEM_stage_inst_dmem_n3834) );
NAND2_X1 MEM_stage_inst_dmem_U3978 ( .A1(MEM_stage_inst_dmem_ram_86), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n3832) );
NAND2_X1 MEM_stage_inst_dmem_U3977 ( .A1(MEM_stage_inst_dmem_ram_102), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n3833) );
NAND2_X1 MEM_stage_inst_dmem_U3976 ( .A1(MEM_stage_inst_dmem_n3831), .A2(MEM_stage_inst_dmem_n3830), .ZN(MEM_stage_inst_dmem_n3835) );
NAND2_X1 MEM_stage_inst_dmem_U3975 ( .A1(MEM_stage_inst_dmem_ram_230), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n3830) );
NAND2_X1 MEM_stage_inst_dmem_U3974 ( .A1(MEM_stage_inst_dmem_ram_470), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n3831) );
NOR2_X1 MEM_stage_inst_dmem_U3973 ( .A1(MEM_stage_inst_dmem_n3829), .A2(MEM_stage_inst_dmem_n3828), .ZN(MEM_stage_inst_dmem_n3837) );
NAND2_X1 MEM_stage_inst_dmem_U3972 ( .A1(MEM_stage_inst_dmem_n3827), .A2(MEM_stage_inst_dmem_n3826), .ZN(MEM_stage_inst_dmem_n3828) );
NAND2_X1 MEM_stage_inst_dmem_U3971 ( .A1(MEM_stage_inst_dmem_ram_598), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n3826) );
NAND2_X1 MEM_stage_inst_dmem_U3970 ( .A1(MEM_stage_inst_dmem_ram_6), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n3827) );
NAND2_X1 MEM_stage_inst_dmem_U3969 ( .A1(MEM_stage_inst_dmem_n3825), .A2(MEM_stage_inst_dmem_n3824), .ZN(MEM_stage_inst_dmem_n3829) );
NAND2_X1 MEM_stage_inst_dmem_U3968 ( .A1(MEM_stage_inst_dmem_ram_406), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n3824) );
NAND2_X1 MEM_stage_inst_dmem_U3967 ( .A1(MEM_stage_inst_dmem_ram_38), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n3825) );
NAND2_X1 MEM_stage_inst_dmem_U3966 ( .A1(MEM_stage_inst_dmem_n3823), .A2(MEM_stage_inst_dmem_n3822), .ZN(MEM_stage_inst_dmem_n3839) );
NOR2_X1 MEM_stage_inst_dmem_U3965 ( .A1(MEM_stage_inst_dmem_n3821), .A2(MEM_stage_inst_dmem_n3820), .ZN(MEM_stage_inst_dmem_n3822) );
NAND2_X1 MEM_stage_inst_dmem_U3964 ( .A1(MEM_stage_inst_dmem_n3819), .A2(MEM_stage_inst_dmem_n3818), .ZN(MEM_stage_inst_dmem_n3820) );
NAND2_X1 MEM_stage_inst_dmem_U3963 ( .A1(MEM_stage_inst_dmem_ram_214), .A2(MEM_stage_inst_dmem_n51), .ZN(MEM_stage_inst_dmem_n3818) );
NAND2_X1 MEM_stage_inst_dmem_U3962 ( .A1(MEM_stage_inst_dmem_ram_1014), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n3819) );
NAND2_X1 MEM_stage_inst_dmem_U3961 ( .A1(MEM_stage_inst_dmem_n3817), .A2(MEM_stage_inst_dmem_n3816), .ZN(MEM_stage_inst_dmem_n3821) );
NAND2_X1 MEM_stage_inst_dmem_U3960 ( .A1(MEM_stage_inst_dmem_ram_70), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n3816) );
NAND2_X1 MEM_stage_inst_dmem_U3959 ( .A1(MEM_stage_inst_dmem_ram_278), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n3817) );
NOR2_X1 MEM_stage_inst_dmem_U3958 ( .A1(MEM_stage_inst_dmem_n3815), .A2(MEM_stage_inst_dmem_n3814), .ZN(MEM_stage_inst_dmem_n3823) );
NAND2_X1 MEM_stage_inst_dmem_U3957 ( .A1(MEM_stage_inst_dmem_n3813), .A2(MEM_stage_inst_dmem_n3812), .ZN(MEM_stage_inst_dmem_n3814) );
NAND2_X1 MEM_stage_inst_dmem_U3956 ( .A1(MEM_stage_inst_dmem_ram_294), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n3812) );
NAND2_X1 MEM_stage_inst_dmem_U3955 ( .A1(MEM_stage_inst_dmem_ram_518), .A2(MEM_stage_inst_dmem_n71), .ZN(MEM_stage_inst_dmem_n3813) );
NAND2_X1 MEM_stage_inst_dmem_U3954 ( .A1(MEM_stage_inst_dmem_n3811), .A2(MEM_stage_inst_dmem_n3810), .ZN(MEM_stage_inst_dmem_n3815) );
NAND2_X1 MEM_stage_inst_dmem_U3953 ( .A1(MEM_stage_inst_dmem_ram_998), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n3810) );
NAND2_X1 MEM_stage_inst_dmem_U3952 ( .A1(MEM_stage_inst_dmem_ram_422), .A2(MEM_stage_inst_dmem_n4772), .ZN(MEM_stage_inst_dmem_n3811) );
NAND2_X1 MEM_stage_inst_dmem_U3951 ( .A1(MEM_stage_inst_dmem_n3809), .A2(MEM_stage_inst_dmem_n3808), .ZN(MEM_stage_inst_dmem_n3873) );
NOR2_X1 MEM_stage_inst_dmem_U3950 ( .A1(MEM_stage_inst_dmem_n3807), .A2(MEM_stage_inst_dmem_n3806), .ZN(MEM_stage_inst_dmem_n3808) );
NAND2_X1 MEM_stage_inst_dmem_U3949 ( .A1(MEM_stage_inst_dmem_n3805), .A2(MEM_stage_inst_dmem_n3804), .ZN(MEM_stage_inst_dmem_n3806) );
NOR2_X1 MEM_stage_inst_dmem_U3948 ( .A1(MEM_stage_inst_dmem_n3803), .A2(MEM_stage_inst_dmem_n3802), .ZN(MEM_stage_inst_dmem_n3804) );
NAND2_X1 MEM_stage_inst_dmem_U3947 ( .A1(MEM_stage_inst_dmem_n3801), .A2(MEM_stage_inst_dmem_n3800), .ZN(MEM_stage_inst_dmem_n3802) );
NAND2_X1 MEM_stage_inst_dmem_U3946 ( .A1(MEM_stage_inst_dmem_ram_134), .A2(MEM_stage_inst_dmem_n61), .ZN(MEM_stage_inst_dmem_n3800) );
NAND2_X1 MEM_stage_inst_dmem_U3945 ( .A1(MEM_stage_inst_dmem_ram_550), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n3801) );
NAND2_X1 MEM_stage_inst_dmem_U3944 ( .A1(MEM_stage_inst_dmem_n3799), .A2(MEM_stage_inst_dmem_n3798), .ZN(MEM_stage_inst_dmem_n3803) );
NAND2_X1 MEM_stage_inst_dmem_U3943 ( .A1(MEM_stage_inst_dmem_ram_438), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n3798) );
NAND2_X1 MEM_stage_inst_dmem_U3942 ( .A1(MEM_stage_inst_dmem_ram_150), .A2(MEM_stage_inst_dmem_n5807), .ZN(MEM_stage_inst_dmem_n3799) );
NOR2_X1 MEM_stage_inst_dmem_U3941 ( .A1(MEM_stage_inst_dmem_n3797), .A2(MEM_stage_inst_dmem_n3796), .ZN(MEM_stage_inst_dmem_n3805) );
NAND2_X1 MEM_stage_inst_dmem_U3940 ( .A1(MEM_stage_inst_dmem_n3795), .A2(MEM_stage_inst_dmem_n3794), .ZN(MEM_stage_inst_dmem_n3796) );
NAND2_X1 MEM_stage_inst_dmem_U3939 ( .A1(MEM_stage_inst_dmem_ram_870), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n3794) );
NAND2_X1 MEM_stage_inst_dmem_U3938 ( .A1(MEM_stage_inst_dmem_ram_534), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n3795) );
NAND2_X1 MEM_stage_inst_dmem_U3937 ( .A1(MEM_stage_inst_dmem_n3793), .A2(MEM_stage_inst_dmem_n3792), .ZN(MEM_stage_inst_dmem_n3797) );
NAND2_X1 MEM_stage_inst_dmem_U3936 ( .A1(MEM_stage_inst_dmem_ram_886), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n3792) );
NAND2_X1 MEM_stage_inst_dmem_U3935 ( .A1(MEM_stage_inst_dmem_ram_646), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n3793) );
NAND2_X1 MEM_stage_inst_dmem_U3934 ( .A1(MEM_stage_inst_dmem_n3791), .A2(MEM_stage_inst_dmem_n3790), .ZN(MEM_stage_inst_dmem_n3807) );
NOR2_X1 MEM_stage_inst_dmem_U3933 ( .A1(MEM_stage_inst_dmem_n3789), .A2(MEM_stage_inst_dmem_n3788), .ZN(MEM_stage_inst_dmem_n3790) );
NAND2_X1 MEM_stage_inst_dmem_U3932 ( .A1(MEM_stage_inst_dmem_n3787), .A2(MEM_stage_inst_dmem_n3786), .ZN(MEM_stage_inst_dmem_n3788) );
NAND2_X1 MEM_stage_inst_dmem_U3931 ( .A1(MEM_stage_inst_dmem_ram_166), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n3786) );
NAND2_X1 MEM_stage_inst_dmem_U3930 ( .A1(MEM_stage_inst_dmem_ram_374), .A2(MEM_stage_inst_dmem_n4721), .ZN(MEM_stage_inst_dmem_n3787) );
NAND2_X1 MEM_stage_inst_dmem_U3929 ( .A1(MEM_stage_inst_dmem_n3785), .A2(MEM_stage_inst_dmem_n3784), .ZN(MEM_stage_inst_dmem_n3789) );
NAND2_X1 MEM_stage_inst_dmem_U3928 ( .A1(MEM_stage_inst_dmem_ram_198), .A2(MEM_stage_inst_dmem_n36), .ZN(MEM_stage_inst_dmem_n3784) );
NAND2_X1 MEM_stage_inst_dmem_U3927 ( .A1(MEM_stage_inst_dmem_ram_662), .A2(MEM_stage_inst_dmem_n3076), .ZN(MEM_stage_inst_dmem_n3785) );
NOR2_X1 MEM_stage_inst_dmem_U3926 ( .A1(MEM_stage_inst_dmem_n3783), .A2(MEM_stage_inst_dmem_n3782), .ZN(MEM_stage_inst_dmem_n3791) );
NAND2_X1 MEM_stage_inst_dmem_U3925 ( .A1(MEM_stage_inst_dmem_n3781), .A2(MEM_stage_inst_dmem_n3780), .ZN(MEM_stage_inst_dmem_n3782) );
NAND2_X1 MEM_stage_inst_dmem_U3924 ( .A1(MEM_stage_inst_dmem_ram_358), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n3780) );
NAND2_X1 MEM_stage_inst_dmem_U3923 ( .A1(MEM_stage_inst_dmem_ram_630), .A2(MEM_stage_inst_dmem_n4652), .ZN(MEM_stage_inst_dmem_n3781) );
NAND2_X1 MEM_stage_inst_dmem_U3922 ( .A1(MEM_stage_inst_dmem_n3779), .A2(MEM_stage_inst_dmem_n3778), .ZN(MEM_stage_inst_dmem_n3783) );
NAND2_X1 MEM_stage_inst_dmem_U3921 ( .A1(MEM_stage_inst_dmem_ram_966), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n3778) );
NAND2_X1 MEM_stage_inst_dmem_U3920 ( .A1(MEM_stage_inst_dmem_ram_182), .A2(MEM_stage_inst_dmem_n55), .ZN(MEM_stage_inst_dmem_n3779) );
NOR2_X1 MEM_stage_inst_dmem_U3919 ( .A1(MEM_stage_inst_dmem_n3777), .A2(MEM_stage_inst_dmem_n3776), .ZN(MEM_stage_inst_dmem_n3809) );
NAND2_X1 MEM_stage_inst_dmem_U3918 ( .A1(MEM_stage_inst_dmem_n3775), .A2(MEM_stage_inst_dmem_n3774), .ZN(MEM_stage_inst_dmem_n3776) );
NOR2_X1 MEM_stage_inst_dmem_U3917 ( .A1(MEM_stage_inst_dmem_n3773), .A2(MEM_stage_inst_dmem_n3772), .ZN(MEM_stage_inst_dmem_n3774) );
NAND2_X1 MEM_stage_inst_dmem_U3916 ( .A1(MEM_stage_inst_dmem_n3771), .A2(MEM_stage_inst_dmem_n3770), .ZN(MEM_stage_inst_dmem_n3772) );
NAND2_X1 MEM_stage_inst_dmem_U3915 ( .A1(MEM_stage_inst_dmem_ram_838), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n3770) );
NAND2_X1 MEM_stage_inst_dmem_U3914 ( .A1(MEM_stage_inst_dmem_ram_118), .A2(MEM_stage_inst_dmem_n4710), .ZN(MEM_stage_inst_dmem_n3771) );
NAND2_X1 MEM_stage_inst_dmem_U3913 ( .A1(MEM_stage_inst_dmem_n3769), .A2(MEM_stage_inst_dmem_n3768), .ZN(MEM_stage_inst_dmem_n3773) );
NAND2_X1 MEM_stage_inst_dmem_U3912 ( .A1(MEM_stage_inst_dmem_ram_54), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n3768) );
NAND2_X1 MEM_stage_inst_dmem_U3911 ( .A1(MEM_stage_inst_dmem_ram_902), .A2(MEM_stage_inst_dmem_n72), .ZN(MEM_stage_inst_dmem_n3769) );
NOR2_X1 MEM_stage_inst_dmem_U3910 ( .A1(MEM_stage_inst_dmem_n3767), .A2(MEM_stage_inst_dmem_n3766), .ZN(MEM_stage_inst_dmem_n3775) );
NAND2_X1 MEM_stage_inst_dmem_U3909 ( .A1(MEM_stage_inst_dmem_n3765), .A2(MEM_stage_inst_dmem_n3764), .ZN(MEM_stage_inst_dmem_n3766) );
NAND2_X1 MEM_stage_inst_dmem_U3908 ( .A1(MEM_stage_inst_dmem_ram_710), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n3764) );
NAND2_X1 MEM_stage_inst_dmem_U3907 ( .A1(MEM_stage_inst_dmem_ram_390), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n3765) );
NAND2_X1 MEM_stage_inst_dmem_U3906 ( .A1(MEM_stage_inst_dmem_n3763), .A2(MEM_stage_inst_dmem_n3762), .ZN(MEM_stage_inst_dmem_n3767) );
NAND2_X1 MEM_stage_inst_dmem_U3905 ( .A1(MEM_stage_inst_dmem_ram_758), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n3762) );
NAND2_X1 MEM_stage_inst_dmem_U3904 ( .A1(MEM_stage_inst_dmem_ram_694), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n3763) );
NAND2_X1 MEM_stage_inst_dmem_U3903 ( .A1(MEM_stage_inst_dmem_n3761), .A2(MEM_stage_inst_dmem_n3760), .ZN(MEM_stage_inst_dmem_n3777) );
NOR2_X1 MEM_stage_inst_dmem_U3902 ( .A1(MEM_stage_inst_dmem_n3759), .A2(MEM_stage_inst_dmem_n3758), .ZN(MEM_stage_inst_dmem_n3760) );
NAND2_X1 MEM_stage_inst_dmem_U3901 ( .A1(MEM_stage_inst_dmem_n3757), .A2(MEM_stage_inst_dmem_n3756), .ZN(MEM_stage_inst_dmem_n3758) );
NAND2_X1 MEM_stage_inst_dmem_U3900 ( .A1(MEM_stage_inst_dmem_ram_806), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n3756) );
NAND2_X1 MEM_stage_inst_dmem_U3899 ( .A1(MEM_stage_inst_dmem_ram_342), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n3757) );
NAND2_X1 MEM_stage_inst_dmem_U3898 ( .A1(MEM_stage_inst_dmem_n3755), .A2(MEM_stage_inst_dmem_n3754), .ZN(MEM_stage_inst_dmem_n3759) );
NAND2_X1 MEM_stage_inst_dmem_U3897 ( .A1(MEM_stage_inst_dmem_ram_774), .A2(MEM_stage_inst_dmem_n37), .ZN(MEM_stage_inst_dmem_n3754) );
NAND2_X1 MEM_stage_inst_dmem_U3896 ( .A1(MEM_stage_inst_dmem_ram_502), .A2(MEM_stage_inst_dmem_n8535), .ZN(MEM_stage_inst_dmem_n3755) );
NOR2_X1 MEM_stage_inst_dmem_U3895 ( .A1(MEM_stage_inst_dmem_n3753), .A2(MEM_stage_inst_dmem_n3752), .ZN(MEM_stage_inst_dmem_n3761) );
NAND2_X1 MEM_stage_inst_dmem_U3894 ( .A1(MEM_stage_inst_dmem_n3751), .A2(MEM_stage_inst_dmem_n3750), .ZN(MEM_stage_inst_dmem_n3752) );
NAND2_X1 MEM_stage_inst_dmem_U3893 ( .A1(MEM_stage_inst_dmem_ram_854), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n3750) );
NAND2_X1 MEM_stage_inst_dmem_U3892 ( .A1(MEM_stage_inst_dmem_ram_22), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n3751) );
NAND2_X1 MEM_stage_inst_dmem_U3891 ( .A1(MEM_stage_inst_dmem_n3749), .A2(MEM_stage_inst_dmem_n3748), .ZN(MEM_stage_inst_dmem_n3753) );
NAND2_X1 MEM_stage_inst_dmem_U3890 ( .A1(MEM_stage_inst_dmem_ram_262), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n3748) );
NAND2_X1 MEM_stage_inst_dmem_U3889 ( .A1(MEM_stage_inst_dmem_ram_582), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n3749) );
NOR2_X1 MEM_stage_inst_dmem_U3888 ( .A1(MEM_stage_inst_dmem_n3747), .A2(MEM_stage_inst_dmem_n8417), .ZN(MEM_stage_inst_dmem_n3876) );
NOR2_X1 MEM_stage_inst_dmem_U3887 ( .A1(MEM_stage_inst_dmem_n3746), .A2(MEM_stage_inst_dmem_n3745), .ZN(MEM_stage_inst_dmem_n3747) );
NAND2_X1 MEM_stage_inst_dmem_U3886 ( .A1(MEM_stage_inst_dmem_n3744), .A2(MEM_stage_inst_dmem_n3743), .ZN(MEM_stage_inst_dmem_n3745) );
NOR2_X1 MEM_stage_inst_dmem_U3885 ( .A1(MEM_stage_inst_dmem_n3742), .A2(MEM_stage_inst_dmem_n3741), .ZN(MEM_stage_inst_dmem_n3743) );
NAND2_X1 MEM_stage_inst_dmem_U3884 ( .A1(MEM_stage_inst_dmem_n3740), .A2(MEM_stage_inst_dmem_n3739), .ZN(MEM_stage_inst_dmem_n3741) );
NOR2_X1 MEM_stage_inst_dmem_U3883 ( .A1(MEM_stage_inst_dmem_n3738), .A2(MEM_stage_inst_dmem_n3737), .ZN(MEM_stage_inst_dmem_n3739) );
NAND2_X1 MEM_stage_inst_dmem_U3882 ( .A1(MEM_stage_inst_dmem_n3736), .A2(MEM_stage_inst_dmem_n3735), .ZN(MEM_stage_inst_dmem_n3737) );
NAND2_X1 MEM_stage_inst_dmem_U3881 ( .A1(MEM_stage_inst_dmem_ram_4022), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n3735) );
NAND2_X1 MEM_stage_inst_dmem_U3880 ( .A1(MEM_stage_inst_dmem_ram_3750), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n3736) );
NAND2_X1 MEM_stage_inst_dmem_U3879 ( .A1(MEM_stage_inst_dmem_n3734), .A2(MEM_stage_inst_dmem_n3733), .ZN(MEM_stage_inst_dmem_n3738) );
NAND2_X1 MEM_stage_inst_dmem_U3878 ( .A1(MEM_stage_inst_dmem_ram_3846), .A2(MEM_stage_inst_dmem_n37), .ZN(MEM_stage_inst_dmem_n3733) );
NAND2_X1 MEM_stage_inst_dmem_U3877 ( .A1(MEM_stage_inst_dmem_ram_3334), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n3734) );
NOR2_X1 MEM_stage_inst_dmem_U3876 ( .A1(MEM_stage_inst_dmem_n3732), .A2(MEM_stage_inst_dmem_n3731), .ZN(MEM_stage_inst_dmem_n3740) );
NAND2_X1 MEM_stage_inst_dmem_U3875 ( .A1(MEM_stage_inst_dmem_n3730), .A2(MEM_stage_inst_dmem_n3729), .ZN(MEM_stage_inst_dmem_n3731) );
NAND2_X1 MEM_stage_inst_dmem_U3874 ( .A1(MEM_stage_inst_dmem_ram_3958), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n3729) );
NAND2_X1 MEM_stage_inst_dmem_U3873 ( .A1(MEM_stage_inst_dmem_ram_3574), .A2(MEM_stage_inst_dmem_n64), .ZN(MEM_stage_inst_dmem_n3730) );
NAND2_X1 MEM_stage_inst_dmem_U3872 ( .A1(MEM_stage_inst_dmem_n3728), .A2(MEM_stage_inst_dmem_n3727), .ZN(MEM_stage_inst_dmem_n3732) );
NAND2_X1 MEM_stage_inst_dmem_U3871 ( .A1(MEM_stage_inst_dmem_ram_3622), .A2(MEM_stage_inst_dmem_n4692), .ZN(MEM_stage_inst_dmem_n3727) );
NAND2_X1 MEM_stage_inst_dmem_U3870 ( .A1(MEM_stage_inst_dmem_ram_3078), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n3728) );
NAND2_X1 MEM_stage_inst_dmem_U3869 ( .A1(MEM_stage_inst_dmem_n3726), .A2(MEM_stage_inst_dmem_n3725), .ZN(MEM_stage_inst_dmem_n3742) );
NOR2_X1 MEM_stage_inst_dmem_U3868 ( .A1(MEM_stage_inst_dmem_n3724), .A2(MEM_stage_inst_dmem_n3723), .ZN(MEM_stage_inst_dmem_n3725) );
NAND2_X1 MEM_stage_inst_dmem_U3867 ( .A1(MEM_stage_inst_dmem_n3722), .A2(MEM_stage_inst_dmem_n3721), .ZN(MEM_stage_inst_dmem_n3723) );
NAND2_X1 MEM_stage_inst_dmem_U3866 ( .A1(MEM_stage_inst_dmem_ram_4070), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n3721) );
NAND2_X1 MEM_stage_inst_dmem_U3865 ( .A1(MEM_stage_inst_dmem_ram_3238), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n3722) );
NAND2_X1 MEM_stage_inst_dmem_U3864 ( .A1(MEM_stage_inst_dmem_n3720), .A2(MEM_stage_inst_dmem_n3719), .ZN(MEM_stage_inst_dmem_n3724) );
NAND2_X1 MEM_stage_inst_dmem_U3863 ( .A1(MEM_stage_inst_dmem_ram_3830), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n3719) );
NAND2_X1 MEM_stage_inst_dmem_U3862 ( .A1(MEM_stage_inst_dmem_ram_3814), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n3720) );
NOR2_X1 MEM_stage_inst_dmem_U3861 ( .A1(MEM_stage_inst_dmem_n3718), .A2(MEM_stage_inst_dmem_n3717), .ZN(MEM_stage_inst_dmem_n3726) );
NAND2_X1 MEM_stage_inst_dmem_U3860 ( .A1(MEM_stage_inst_dmem_n3716), .A2(MEM_stage_inst_dmem_n3715), .ZN(MEM_stage_inst_dmem_n3717) );
NAND2_X1 MEM_stage_inst_dmem_U3859 ( .A1(MEM_stage_inst_dmem_ram_3126), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n3715) );
NAND2_X1 MEM_stage_inst_dmem_U3858 ( .A1(MEM_stage_inst_dmem_ram_3894), .A2(MEM_stage_inst_dmem_n4740), .ZN(MEM_stage_inst_dmem_n3716) );
NAND2_X1 MEM_stage_inst_dmem_U3857 ( .A1(MEM_stage_inst_dmem_n3714), .A2(MEM_stage_inst_dmem_n3713), .ZN(MEM_stage_inst_dmem_n3718) );
NAND2_X1 MEM_stage_inst_dmem_U3856 ( .A1(MEM_stage_inst_dmem_ram_3878), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n3713) );
NAND2_X1 MEM_stage_inst_dmem_U3855 ( .A1(MEM_stage_inst_dmem_ram_3190), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n3714) );
NOR2_X1 MEM_stage_inst_dmem_U3854 ( .A1(MEM_stage_inst_dmem_n3712), .A2(MEM_stage_inst_dmem_n3711), .ZN(MEM_stage_inst_dmem_n3744) );
NAND2_X1 MEM_stage_inst_dmem_U3853 ( .A1(MEM_stage_inst_dmem_n3710), .A2(MEM_stage_inst_dmem_n3709), .ZN(MEM_stage_inst_dmem_n3711) );
NOR2_X1 MEM_stage_inst_dmem_U3852 ( .A1(MEM_stage_inst_dmem_n3708), .A2(MEM_stage_inst_dmem_n3707), .ZN(MEM_stage_inst_dmem_n3709) );
NAND2_X1 MEM_stage_inst_dmem_U3851 ( .A1(MEM_stage_inst_dmem_n3706), .A2(MEM_stage_inst_dmem_n3705), .ZN(MEM_stage_inst_dmem_n3707) );
NAND2_X1 MEM_stage_inst_dmem_U3850 ( .A1(MEM_stage_inst_dmem_ram_3478), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n3705) );
NAND2_X1 MEM_stage_inst_dmem_U3849 ( .A1(MEM_stage_inst_dmem_ram_3318), .A2(MEM_stage_inst_dmem_n4649), .ZN(MEM_stage_inst_dmem_n3706) );
NAND2_X1 MEM_stage_inst_dmem_U3848 ( .A1(MEM_stage_inst_dmem_n3704), .A2(MEM_stage_inst_dmem_n3703), .ZN(MEM_stage_inst_dmem_n3708) );
NAND2_X1 MEM_stage_inst_dmem_U3847 ( .A1(MEM_stage_inst_dmem_ram_3638), .A2(MEM_stage_inst_dmem_n41), .ZN(MEM_stage_inst_dmem_n3703) );
NAND2_X1 MEM_stage_inst_dmem_U3846 ( .A1(MEM_stage_inst_dmem_ram_3350), .A2(MEM_stage_inst_dmem_n4672), .ZN(MEM_stage_inst_dmem_n3704) );
NOR2_X1 MEM_stage_inst_dmem_U3845 ( .A1(MEM_stage_inst_dmem_n3702), .A2(MEM_stage_inst_dmem_n3701), .ZN(MEM_stage_inst_dmem_n3710) );
NAND2_X1 MEM_stage_inst_dmem_U3844 ( .A1(MEM_stage_inst_dmem_n3700), .A2(MEM_stage_inst_dmem_n3699), .ZN(MEM_stage_inst_dmem_n3701) );
NAND2_X1 MEM_stage_inst_dmem_U3843 ( .A1(MEM_stage_inst_dmem_ram_3990), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n3699) );
NAND2_X1 MEM_stage_inst_dmem_U3842 ( .A1(MEM_stage_inst_dmem_ram_3158), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n3700) );
NAND2_X1 MEM_stage_inst_dmem_U3841 ( .A1(MEM_stage_inst_dmem_n3698), .A2(MEM_stage_inst_dmem_n3697), .ZN(MEM_stage_inst_dmem_n3702) );
NAND2_X1 MEM_stage_inst_dmem_U3840 ( .A1(MEM_stage_inst_dmem_ram_3686), .A2(MEM_stage_inst_dmem_n4701), .ZN(MEM_stage_inst_dmem_n3697) );
NAND2_X1 MEM_stage_inst_dmem_U3839 ( .A1(MEM_stage_inst_dmem_ram_3654), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n3698) );
NAND2_X1 MEM_stage_inst_dmem_U3838 ( .A1(MEM_stage_inst_dmem_n3696), .A2(MEM_stage_inst_dmem_n3695), .ZN(MEM_stage_inst_dmem_n3712) );
NOR2_X1 MEM_stage_inst_dmem_U3837 ( .A1(MEM_stage_inst_dmem_n3694), .A2(MEM_stage_inst_dmem_n3693), .ZN(MEM_stage_inst_dmem_n3695) );
NAND2_X1 MEM_stage_inst_dmem_U3836 ( .A1(MEM_stage_inst_dmem_n3692), .A2(MEM_stage_inst_dmem_n3691), .ZN(MEM_stage_inst_dmem_n3693) );
NAND2_X1 MEM_stage_inst_dmem_U3835 ( .A1(MEM_stage_inst_dmem_ram_3494), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n3691) );
NAND2_X1 MEM_stage_inst_dmem_U3834 ( .A1(MEM_stage_inst_dmem_ram_3798), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n3692) );
NAND2_X1 MEM_stage_inst_dmem_U3833 ( .A1(MEM_stage_inst_dmem_n3690), .A2(MEM_stage_inst_dmem_n3689), .ZN(MEM_stage_inst_dmem_n3694) );
NAND2_X1 MEM_stage_inst_dmem_U3832 ( .A1(MEM_stage_inst_dmem_ram_3382), .A2(MEM_stage_inst_dmem_n4731), .ZN(MEM_stage_inst_dmem_n3689) );
NAND2_X1 MEM_stage_inst_dmem_U3831 ( .A1(MEM_stage_inst_dmem_ram_3702), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n3690) );
NOR2_X1 MEM_stage_inst_dmem_U3830 ( .A1(MEM_stage_inst_dmem_n3688), .A2(MEM_stage_inst_dmem_n3687), .ZN(MEM_stage_inst_dmem_n3696) );
NAND2_X1 MEM_stage_inst_dmem_U3829 ( .A1(MEM_stage_inst_dmem_n3686), .A2(MEM_stage_inst_dmem_n3685), .ZN(MEM_stage_inst_dmem_n3687) );
NAND2_X1 MEM_stage_inst_dmem_U3828 ( .A1(MEM_stage_inst_dmem_ram_3782), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n3685) );
NAND2_X1 MEM_stage_inst_dmem_U3827 ( .A1(MEM_stage_inst_dmem_ram_3718), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n3686) );
NAND2_X1 MEM_stage_inst_dmem_U3826 ( .A1(MEM_stage_inst_dmem_n3684), .A2(MEM_stage_inst_dmem_n3683), .ZN(MEM_stage_inst_dmem_n3688) );
NAND2_X1 MEM_stage_inst_dmem_U3825 ( .A1(MEM_stage_inst_dmem_ram_3942), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n3683) );
NAND2_X1 MEM_stage_inst_dmem_U3824 ( .A1(MEM_stage_inst_dmem_ram_3110), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n3684) );
NAND2_X1 MEM_stage_inst_dmem_U3823 ( .A1(MEM_stage_inst_dmem_n3682), .A2(MEM_stage_inst_dmem_n3681), .ZN(MEM_stage_inst_dmem_n3746) );
NOR2_X1 MEM_stage_inst_dmem_U3822 ( .A1(MEM_stage_inst_dmem_n3680), .A2(MEM_stage_inst_dmem_n3679), .ZN(MEM_stage_inst_dmem_n3681) );
NAND2_X1 MEM_stage_inst_dmem_U3821 ( .A1(MEM_stage_inst_dmem_n3678), .A2(MEM_stage_inst_dmem_n3677), .ZN(MEM_stage_inst_dmem_n3679) );
NOR2_X1 MEM_stage_inst_dmem_U3820 ( .A1(MEM_stage_inst_dmem_n3676), .A2(MEM_stage_inst_dmem_n3675), .ZN(MEM_stage_inst_dmem_n3677) );
NAND2_X1 MEM_stage_inst_dmem_U3819 ( .A1(MEM_stage_inst_dmem_n3674), .A2(MEM_stage_inst_dmem_n3673), .ZN(MEM_stage_inst_dmem_n3675) );
NAND2_X1 MEM_stage_inst_dmem_U3818 ( .A1(MEM_stage_inst_dmem_ram_3526), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n3673) );
NAND2_X1 MEM_stage_inst_dmem_U3817 ( .A1(MEM_stage_inst_dmem_ram_3222), .A2(MEM_stage_inst_dmem_n5807), .ZN(MEM_stage_inst_dmem_n3674) );
NAND2_X1 MEM_stage_inst_dmem_U3816 ( .A1(MEM_stage_inst_dmem_n3672), .A2(MEM_stage_inst_dmem_n3671), .ZN(MEM_stage_inst_dmem_n3676) );
NAND2_X1 MEM_stage_inst_dmem_U3815 ( .A1(MEM_stage_inst_dmem_ram_3414), .A2(MEM_stage_inst_dmem_n3216), .ZN(MEM_stage_inst_dmem_n3671) );
NAND2_X1 MEM_stage_inst_dmem_U3814 ( .A1(MEM_stage_inst_dmem_ram_3670), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n3672) );
NOR2_X1 MEM_stage_inst_dmem_U3813 ( .A1(MEM_stage_inst_dmem_n3670), .A2(MEM_stage_inst_dmem_n3669), .ZN(MEM_stage_inst_dmem_n3678) );
NAND2_X1 MEM_stage_inst_dmem_U3812 ( .A1(MEM_stage_inst_dmem_n3668), .A2(MEM_stage_inst_dmem_n3667), .ZN(MEM_stage_inst_dmem_n3669) );
NAND2_X1 MEM_stage_inst_dmem_U3811 ( .A1(MEM_stage_inst_dmem_ram_3558), .A2(MEM_stage_inst_dmem_n4667), .ZN(MEM_stage_inst_dmem_n3667) );
NAND2_X1 MEM_stage_inst_dmem_U3810 ( .A1(MEM_stage_inst_dmem_ram_4054), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n3668) );
NAND2_X1 MEM_stage_inst_dmem_U3809 ( .A1(MEM_stage_inst_dmem_n3666), .A2(MEM_stage_inst_dmem_n3665), .ZN(MEM_stage_inst_dmem_n3670) );
NAND2_X1 MEM_stage_inst_dmem_U3808 ( .A1(MEM_stage_inst_dmem_ram_3510), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n3665) );
NAND2_X1 MEM_stage_inst_dmem_U3807 ( .A1(MEM_stage_inst_dmem_ram_3366), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n3666) );
NAND2_X1 MEM_stage_inst_dmem_U3806 ( .A1(MEM_stage_inst_dmem_n3664), .A2(MEM_stage_inst_dmem_n3663), .ZN(MEM_stage_inst_dmem_n3680) );
NOR2_X1 MEM_stage_inst_dmem_U3805 ( .A1(MEM_stage_inst_dmem_n3662), .A2(MEM_stage_inst_dmem_n3661), .ZN(MEM_stage_inst_dmem_n3663) );
NAND2_X1 MEM_stage_inst_dmem_U3804 ( .A1(MEM_stage_inst_dmem_n3660), .A2(MEM_stage_inst_dmem_n3659), .ZN(MEM_stage_inst_dmem_n3661) );
NAND2_X1 MEM_stage_inst_dmem_U3803 ( .A1(MEM_stage_inst_dmem_ram_3270), .A2(MEM_stage_inst_dmem_n36), .ZN(MEM_stage_inst_dmem_n3659) );
NAND2_X1 MEM_stage_inst_dmem_U3802 ( .A1(MEM_stage_inst_dmem_ram_3734), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n3660) );
NAND2_X1 MEM_stage_inst_dmem_U3801 ( .A1(MEM_stage_inst_dmem_n3658), .A2(MEM_stage_inst_dmem_n3657), .ZN(MEM_stage_inst_dmem_n3662) );
NAND2_X1 MEM_stage_inst_dmem_U3800 ( .A1(MEM_stage_inst_dmem_ram_3766), .A2(MEM_stage_inst_dmem_n4709), .ZN(MEM_stage_inst_dmem_n3657) );
NAND2_X1 MEM_stage_inst_dmem_U3799 ( .A1(MEM_stage_inst_dmem_ram_3462), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n3658) );
NOR2_X1 MEM_stage_inst_dmem_U3798 ( .A1(MEM_stage_inst_dmem_n3656), .A2(MEM_stage_inst_dmem_n3655), .ZN(MEM_stage_inst_dmem_n3664) );
NAND2_X1 MEM_stage_inst_dmem_U3797 ( .A1(MEM_stage_inst_dmem_n3654), .A2(MEM_stage_inst_dmem_n3653), .ZN(MEM_stage_inst_dmem_n3655) );
NAND2_X1 MEM_stage_inst_dmem_U3796 ( .A1(MEM_stage_inst_dmem_ram_3206), .A2(MEM_stage_inst_dmem_n61), .ZN(MEM_stage_inst_dmem_n3653) );
NAND2_X1 MEM_stage_inst_dmem_U3795 ( .A1(MEM_stage_inst_dmem_ram_3974), .A2(MEM_stage_inst_dmem_n72), .ZN(MEM_stage_inst_dmem_n3654) );
NAND2_X1 MEM_stage_inst_dmem_U3794 ( .A1(MEM_stage_inst_dmem_n3652), .A2(MEM_stage_inst_dmem_n3651), .ZN(MEM_stage_inst_dmem_n3656) );
NAND2_X1 MEM_stage_inst_dmem_U3793 ( .A1(MEM_stage_inst_dmem_ram_3398), .A2(MEM_stage_inst_dmem_n4706), .ZN(MEM_stage_inst_dmem_n3651) );
NAND2_X1 MEM_stage_inst_dmem_U3792 ( .A1(MEM_stage_inst_dmem_ram_3926), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n3652) );
NOR2_X1 MEM_stage_inst_dmem_U3791 ( .A1(MEM_stage_inst_dmem_n3650), .A2(MEM_stage_inst_dmem_n3649), .ZN(MEM_stage_inst_dmem_n3682) );
NAND2_X1 MEM_stage_inst_dmem_U3790 ( .A1(MEM_stage_inst_dmem_n3648), .A2(MEM_stage_inst_dmem_n3647), .ZN(MEM_stage_inst_dmem_n3649) );
NOR2_X1 MEM_stage_inst_dmem_U3789 ( .A1(MEM_stage_inst_dmem_n3646), .A2(MEM_stage_inst_dmem_n3645), .ZN(MEM_stage_inst_dmem_n3647) );
NAND2_X1 MEM_stage_inst_dmem_U3788 ( .A1(MEM_stage_inst_dmem_n3644), .A2(MEM_stage_inst_dmem_n3643), .ZN(MEM_stage_inst_dmem_n3645) );
NAND2_X1 MEM_stage_inst_dmem_U3787 ( .A1(MEM_stage_inst_dmem_ram_4006), .A2(MEM_stage_inst_dmem_n4675), .ZN(MEM_stage_inst_dmem_n3643) );
NAND2_X1 MEM_stage_inst_dmem_U3786 ( .A1(MEM_stage_inst_dmem_ram_3862), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n3644) );
NAND2_X1 MEM_stage_inst_dmem_U3785 ( .A1(MEM_stage_inst_dmem_n3642), .A2(MEM_stage_inst_dmem_n3641), .ZN(MEM_stage_inst_dmem_n3646) );
NAND2_X1 MEM_stage_inst_dmem_U3784 ( .A1(MEM_stage_inst_dmem_ram_3910), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n3641) );
NAND2_X1 MEM_stage_inst_dmem_U3783 ( .A1(MEM_stage_inst_dmem_ram_3286), .A2(MEM_stage_inst_dmem_n51), .ZN(MEM_stage_inst_dmem_n3642) );
NOR2_X1 MEM_stage_inst_dmem_U3782 ( .A1(MEM_stage_inst_dmem_n3640), .A2(MEM_stage_inst_dmem_n3639), .ZN(MEM_stage_inst_dmem_n3648) );
NAND2_X1 MEM_stage_inst_dmem_U3781 ( .A1(MEM_stage_inst_dmem_n3638), .A2(MEM_stage_inst_dmem_n3637), .ZN(MEM_stage_inst_dmem_n3639) );
NAND2_X1 MEM_stage_inst_dmem_U3780 ( .A1(MEM_stage_inst_dmem_ram_3142), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n3637) );
NAND2_X1 MEM_stage_inst_dmem_U3779 ( .A1(MEM_stage_inst_dmem_ram_4086), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n3638) );
NAND2_X1 MEM_stage_inst_dmem_U3778 ( .A1(MEM_stage_inst_dmem_n3636), .A2(MEM_stage_inst_dmem_n3635), .ZN(MEM_stage_inst_dmem_n3640) );
NAND2_X1 MEM_stage_inst_dmem_U3777 ( .A1(MEM_stage_inst_dmem_ram_3606), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n3635) );
NAND2_X1 MEM_stage_inst_dmem_U3776 ( .A1(MEM_stage_inst_dmem_ram_3446), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n3636) );
NAND2_X1 MEM_stage_inst_dmem_U3775 ( .A1(MEM_stage_inst_dmem_n3634), .A2(MEM_stage_inst_dmem_n3633), .ZN(MEM_stage_inst_dmem_n3650) );
NOR2_X1 MEM_stage_inst_dmem_U3774 ( .A1(MEM_stage_inst_dmem_n3632), .A2(MEM_stage_inst_dmem_n3631), .ZN(MEM_stage_inst_dmem_n3633) );
NAND2_X1 MEM_stage_inst_dmem_U3773 ( .A1(MEM_stage_inst_dmem_n3630), .A2(MEM_stage_inst_dmem_n3629), .ZN(MEM_stage_inst_dmem_n3631) );
NAND2_X1 MEM_stage_inst_dmem_U3772 ( .A1(MEM_stage_inst_dmem_ram_3094), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n3629) );
NAND2_X1 MEM_stage_inst_dmem_U3771 ( .A1(MEM_stage_inst_dmem_ram_3254), .A2(MEM_stage_inst_dmem_n55), .ZN(MEM_stage_inst_dmem_n3630) );
NAND2_X1 MEM_stage_inst_dmem_U3770 ( .A1(MEM_stage_inst_dmem_n3628), .A2(MEM_stage_inst_dmem_n3627), .ZN(MEM_stage_inst_dmem_n3632) );
NAND2_X1 MEM_stage_inst_dmem_U3769 ( .A1(MEM_stage_inst_dmem_ram_3302), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n3627) );
NAND2_X1 MEM_stage_inst_dmem_U3768 ( .A1(MEM_stage_inst_dmem_ram_3174), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n3628) );
NOR2_X1 MEM_stage_inst_dmem_U3767 ( .A1(MEM_stage_inst_dmem_n3626), .A2(MEM_stage_inst_dmem_n3625), .ZN(MEM_stage_inst_dmem_n3634) );
NAND2_X1 MEM_stage_inst_dmem_U3766 ( .A1(MEM_stage_inst_dmem_n3624), .A2(MEM_stage_inst_dmem_n3623), .ZN(MEM_stage_inst_dmem_n3625) );
NAND2_X1 MEM_stage_inst_dmem_U3765 ( .A1(MEM_stage_inst_dmem_ram_3542), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n3623) );
NAND2_X1 MEM_stage_inst_dmem_U3764 ( .A1(MEM_stage_inst_dmem_ram_3590), .A2(MEM_stage_inst_dmem_n71), .ZN(MEM_stage_inst_dmem_n3624) );
NAND2_X1 MEM_stage_inst_dmem_U3763 ( .A1(MEM_stage_inst_dmem_n3622), .A2(MEM_stage_inst_dmem_n3621), .ZN(MEM_stage_inst_dmem_n3626) );
NAND2_X1 MEM_stage_inst_dmem_U3762 ( .A1(MEM_stage_inst_dmem_ram_3430), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n3621) );
NAND2_X1 MEM_stage_inst_dmem_U3761 ( .A1(MEM_stage_inst_dmem_ram_4038), .A2(MEM_stage_inst_dmem_n4728), .ZN(MEM_stage_inst_dmem_n3622) );
NOR2_X1 MEM_stage_inst_dmem_U3760 ( .A1(MEM_stage_inst_dmem_n3620), .A2(MEM_stage_inst_dmem_n3619), .ZN(MEM_stage_inst_dmem_n3878) );
NOR2_X1 MEM_stage_inst_dmem_U3759 ( .A1(MEM_stage_inst_dmem_n3618), .A2(MEM_stage_inst_dmem_n8286), .ZN(MEM_stage_inst_dmem_n3619) );
NOR2_X1 MEM_stage_inst_dmem_U3758 ( .A1(MEM_stage_inst_dmem_n3617), .A2(MEM_stage_inst_dmem_n3616), .ZN(MEM_stage_inst_dmem_n3618) );
NAND2_X1 MEM_stage_inst_dmem_U3757 ( .A1(MEM_stage_inst_dmem_n3615), .A2(MEM_stage_inst_dmem_n3614), .ZN(MEM_stage_inst_dmem_n3616) );
NOR2_X1 MEM_stage_inst_dmem_U3756 ( .A1(MEM_stage_inst_dmem_n3613), .A2(MEM_stage_inst_dmem_n3612), .ZN(MEM_stage_inst_dmem_n3614) );
NAND2_X1 MEM_stage_inst_dmem_U3755 ( .A1(MEM_stage_inst_dmem_n3611), .A2(MEM_stage_inst_dmem_n3610), .ZN(MEM_stage_inst_dmem_n3612) );
NOR2_X1 MEM_stage_inst_dmem_U3754 ( .A1(MEM_stage_inst_dmem_n3609), .A2(MEM_stage_inst_dmem_n3608), .ZN(MEM_stage_inst_dmem_n3610) );
NAND2_X1 MEM_stage_inst_dmem_U3753 ( .A1(MEM_stage_inst_dmem_n3607), .A2(MEM_stage_inst_dmem_n3606), .ZN(MEM_stage_inst_dmem_n3608) );
NAND2_X1 MEM_stage_inst_dmem_U3752 ( .A1(MEM_stage_inst_dmem_ram_2246), .A2(MEM_stage_inst_dmem_n8256), .ZN(MEM_stage_inst_dmem_n3606) );
NAND2_X1 MEM_stage_inst_dmem_U3751 ( .A1(MEM_stage_inst_dmem_ram_2150), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n3607) );
NAND2_X1 MEM_stage_inst_dmem_U3750 ( .A1(MEM_stage_inst_dmem_n3605), .A2(MEM_stage_inst_dmem_n3604), .ZN(MEM_stage_inst_dmem_n3609) );
NAND2_X1 MEM_stage_inst_dmem_U3749 ( .A1(MEM_stage_inst_dmem_ram_2070), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n3604) );
NAND2_X1 MEM_stage_inst_dmem_U3748 ( .A1(MEM_stage_inst_dmem_ram_2630), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n3605) );
NOR2_X1 MEM_stage_inst_dmem_U3747 ( .A1(MEM_stage_inst_dmem_n3603), .A2(MEM_stage_inst_dmem_n3602), .ZN(MEM_stage_inst_dmem_n3611) );
NAND2_X1 MEM_stage_inst_dmem_U3746 ( .A1(MEM_stage_inst_dmem_n3601), .A2(MEM_stage_inst_dmem_n3600), .ZN(MEM_stage_inst_dmem_n3602) );
NAND2_X1 MEM_stage_inst_dmem_U3745 ( .A1(MEM_stage_inst_dmem_ram_2134), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n3600) );
NAND2_X1 MEM_stage_inst_dmem_U3744 ( .A1(MEM_stage_inst_dmem_ram_2790), .A2(MEM_stage_inst_dmem_n4769), .ZN(MEM_stage_inst_dmem_n3601) );
NAND2_X1 MEM_stage_inst_dmem_U3743 ( .A1(MEM_stage_inst_dmem_n3599), .A2(MEM_stage_inst_dmem_n3598), .ZN(MEM_stage_inst_dmem_n3603) );
NAND2_X1 MEM_stage_inst_dmem_U3742 ( .A1(MEM_stage_inst_dmem_ram_2534), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n3598) );
NAND2_X1 MEM_stage_inst_dmem_U3741 ( .A1(MEM_stage_inst_dmem_ram_2086), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n3599) );
NAND2_X1 MEM_stage_inst_dmem_U3740 ( .A1(MEM_stage_inst_dmem_n3597), .A2(MEM_stage_inst_dmem_n3596), .ZN(MEM_stage_inst_dmem_n3613) );
NOR2_X1 MEM_stage_inst_dmem_U3739 ( .A1(MEM_stage_inst_dmem_n3595), .A2(MEM_stage_inst_dmem_n3594), .ZN(MEM_stage_inst_dmem_n3596) );
NAND2_X1 MEM_stage_inst_dmem_U3738 ( .A1(MEM_stage_inst_dmem_n3593), .A2(MEM_stage_inst_dmem_n3592), .ZN(MEM_stage_inst_dmem_n3594) );
NAND2_X1 MEM_stage_inst_dmem_U3737 ( .A1(MEM_stage_inst_dmem_ram_2358), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n3592) );
NAND2_X1 MEM_stage_inst_dmem_U3736 ( .A1(MEM_stage_inst_dmem_ram_2214), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n3593) );
NAND2_X1 MEM_stage_inst_dmem_U3735 ( .A1(MEM_stage_inst_dmem_n3591), .A2(MEM_stage_inst_dmem_n3590), .ZN(MEM_stage_inst_dmem_n3595) );
NAND2_X1 MEM_stage_inst_dmem_U3734 ( .A1(MEM_stage_inst_dmem_ram_2758), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n3590) );
NAND2_X1 MEM_stage_inst_dmem_U3733 ( .A1(MEM_stage_inst_dmem_ram_2438), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n3591) );
NOR2_X1 MEM_stage_inst_dmem_U3732 ( .A1(MEM_stage_inst_dmem_n3589), .A2(MEM_stage_inst_dmem_n3588), .ZN(MEM_stage_inst_dmem_n3597) );
NAND2_X1 MEM_stage_inst_dmem_U3731 ( .A1(MEM_stage_inst_dmem_n3587), .A2(MEM_stage_inst_dmem_n3586), .ZN(MEM_stage_inst_dmem_n3588) );
NAND2_X1 MEM_stage_inst_dmem_U3730 ( .A1(MEM_stage_inst_dmem_ram_2518), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n3586) );
NAND2_X1 MEM_stage_inst_dmem_U3729 ( .A1(MEM_stage_inst_dmem_ram_2774), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n3587) );
NAND2_X1 MEM_stage_inst_dmem_U3728 ( .A1(MEM_stage_inst_dmem_n3585), .A2(MEM_stage_inst_dmem_n3584), .ZN(MEM_stage_inst_dmem_n3589) );
NAND2_X1 MEM_stage_inst_dmem_U3727 ( .A1(MEM_stage_inst_dmem_ram_2902), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n3584) );
NAND2_X1 MEM_stage_inst_dmem_U3726 ( .A1(MEM_stage_inst_dmem_ram_3014), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n3585) );
NOR2_X1 MEM_stage_inst_dmem_U3725 ( .A1(MEM_stage_inst_dmem_n3583), .A2(MEM_stage_inst_dmem_n3582), .ZN(MEM_stage_inst_dmem_n3615) );
NAND2_X1 MEM_stage_inst_dmem_U3724 ( .A1(MEM_stage_inst_dmem_n3581), .A2(MEM_stage_inst_dmem_n3580), .ZN(MEM_stage_inst_dmem_n3582) );
NOR2_X1 MEM_stage_inst_dmem_U3723 ( .A1(MEM_stage_inst_dmem_n3579), .A2(MEM_stage_inst_dmem_n3578), .ZN(MEM_stage_inst_dmem_n3580) );
NAND2_X1 MEM_stage_inst_dmem_U3722 ( .A1(MEM_stage_inst_dmem_n3577), .A2(MEM_stage_inst_dmem_n3576), .ZN(MEM_stage_inst_dmem_n3578) );
NAND2_X1 MEM_stage_inst_dmem_U3721 ( .A1(MEM_stage_inst_dmem_ram_2374), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n3576) );
NAND2_X1 MEM_stage_inst_dmem_U3720 ( .A1(MEM_stage_inst_dmem_ram_2886), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n3577) );
NAND2_X1 MEM_stage_inst_dmem_U3719 ( .A1(MEM_stage_inst_dmem_n3575), .A2(MEM_stage_inst_dmem_n3574), .ZN(MEM_stage_inst_dmem_n3579) );
NAND2_X1 MEM_stage_inst_dmem_U3718 ( .A1(MEM_stage_inst_dmem_ram_2342), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n3574) );
NAND2_X1 MEM_stage_inst_dmem_U3717 ( .A1(MEM_stage_inst_dmem_ram_2390), .A2(MEM_stage_inst_dmem_n3216), .ZN(MEM_stage_inst_dmem_n3575) );
NOR2_X1 MEM_stage_inst_dmem_U3716 ( .A1(MEM_stage_inst_dmem_n3573), .A2(MEM_stage_inst_dmem_n3572), .ZN(MEM_stage_inst_dmem_n3581) );
NAND2_X1 MEM_stage_inst_dmem_U3715 ( .A1(MEM_stage_inst_dmem_n3571), .A2(MEM_stage_inst_dmem_n3570), .ZN(MEM_stage_inst_dmem_n3572) );
NAND2_X1 MEM_stage_inst_dmem_U3714 ( .A1(MEM_stage_inst_dmem_ram_2486), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n3570) );
NAND2_X1 MEM_stage_inst_dmem_U3713 ( .A1(MEM_stage_inst_dmem_ram_2998), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n3571) );
NAND2_X1 MEM_stage_inst_dmem_U3712 ( .A1(MEM_stage_inst_dmem_n3569), .A2(MEM_stage_inst_dmem_n3568), .ZN(MEM_stage_inst_dmem_n3573) );
NAND2_X1 MEM_stage_inst_dmem_U3711 ( .A1(MEM_stage_inst_dmem_ram_2230), .A2(MEM_stage_inst_dmem_n55), .ZN(MEM_stage_inst_dmem_n3568) );
NAND2_X1 MEM_stage_inst_dmem_U3710 ( .A1(MEM_stage_inst_dmem_ram_2646), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n3569) );
NAND2_X1 MEM_stage_inst_dmem_U3709 ( .A1(MEM_stage_inst_dmem_n3567), .A2(MEM_stage_inst_dmem_n3566), .ZN(MEM_stage_inst_dmem_n3583) );
NOR2_X1 MEM_stage_inst_dmem_U3708 ( .A1(MEM_stage_inst_dmem_n3565), .A2(MEM_stage_inst_dmem_n3564), .ZN(MEM_stage_inst_dmem_n3566) );
NAND2_X1 MEM_stage_inst_dmem_U3707 ( .A1(MEM_stage_inst_dmem_n3563), .A2(MEM_stage_inst_dmem_n3562), .ZN(MEM_stage_inst_dmem_n3564) );
NAND2_X1 MEM_stage_inst_dmem_U3706 ( .A1(MEM_stage_inst_dmem_ram_3062), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n3562) );
NAND2_X1 MEM_stage_inst_dmem_U3705 ( .A1(MEM_stage_inst_dmem_ram_2198), .A2(MEM_stage_inst_dmem_n5807), .ZN(MEM_stage_inst_dmem_n3563) );
NAND2_X1 MEM_stage_inst_dmem_U3704 ( .A1(MEM_stage_inst_dmem_n3561), .A2(MEM_stage_inst_dmem_n3560), .ZN(MEM_stage_inst_dmem_n3565) );
NAND2_X1 MEM_stage_inst_dmem_U3703 ( .A1(MEM_stage_inst_dmem_ram_2406), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n3560) );
NAND2_X1 MEM_stage_inst_dmem_U3702 ( .A1(MEM_stage_inst_dmem_ram_2278), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n3561) );
NOR2_X1 MEM_stage_inst_dmem_U3701 ( .A1(MEM_stage_inst_dmem_n3559), .A2(MEM_stage_inst_dmem_n3558), .ZN(MEM_stage_inst_dmem_n3567) );
NAND2_X1 MEM_stage_inst_dmem_U3700 ( .A1(MEM_stage_inst_dmem_n3557), .A2(MEM_stage_inst_dmem_n3556), .ZN(MEM_stage_inst_dmem_n3558) );
NAND2_X1 MEM_stage_inst_dmem_U3699 ( .A1(MEM_stage_inst_dmem_ram_2982), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n3556) );
NAND2_X1 MEM_stage_inst_dmem_U3698 ( .A1(MEM_stage_inst_dmem_ram_2054), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n3557) );
NAND2_X1 MEM_stage_inst_dmem_U3697 ( .A1(MEM_stage_inst_dmem_n3555), .A2(MEM_stage_inst_dmem_n3554), .ZN(MEM_stage_inst_dmem_n3559) );
NAND2_X1 MEM_stage_inst_dmem_U3696 ( .A1(MEM_stage_inst_dmem_ram_2934), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n3554) );
NAND2_X1 MEM_stage_inst_dmem_U3695 ( .A1(MEM_stage_inst_dmem_ram_3030), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n3555) );
NAND2_X1 MEM_stage_inst_dmem_U3694 ( .A1(MEM_stage_inst_dmem_n3553), .A2(MEM_stage_inst_dmem_n3552), .ZN(MEM_stage_inst_dmem_n3617) );
NOR2_X1 MEM_stage_inst_dmem_U3693 ( .A1(MEM_stage_inst_dmem_n3551), .A2(MEM_stage_inst_dmem_n3550), .ZN(MEM_stage_inst_dmem_n3552) );
NAND2_X1 MEM_stage_inst_dmem_U3692 ( .A1(MEM_stage_inst_dmem_n3549), .A2(MEM_stage_inst_dmem_n3548), .ZN(MEM_stage_inst_dmem_n3550) );
NOR2_X1 MEM_stage_inst_dmem_U3691 ( .A1(MEM_stage_inst_dmem_n3547), .A2(MEM_stage_inst_dmem_n3546), .ZN(MEM_stage_inst_dmem_n3548) );
NAND2_X1 MEM_stage_inst_dmem_U3690 ( .A1(MEM_stage_inst_dmem_n3545), .A2(MEM_stage_inst_dmem_n3544), .ZN(MEM_stage_inst_dmem_n3546) );
NAND2_X1 MEM_stage_inst_dmem_U3689 ( .A1(MEM_stage_inst_dmem_ram_2822), .A2(MEM_stage_inst_dmem_n37), .ZN(MEM_stage_inst_dmem_n3544) );
NAND2_X1 MEM_stage_inst_dmem_U3688 ( .A1(MEM_stage_inst_dmem_ram_2854), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n3545) );
NAND2_X1 MEM_stage_inst_dmem_U3687 ( .A1(MEM_stage_inst_dmem_n3543), .A2(MEM_stage_inst_dmem_n3542), .ZN(MEM_stage_inst_dmem_n3547) );
NAND2_X1 MEM_stage_inst_dmem_U3686 ( .A1(MEM_stage_inst_dmem_ram_2326), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n3542) );
NAND2_X1 MEM_stage_inst_dmem_U3685 ( .A1(MEM_stage_inst_dmem_ram_2726), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n3543) );
NOR2_X1 MEM_stage_inst_dmem_U3684 ( .A1(MEM_stage_inst_dmem_n3541), .A2(MEM_stage_inst_dmem_n3540), .ZN(MEM_stage_inst_dmem_n3549) );
NAND2_X1 MEM_stage_inst_dmem_U3683 ( .A1(MEM_stage_inst_dmem_n3539), .A2(MEM_stage_inst_dmem_n3538), .ZN(MEM_stage_inst_dmem_n3540) );
NAND2_X1 MEM_stage_inst_dmem_U3682 ( .A1(MEM_stage_inst_dmem_ram_2966), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n3538) );
NAND2_X1 MEM_stage_inst_dmem_U3681 ( .A1(MEM_stage_inst_dmem_ram_2838), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n3539) );
NAND2_X1 MEM_stage_inst_dmem_U3680 ( .A1(MEM_stage_inst_dmem_n3537), .A2(MEM_stage_inst_dmem_n3536), .ZN(MEM_stage_inst_dmem_n3541) );
NAND2_X1 MEM_stage_inst_dmem_U3679 ( .A1(MEM_stage_inst_dmem_ram_3046), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n3536) );
NAND2_X1 MEM_stage_inst_dmem_U3678 ( .A1(MEM_stage_inst_dmem_ram_2502), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n3537) );
NAND2_X1 MEM_stage_inst_dmem_U3677 ( .A1(MEM_stage_inst_dmem_n3535), .A2(MEM_stage_inst_dmem_n3534), .ZN(MEM_stage_inst_dmem_n3551) );
NOR2_X1 MEM_stage_inst_dmem_U3676 ( .A1(MEM_stage_inst_dmem_n3533), .A2(MEM_stage_inst_dmem_n3532), .ZN(MEM_stage_inst_dmem_n3534) );
NAND2_X1 MEM_stage_inst_dmem_U3675 ( .A1(MEM_stage_inst_dmem_n3531), .A2(MEM_stage_inst_dmem_n3530), .ZN(MEM_stage_inst_dmem_n3532) );
NAND2_X1 MEM_stage_inst_dmem_U3674 ( .A1(MEM_stage_inst_dmem_ram_2614), .A2(MEM_stage_inst_dmem_n8169), .ZN(MEM_stage_inst_dmem_n3530) );
NAND2_X1 MEM_stage_inst_dmem_U3673 ( .A1(MEM_stage_inst_dmem_ram_2678), .A2(MEM_stage_inst_dmem_n4652), .ZN(MEM_stage_inst_dmem_n3531) );
NAND2_X1 MEM_stage_inst_dmem_U3672 ( .A1(MEM_stage_inst_dmem_n3529), .A2(MEM_stage_inst_dmem_n3528), .ZN(MEM_stage_inst_dmem_n3533) );
NAND2_X1 MEM_stage_inst_dmem_U3671 ( .A1(MEM_stage_inst_dmem_ram_2118), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n3528) );
NAND2_X1 MEM_stage_inst_dmem_U3670 ( .A1(MEM_stage_inst_dmem_ram_2166), .A2(MEM_stage_inst_dmem_n4710), .ZN(MEM_stage_inst_dmem_n3529) );
NOR2_X1 MEM_stage_inst_dmem_U3669 ( .A1(MEM_stage_inst_dmem_n3527), .A2(MEM_stage_inst_dmem_n3526), .ZN(MEM_stage_inst_dmem_n3535) );
NAND2_X1 MEM_stage_inst_dmem_U3668 ( .A1(MEM_stage_inst_dmem_n3525), .A2(MEM_stage_inst_dmem_n3524), .ZN(MEM_stage_inst_dmem_n3526) );
NAND2_X1 MEM_stage_inst_dmem_U3667 ( .A1(MEM_stage_inst_dmem_ram_2470), .A2(MEM_stage_inst_dmem_n4772), .ZN(MEM_stage_inst_dmem_n3524) );
NAND2_X1 MEM_stage_inst_dmem_U3666 ( .A1(MEM_stage_inst_dmem_ram_2662), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n3525) );
NAND2_X1 MEM_stage_inst_dmem_U3665 ( .A1(MEM_stage_inst_dmem_n3523), .A2(MEM_stage_inst_dmem_n3522), .ZN(MEM_stage_inst_dmem_n3527) );
NAND2_X1 MEM_stage_inst_dmem_U3664 ( .A1(MEM_stage_inst_dmem_ram_2550), .A2(MEM_stage_inst_dmem_n64), .ZN(MEM_stage_inst_dmem_n3522) );
NAND2_X1 MEM_stage_inst_dmem_U3663 ( .A1(MEM_stage_inst_dmem_ram_2950), .A2(MEM_stage_inst_dmem_n8193), .ZN(MEM_stage_inst_dmem_n3523) );
NOR2_X1 MEM_stage_inst_dmem_U3662 ( .A1(MEM_stage_inst_dmem_n3521), .A2(MEM_stage_inst_dmem_n3520), .ZN(MEM_stage_inst_dmem_n3553) );
NAND2_X1 MEM_stage_inst_dmem_U3661 ( .A1(MEM_stage_inst_dmem_n3519), .A2(MEM_stage_inst_dmem_n3518), .ZN(MEM_stage_inst_dmem_n3520) );
NOR2_X1 MEM_stage_inst_dmem_U3660 ( .A1(MEM_stage_inst_dmem_n3517), .A2(MEM_stage_inst_dmem_n3516), .ZN(MEM_stage_inst_dmem_n3518) );
NAND2_X1 MEM_stage_inst_dmem_U3659 ( .A1(MEM_stage_inst_dmem_n3515), .A2(MEM_stage_inst_dmem_n3514), .ZN(MEM_stage_inst_dmem_n3516) );
NAND2_X1 MEM_stage_inst_dmem_U3658 ( .A1(MEM_stage_inst_dmem_ram_2694), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n3514) );
NAND2_X1 MEM_stage_inst_dmem_U3657 ( .A1(MEM_stage_inst_dmem_ram_2566), .A2(MEM_stage_inst_dmem_n8225), .ZN(MEM_stage_inst_dmem_n3515) );
NAND2_X1 MEM_stage_inst_dmem_U3656 ( .A1(MEM_stage_inst_dmem_n3513), .A2(MEM_stage_inst_dmem_n3512), .ZN(MEM_stage_inst_dmem_n3517) );
NAND2_X1 MEM_stage_inst_dmem_U3655 ( .A1(MEM_stage_inst_dmem_ram_2102), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n3512) );
NAND2_X1 MEM_stage_inst_dmem_U3654 ( .A1(MEM_stage_inst_dmem_ram_2870), .A2(MEM_stage_inst_dmem_n46), .ZN(MEM_stage_inst_dmem_n3513) );
NOR2_X1 MEM_stage_inst_dmem_U3653 ( .A1(MEM_stage_inst_dmem_n3511), .A2(MEM_stage_inst_dmem_n3510), .ZN(MEM_stage_inst_dmem_n3519) );
NAND2_X1 MEM_stage_inst_dmem_U3652 ( .A1(MEM_stage_inst_dmem_n3509), .A2(MEM_stage_inst_dmem_n3508), .ZN(MEM_stage_inst_dmem_n3510) );
NAND2_X1 MEM_stage_inst_dmem_U3651 ( .A1(MEM_stage_inst_dmem_ram_2582), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n3508) );
NAND2_X1 MEM_stage_inst_dmem_U3650 ( .A1(MEM_stage_inst_dmem_ram_2422), .A2(MEM_stage_inst_dmem_n4721), .ZN(MEM_stage_inst_dmem_n3509) );
NAND2_X1 MEM_stage_inst_dmem_U3649 ( .A1(MEM_stage_inst_dmem_n3507), .A2(MEM_stage_inst_dmem_n3506), .ZN(MEM_stage_inst_dmem_n3511) );
NAND2_X1 MEM_stage_inst_dmem_U3648 ( .A1(MEM_stage_inst_dmem_ram_2806), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n3506) );
NAND2_X1 MEM_stage_inst_dmem_U3647 ( .A1(MEM_stage_inst_dmem_ram_2182), .A2(MEM_stage_inst_dmem_n8174), .ZN(MEM_stage_inst_dmem_n3507) );
NAND2_X1 MEM_stage_inst_dmem_U3646 ( .A1(MEM_stage_inst_dmem_n3505), .A2(MEM_stage_inst_dmem_n3504), .ZN(MEM_stage_inst_dmem_n3521) );
NOR2_X1 MEM_stage_inst_dmem_U3645 ( .A1(MEM_stage_inst_dmem_n3503), .A2(MEM_stage_inst_dmem_n3502), .ZN(MEM_stage_inst_dmem_n3504) );
NAND2_X1 MEM_stage_inst_dmem_U3644 ( .A1(MEM_stage_inst_dmem_n3501), .A2(MEM_stage_inst_dmem_n3500), .ZN(MEM_stage_inst_dmem_n3502) );
NAND2_X1 MEM_stage_inst_dmem_U3643 ( .A1(MEM_stage_inst_dmem_ram_2454), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n3500) );
NAND2_X1 MEM_stage_inst_dmem_U3642 ( .A1(MEM_stage_inst_dmem_ram_2598), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n3501) );
NAND2_X1 MEM_stage_inst_dmem_U3641 ( .A1(MEM_stage_inst_dmem_n3499), .A2(MEM_stage_inst_dmem_n3498), .ZN(MEM_stage_inst_dmem_n3503) );
NAND2_X1 MEM_stage_inst_dmem_U3640 ( .A1(MEM_stage_inst_dmem_ram_2918), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n3498) );
NAND2_X1 MEM_stage_inst_dmem_U3639 ( .A1(MEM_stage_inst_dmem_ram_2294), .A2(MEM_stage_inst_dmem_n39), .ZN(MEM_stage_inst_dmem_n3499) );
NOR2_X1 MEM_stage_inst_dmem_U3638 ( .A1(MEM_stage_inst_dmem_n3497), .A2(MEM_stage_inst_dmem_n3496), .ZN(MEM_stage_inst_dmem_n3505) );
NAND2_X1 MEM_stage_inst_dmem_U3637 ( .A1(MEM_stage_inst_dmem_n3495), .A2(MEM_stage_inst_dmem_n3494), .ZN(MEM_stage_inst_dmem_n3496) );
NAND2_X1 MEM_stage_inst_dmem_U3636 ( .A1(MEM_stage_inst_dmem_ram_2262), .A2(MEM_stage_inst_dmem_n8206), .ZN(MEM_stage_inst_dmem_n3494) );
NAND2_X1 MEM_stage_inst_dmem_U3635 ( .A1(MEM_stage_inst_dmem_ram_2310), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n3495) );
NAND2_X1 MEM_stage_inst_dmem_U3634 ( .A1(MEM_stage_inst_dmem_n3493), .A2(MEM_stage_inst_dmem_n3492), .ZN(MEM_stage_inst_dmem_n3497) );
NAND2_X1 MEM_stage_inst_dmem_U3633 ( .A1(MEM_stage_inst_dmem_ram_2742), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n3492) );
NAND2_X1 MEM_stage_inst_dmem_U3632 ( .A1(MEM_stage_inst_dmem_ram_2710), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n3493) );
NOR2_X1 MEM_stage_inst_dmem_U3631 ( .A1(MEM_stage_inst_dmem_n3491), .A2(MEM_stage_inst_dmem_n8152), .ZN(MEM_stage_inst_dmem_n3620) );
NOR2_X1 MEM_stage_inst_dmem_U3630 ( .A1(MEM_stage_inst_dmem_n3490), .A2(MEM_stage_inst_dmem_n3489), .ZN(MEM_stage_inst_dmem_n3491) );
NAND2_X1 MEM_stage_inst_dmem_U3629 ( .A1(MEM_stage_inst_dmem_n3488), .A2(MEM_stage_inst_dmem_n3487), .ZN(MEM_stage_inst_dmem_n3489) );
NOR2_X1 MEM_stage_inst_dmem_U3628 ( .A1(MEM_stage_inst_dmem_n3486), .A2(MEM_stage_inst_dmem_n3485), .ZN(MEM_stage_inst_dmem_n3487) );
NAND2_X1 MEM_stage_inst_dmem_U3627 ( .A1(MEM_stage_inst_dmem_n3484), .A2(MEM_stage_inst_dmem_n3483), .ZN(MEM_stage_inst_dmem_n3485) );
NOR2_X1 MEM_stage_inst_dmem_U3626 ( .A1(MEM_stage_inst_dmem_n3482), .A2(MEM_stage_inst_dmem_n3481), .ZN(MEM_stage_inst_dmem_n3483) );
NAND2_X1 MEM_stage_inst_dmem_U3625 ( .A1(MEM_stage_inst_dmem_n3480), .A2(MEM_stage_inst_dmem_n3479), .ZN(MEM_stage_inst_dmem_n3481) );
NAND2_X1 MEM_stage_inst_dmem_U3624 ( .A1(MEM_stage_inst_dmem_ram_1158), .A2(MEM_stage_inst_dmem_n61), .ZN(MEM_stage_inst_dmem_n3479) );
NAND2_X1 MEM_stage_inst_dmem_U3623 ( .A1(MEM_stage_inst_dmem_ram_2038), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n3480) );
NAND2_X1 MEM_stage_inst_dmem_U3622 ( .A1(MEM_stage_inst_dmem_n3478), .A2(MEM_stage_inst_dmem_n3477), .ZN(MEM_stage_inst_dmem_n3482) );
NAND2_X1 MEM_stage_inst_dmem_U3621 ( .A1(MEM_stage_inst_dmem_ram_1574), .A2(MEM_stage_inst_dmem_n4692), .ZN(MEM_stage_inst_dmem_n3477) );
NAND2_X1 MEM_stage_inst_dmem_U3620 ( .A1(MEM_stage_inst_dmem_ram_1638), .A2(MEM_stage_inst_dmem_n4701), .ZN(MEM_stage_inst_dmem_n3478) );
NOR2_X1 MEM_stage_inst_dmem_U3619 ( .A1(MEM_stage_inst_dmem_n3476), .A2(MEM_stage_inst_dmem_n3475), .ZN(MEM_stage_inst_dmem_n3484) );
NAND2_X1 MEM_stage_inst_dmem_U3618 ( .A1(MEM_stage_inst_dmem_n3474), .A2(MEM_stage_inst_dmem_n3473), .ZN(MEM_stage_inst_dmem_n3475) );
NAND2_X1 MEM_stage_inst_dmem_U3617 ( .A1(MEM_stage_inst_dmem_ram_1270), .A2(MEM_stage_inst_dmem_n4649), .ZN(MEM_stage_inst_dmem_n3473) );
NAND2_X1 MEM_stage_inst_dmem_U3616 ( .A1(MEM_stage_inst_dmem_ram_1622), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n3474) );
NAND2_X1 MEM_stage_inst_dmem_U3615 ( .A1(MEM_stage_inst_dmem_n3472), .A2(MEM_stage_inst_dmem_n3471), .ZN(MEM_stage_inst_dmem_n3476) );
NAND2_X1 MEM_stage_inst_dmem_U3614 ( .A1(MEM_stage_inst_dmem_ram_1782), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n3471) );
NAND2_X1 MEM_stage_inst_dmem_U3613 ( .A1(MEM_stage_inst_dmem_ram_1126), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n3472) );
NAND2_X1 MEM_stage_inst_dmem_U3612 ( .A1(MEM_stage_inst_dmem_n3470), .A2(MEM_stage_inst_dmem_n3469), .ZN(MEM_stage_inst_dmem_n3486) );
NOR2_X1 MEM_stage_inst_dmem_U3611 ( .A1(MEM_stage_inst_dmem_n3468), .A2(MEM_stage_inst_dmem_n3467), .ZN(MEM_stage_inst_dmem_n3469) );
NAND2_X1 MEM_stage_inst_dmem_U3610 ( .A1(MEM_stage_inst_dmem_n3466), .A2(MEM_stage_inst_dmem_n3465), .ZN(MEM_stage_inst_dmem_n3467) );
NAND2_X1 MEM_stage_inst_dmem_U3609 ( .A1(MEM_stage_inst_dmem_ram_1238), .A2(MEM_stage_inst_dmem_n51), .ZN(MEM_stage_inst_dmem_n3465) );
NAND2_X1 MEM_stage_inst_dmem_U3608 ( .A1(MEM_stage_inst_dmem_ram_1190), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n3466) );
NAND2_X1 MEM_stage_inst_dmem_U3607 ( .A1(MEM_stage_inst_dmem_n3464), .A2(MEM_stage_inst_dmem_n3463), .ZN(MEM_stage_inst_dmem_n3468) );
NAND2_X1 MEM_stage_inst_dmem_U3606 ( .A1(MEM_stage_inst_dmem_ram_1878), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n3463) );
NAND2_X1 MEM_stage_inst_dmem_U3605 ( .A1(MEM_stage_inst_dmem_ram_1974), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n3464) );
NOR2_X1 MEM_stage_inst_dmem_U3604 ( .A1(MEM_stage_inst_dmem_n3462), .A2(MEM_stage_inst_dmem_n3461), .ZN(MEM_stage_inst_dmem_n3470) );
NAND2_X1 MEM_stage_inst_dmem_U3603 ( .A1(MEM_stage_inst_dmem_n3460), .A2(MEM_stage_inst_dmem_n3459), .ZN(MEM_stage_inst_dmem_n3461) );
NAND2_X1 MEM_stage_inst_dmem_U3602 ( .A1(MEM_stage_inst_dmem_ram_1222), .A2(MEM_stage_inst_dmem_n36), .ZN(MEM_stage_inst_dmem_n3459) );
NAND2_X1 MEM_stage_inst_dmem_U3601 ( .A1(MEM_stage_inst_dmem_ram_1302), .A2(MEM_stage_inst_dmem_n4672), .ZN(MEM_stage_inst_dmem_n3460) );
NAND2_X1 MEM_stage_inst_dmem_U3600 ( .A1(MEM_stage_inst_dmem_n3458), .A2(MEM_stage_inst_dmem_n3457), .ZN(MEM_stage_inst_dmem_n3462) );
NAND2_X1 MEM_stage_inst_dmem_U3599 ( .A1(MEM_stage_inst_dmem_ram_1910), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n3457) );
NAND2_X1 MEM_stage_inst_dmem_U3598 ( .A1(MEM_stage_inst_dmem_ram_1062), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n3458) );
NOR2_X1 MEM_stage_inst_dmem_U3597 ( .A1(MEM_stage_inst_dmem_n3456), .A2(MEM_stage_inst_dmem_n3455), .ZN(MEM_stage_inst_dmem_n3488) );
NAND2_X1 MEM_stage_inst_dmem_U3596 ( .A1(MEM_stage_inst_dmem_n3454), .A2(MEM_stage_inst_dmem_n3453), .ZN(MEM_stage_inst_dmem_n3455) );
NOR2_X1 MEM_stage_inst_dmem_U3595 ( .A1(MEM_stage_inst_dmem_n3452), .A2(MEM_stage_inst_dmem_n3451), .ZN(MEM_stage_inst_dmem_n3453) );
NAND2_X1 MEM_stage_inst_dmem_U3594 ( .A1(MEM_stage_inst_dmem_n3450), .A2(MEM_stage_inst_dmem_n3449), .ZN(MEM_stage_inst_dmem_n3451) );
NAND2_X1 MEM_stage_inst_dmem_U3593 ( .A1(MEM_stage_inst_dmem_ram_1494), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n3449) );
NAND2_X1 MEM_stage_inst_dmem_U3592 ( .A1(MEM_stage_inst_dmem_ram_1206), .A2(MEM_stage_inst_dmem_n55), .ZN(MEM_stage_inst_dmem_n3450) );
NAND2_X1 MEM_stage_inst_dmem_U3591 ( .A1(MEM_stage_inst_dmem_n3448), .A2(MEM_stage_inst_dmem_n3447), .ZN(MEM_stage_inst_dmem_n3452) );
NAND2_X1 MEM_stage_inst_dmem_U3590 ( .A1(MEM_stage_inst_dmem_ram_1094), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n3447) );
NAND2_X1 MEM_stage_inst_dmem_U3589 ( .A1(MEM_stage_inst_dmem_ram_1110), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n3448) );
NOR2_X1 MEM_stage_inst_dmem_U3588 ( .A1(MEM_stage_inst_dmem_n3446), .A2(MEM_stage_inst_dmem_n3445), .ZN(MEM_stage_inst_dmem_n3454) );
NAND2_X1 MEM_stage_inst_dmem_U3587 ( .A1(MEM_stage_inst_dmem_n3444), .A2(MEM_stage_inst_dmem_n3443), .ZN(MEM_stage_inst_dmem_n3445) );
NAND2_X1 MEM_stage_inst_dmem_U3586 ( .A1(MEM_stage_inst_dmem_ram_1462), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n3443) );
NAND2_X1 MEM_stage_inst_dmem_U3585 ( .A1(MEM_stage_inst_dmem_ram_2006), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n3444) );
NAND2_X1 MEM_stage_inst_dmem_U3584 ( .A1(MEM_stage_inst_dmem_n3442), .A2(MEM_stage_inst_dmem_n3441), .ZN(MEM_stage_inst_dmem_n3446) );
NAND2_X1 MEM_stage_inst_dmem_U3583 ( .A1(MEM_stage_inst_dmem_ram_1702), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n3441) );
NAND2_X1 MEM_stage_inst_dmem_U3582 ( .A1(MEM_stage_inst_dmem_ram_1846), .A2(MEM_stage_inst_dmem_n4740), .ZN(MEM_stage_inst_dmem_n3442) );
NAND2_X1 MEM_stage_inst_dmem_U3581 ( .A1(MEM_stage_inst_dmem_n3440), .A2(MEM_stage_inst_dmem_n3439), .ZN(MEM_stage_inst_dmem_n3456) );
NOR2_X1 MEM_stage_inst_dmem_U3580 ( .A1(MEM_stage_inst_dmem_n3438), .A2(MEM_stage_inst_dmem_n3437), .ZN(MEM_stage_inst_dmem_n3439) );
NAND2_X1 MEM_stage_inst_dmem_U3579 ( .A1(MEM_stage_inst_dmem_n3436), .A2(MEM_stage_inst_dmem_n3435), .ZN(MEM_stage_inst_dmem_n3437) );
NAND2_X1 MEM_stage_inst_dmem_U3578 ( .A1(MEM_stage_inst_dmem_ram_1526), .A2(MEM_stage_inst_dmem_n8535), .ZN(MEM_stage_inst_dmem_n3435) );
NAND2_X1 MEM_stage_inst_dmem_U3577 ( .A1(MEM_stage_inst_dmem_ram_1382), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n3436) );
NAND2_X1 MEM_stage_inst_dmem_U3576 ( .A1(MEM_stage_inst_dmem_n3434), .A2(MEM_stage_inst_dmem_n3433), .ZN(MEM_stage_inst_dmem_n3438) );
NAND2_X1 MEM_stage_inst_dmem_U3575 ( .A1(MEM_stage_inst_dmem_ram_1670), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n3433) );
NAND2_X1 MEM_stage_inst_dmem_U3574 ( .A1(MEM_stage_inst_dmem_ram_1446), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n3434) );
NOR2_X1 MEM_stage_inst_dmem_U3573 ( .A1(MEM_stage_inst_dmem_n3432), .A2(MEM_stage_inst_dmem_n3431), .ZN(MEM_stage_inst_dmem_n3440) );
NAND2_X1 MEM_stage_inst_dmem_U3572 ( .A1(MEM_stage_inst_dmem_n3430), .A2(MEM_stage_inst_dmem_n3429), .ZN(MEM_stage_inst_dmem_n3431) );
NAND2_X1 MEM_stage_inst_dmem_U3571 ( .A1(MEM_stage_inst_dmem_ram_1942), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n3429) );
NAND2_X1 MEM_stage_inst_dmem_U3570 ( .A1(MEM_stage_inst_dmem_ram_1766), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n3430) );
NAND2_X1 MEM_stage_inst_dmem_U3569 ( .A1(MEM_stage_inst_dmem_n3428), .A2(MEM_stage_inst_dmem_n3427), .ZN(MEM_stage_inst_dmem_n3432) );
NAND2_X1 MEM_stage_inst_dmem_U3568 ( .A1(MEM_stage_inst_dmem_ram_1350), .A2(MEM_stage_inst_dmem_n4706), .ZN(MEM_stage_inst_dmem_n3427) );
NAND2_X1 MEM_stage_inst_dmem_U3567 ( .A1(MEM_stage_inst_dmem_ram_1958), .A2(MEM_stage_inst_dmem_n4675), .ZN(MEM_stage_inst_dmem_n3428) );
NAND2_X1 MEM_stage_inst_dmem_U3566 ( .A1(MEM_stage_inst_dmem_n3426), .A2(MEM_stage_inst_dmem_n3425), .ZN(MEM_stage_inst_dmem_n3490) );
NOR2_X1 MEM_stage_inst_dmem_U3565 ( .A1(MEM_stage_inst_dmem_n3424), .A2(MEM_stage_inst_dmem_n3423), .ZN(MEM_stage_inst_dmem_n3425) );
NAND2_X1 MEM_stage_inst_dmem_U3564 ( .A1(MEM_stage_inst_dmem_n3422), .A2(MEM_stage_inst_dmem_n3421), .ZN(MEM_stage_inst_dmem_n3423) );
NOR2_X1 MEM_stage_inst_dmem_U3563 ( .A1(MEM_stage_inst_dmem_n3420), .A2(MEM_stage_inst_dmem_n3419), .ZN(MEM_stage_inst_dmem_n3421) );
NAND2_X1 MEM_stage_inst_dmem_U3562 ( .A1(MEM_stage_inst_dmem_n3418), .A2(MEM_stage_inst_dmem_n3417), .ZN(MEM_stage_inst_dmem_n3419) );
NAND2_X1 MEM_stage_inst_dmem_U3561 ( .A1(MEM_stage_inst_dmem_ram_1078), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n3417) );
NAND2_X1 MEM_stage_inst_dmem_U3560 ( .A1(MEM_stage_inst_dmem_ram_1414), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n3418) );
NAND2_X1 MEM_stage_inst_dmem_U3559 ( .A1(MEM_stage_inst_dmem_n3416), .A2(MEM_stage_inst_dmem_n3415), .ZN(MEM_stage_inst_dmem_n3420) );
NAND2_X1 MEM_stage_inst_dmem_U3558 ( .A1(MEM_stage_inst_dmem_ram_1830), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n3415) );
NAND2_X1 MEM_stage_inst_dmem_U3557 ( .A1(MEM_stage_inst_dmem_ram_1686), .A2(MEM_stage_inst_dmem_n3076), .ZN(MEM_stage_inst_dmem_n3416) );
NOR2_X1 MEM_stage_inst_dmem_U3556 ( .A1(MEM_stage_inst_dmem_n3414), .A2(MEM_stage_inst_dmem_n3413), .ZN(MEM_stage_inst_dmem_n3422) );
NAND2_X1 MEM_stage_inst_dmem_U3555 ( .A1(MEM_stage_inst_dmem_n3412), .A2(MEM_stage_inst_dmem_n3411), .ZN(MEM_stage_inst_dmem_n3413) );
NAND2_X1 MEM_stage_inst_dmem_U3554 ( .A1(MEM_stage_inst_dmem_ram_1334), .A2(MEM_stage_inst_dmem_n4731), .ZN(MEM_stage_inst_dmem_n3411) );
NAND2_X1 MEM_stage_inst_dmem_U3553 ( .A1(MEM_stage_inst_dmem_ram_1510), .A2(MEM_stage_inst_dmem_n4667), .ZN(MEM_stage_inst_dmem_n3412) );
NAND2_X1 MEM_stage_inst_dmem_U3552 ( .A1(MEM_stage_inst_dmem_n3410), .A2(MEM_stage_inst_dmem_n3409), .ZN(MEM_stage_inst_dmem_n3414) );
NAND2_X1 MEM_stage_inst_dmem_U3551 ( .A1(MEM_stage_inst_dmem_ram_1142), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n3409) );
NAND2_X1 MEM_stage_inst_dmem_U3550 ( .A1(MEM_stage_inst_dmem_ram_1654), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n3410) );
NAND2_X1 MEM_stage_inst_dmem_U3549 ( .A1(MEM_stage_inst_dmem_n3408), .A2(MEM_stage_inst_dmem_n3407), .ZN(MEM_stage_inst_dmem_n3424) );
NOR2_X1 MEM_stage_inst_dmem_U3548 ( .A1(MEM_stage_inst_dmem_n3406), .A2(MEM_stage_inst_dmem_n3405), .ZN(MEM_stage_inst_dmem_n3407) );
NAND2_X1 MEM_stage_inst_dmem_U3547 ( .A1(MEM_stage_inst_dmem_n3404), .A2(MEM_stage_inst_dmem_n3403), .ZN(MEM_stage_inst_dmem_n3405) );
NAND2_X1 MEM_stage_inst_dmem_U3546 ( .A1(MEM_stage_inst_dmem_ram_1590), .A2(MEM_stage_inst_dmem_n41), .ZN(MEM_stage_inst_dmem_n3403) );
NAND2_X1 MEM_stage_inst_dmem_U3545 ( .A1(MEM_stage_inst_dmem_ram_1862), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n3404) );
NAND2_X1 MEM_stage_inst_dmem_U3544 ( .A1(MEM_stage_inst_dmem_n3402), .A2(MEM_stage_inst_dmem_n3401), .ZN(MEM_stage_inst_dmem_n3406) );
NAND2_X1 MEM_stage_inst_dmem_U3543 ( .A1(MEM_stage_inst_dmem_ram_1734), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n3401) );
NAND2_X1 MEM_stage_inst_dmem_U3542 ( .A1(MEM_stage_inst_dmem_ram_1718), .A2(MEM_stage_inst_dmem_n4709), .ZN(MEM_stage_inst_dmem_n3402) );
NOR2_X1 MEM_stage_inst_dmem_U3541 ( .A1(MEM_stage_inst_dmem_n3400), .A2(MEM_stage_inst_dmem_n3399), .ZN(MEM_stage_inst_dmem_n3408) );
NAND2_X1 MEM_stage_inst_dmem_U3540 ( .A1(MEM_stage_inst_dmem_n3398), .A2(MEM_stage_inst_dmem_n3397), .ZN(MEM_stage_inst_dmem_n3399) );
NAND2_X1 MEM_stage_inst_dmem_U3539 ( .A1(MEM_stage_inst_dmem_ram_1894), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n3397) );
NAND2_X1 MEM_stage_inst_dmem_U3538 ( .A1(MEM_stage_inst_dmem_ram_1478), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n3398) );
NAND2_X1 MEM_stage_inst_dmem_U3537 ( .A1(MEM_stage_inst_dmem_n3396), .A2(MEM_stage_inst_dmem_n3395), .ZN(MEM_stage_inst_dmem_n3400) );
NAND2_X1 MEM_stage_inst_dmem_U3536 ( .A1(MEM_stage_inst_dmem_ram_1318), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n3395) );
NAND2_X1 MEM_stage_inst_dmem_U3535 ( .A1(MEM_stage_inst_dmem_ram_1814), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n3396) );
NOR2_X1 MEM_stage_inst_dmem_U3534 ( .A1(MEM_stage_inst_dmem_n3394), .A2(MEM_stage_inst_dmem_n3393), .ZN(MEM_stage_inst_dmem_n3426) );
NAND2_X1 MEM_stage_inst_dmem_U3533 ( .A1(MEM_stage_inst_dmem_n3392), .A2(MEM_stage_inst_dmem_n3391), .ZN(MEM_stage_inst_dmem_n3393) );
NOR2_X1 MEM_stage_inst_dmem_U3532 ( .A1(MEM_stage_inst_dmem_n3390), .A2(MEM_stage_inst_dmem_n3389), .ZN(MEM_stage_inst_dmem_n3391) );
NAND2_X1 MEM_stage_inst_dmem_U3531 ( .A1(MEM_stage_inst_dmem_n3388), .A2(MEM_stage_inst_dmem_n3387), .ZN(MEM_stage_inst_dmem_n3389) );
NAND2_X1 MEM_stage_inst_dmem_U3530 ( .A1(MEM_stage_inst_dmem_ram_1254), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n3387) );
NAND2_X1 MEM_stage_inst_dmem_U3529 ( .A1(MEM_stage_inst_dmem_ram_1558), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n3388) );
NAND2_X1 MEM_stage_inst_dmem_U3528 ( .A1(MEM_stage_inst_dmem_n3386), .A2(MEM_stage_inst_dmem_n3385), .ZN(MEM_stage_inst_dmem_n3390) );
NAND2_X1 MEM_stage_inst_dmem_U3527 ( .A1(MEM_stage_inst_dmem_ram_1366), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n3385) );
NAND2_X1 MEM_stage_inst_dmem_U3526 ( .A1(MEM_stage_inst_dmem_ram_1286), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n3386) );
NOR2_X1 MEM_stage_inst_dmem_U3525 ( .A1(MEM_stage_inst_dmem_n3384), .A2(MEM_stage_inst_dmem_n3383), .ZN(MEM_stage_inst_dmem_n3392) );
NAND2_X1 MEM_stage_inst_dmem_U3524 ( .A1(MEM_stage_inst_dmem_n3382), .A2(MEM_stage_inst_dmem_n3381), .ZN(MEM_stage_inst_dmem_n3383) );
NAND2_X1 MEM_stage_inst_dmem_U3523 ( .A1(MEM_stage_inst_dmem_ram_2022), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n3381) );
NAND2_X1 MEM_stage_inst_dmem_U3522 ( .A1(MEM_stage_inst_dmem_ram_1606), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n3382) );
NAND2_X1 MEM_stage_inst_dmem_U3521 ( .A1(MEM_stage_inst_dmem_n3380), .A2(MEM_stage_inst_dmem_n3379), .ZN(MEM_stage_inst_dmem_n3384) );
NAND2_X1 MEM_stage_inst_dmem_U3520 ( .A1(MEM_stage_inst_dmem_ram_1798), .A2(MEM_stage_inst_dmem_n37), .ZN(MEM_stage_inst_dmem_n3379) );
NAND2_X1 MEM_stage_inst_dmem_U3519 ( .A1(MEM_stage_inst_dmem_ram_1430), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n3380) );
NAND2_X1 MEM_stage_inst_dmem_U3518 ( .A1(MEM_stage_inst_dmem_n3378), .A2(MEM_stage_inst_dmem_n3377), .ZN(MEM_stage_inst_dmem_n3394) );
NOR2_X1 MEM_stage_inst_dmem_U3517 ( .A1(MEM_stage_inst_dmem_n3376), .A2(MEM_stage_inst_dmem_n3375), .ZN(MEM_stage_inst_dmem_n3377) );
NAND2_X1 MEM_stage_inst_dmem_U3516 ( .A1(MEM_stage_inst_dmem_n3374), .A2(MEM_stage_inst_dmem_n3373), .ZN(MEM_stage_inst_dmem_n3375) );
NAND2_X1 MEM_stage_inst_dmem_U3515 ( .A1(MEM_stage_inst_dmem_ram_1046), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n3373) );
NAND2_X1 MEM_stage_inst_dmem_U3514 ( .A1(MEM_stage_inst_dmem_ram_1174), .A2(MEM_stage_inst_dmem_n5807), .ZN(MEM_stage_inst_dmem_n3374) );
NAND2_X1 MEM_stage_inst_dmem_U3513 ( .A1(MEM_stage_inst_dmem_n3372), .A2(MEM_stage_inst_dmem_n3371), .ZN(MEM_stage_inst_dmem_n3376) );
NAND2_X1 MEM_stage_inst_dmem_U3512 ( .A1(MEM_stage_inst_dmem_ram_1990), .A2(MEM_stage_inst_dmem_n4728), .ZN(MEM_stage_inst_dmem_n3371) );
NAND2_X1 MEM_stage_inst_dmem_U3511 ( .A1(MEM_stage_inst_dmem_ram_1542), .A2(MEM_stage_inst_dmem_n71), .ZN(MEM_stage_inst_dmem_n3372) );
NOR2_X1 MEM_stage_inst_dmem_U3510 ( .A1(MEM_stage_inst_dmem_n3370), .A2(MEM_stage_inst_dmem_n3369), .ZN(MEM_stage_inst_dmem_n3378) );
NAND2_X1 MEM_stage_inst_dmem_U3509 ( .A1(MEM_stage_inst_dmem_n3368), .A2(MEM_stage_inst_dmem_n3367), .ZN(MEM_stage_inst_dmem_n3369) );
NAND2_X1 MEM_stage_inst_dmem_U3508 ( .A1(MEM_stage_inst_dmem_ram_1750), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n3367) );
NAND2_X1 MEM_stage_inst_dmem_U3507 ( .A1(MEM_stage_inst_dmem_ram_1398), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n3368) );
NAND2_X1 MEM_stage_inst_dmem_U3506 ( .A1(MEM_stage_inst_dmem_n3366), .A2(MEM_stage_inst_dmem_n3365), .ZN(MEM_stage_inst_dmem_n3370) );
NAND2_X1 MEM_stage_inst_dmem_U3505 ( .A1(MEM_stage_inst_dmem_ram_1926), .A2(MEM_stage_inst_dmem_n72), .ZN(MEM_stage_inst_dmem_n3365) );
NAND2_X1 MEM_stage_inst_dmem_U3504 ( .A1(MEM_stage_inst_dmem_ram_1030), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n3366) );
NAND2_X1 MEM_stage_inst_dmem_U3503 ( .A1(MEM_stage_inst_dmem_n3364), .A2(MEM_stage_inst_dmem_n3363), .ZN(MEM_stage_inst_mem_read_data_5) );
NOR2_X1 MEM_stage_inst_dmem_U3502 ( .A1(MEM_stage_inst_dmem_n3362), .A2(MEM_stage_inst_dmem_n3361), .ZN(MEM_stage_inst_dmem_n3363) );
NOR2_X1 MEM_stage_inst_dmem_U3501 ( .A1(MEM_stage_inst_dmem_n3360), .A2(MEM_stage_inst_dmem_n8286), .ZN(MEM_stage_inst_dmem_n3361) );
NOR2_X1 MEM_stage_inst_dmem_U3500 ( .A1(MEM_stage_inst_dmem_n3359), .A2(MEM_stage_inst_dmem_n3358), .ZN(MEM_stage_inst_dmem_n3360) );
NAND2_X1 MEM_stage_inst_dmem_U3499 ( .A1(MEM_stage_inst_dmem_n3357), .A2(MEM_stage_inst_dmem_n3356), .ZN(MEM_stage_inst_dmem_n3358) );
NOR2_X1 MEM_stage_inst_dmem_U3498 ( .A1(MEM_stage_inst_dmem_n3355), .A2(MEM_stage_inst_dmem_n3354), .ZN(MEM_stage_inst_dmem_n3356) );
NAND2_X1 MEM_stage_inst_dmem_U3497 ( .A1(MEM_stage_inst_dmem_n3353), .A2(MEM_stage_inst_dmem_n3352), .ZN(MEM_stage_inst_dmem_n3354) );
NOR2_X1 MEM_stage_inst_dmem_U3496 ( .A1(MEM_stage_inst_dmem_n3351), .A2(MEM_stage_inst_dmem_n3350), .ZN(MEM_stage_inst_dmem_n3352) );
NAND2_X1 MEM_stage_inst_dmem_U3495 ( .A1(MEM_stage_inst_dmem_n3349), .A2(MEM_stage_inst_dmem_n3348), .ZN(MEM_stage_inst_dmem_n3350) );
NAND2_X1 MEM_stage_inst_dmem_U3494 ( .A1(MEM_stage_inst_dmem_ram_2949), .A2(MEM_stage_inst_dmem_n72), .ZN(MEM_stage_inst_dmem_n3348) );
NAND2_X1 MEM_stage_inst_dmem_U3493 ( .A1(MEM_stage_inst_dmem_ram_2165), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n3349) );
NAND2_X1 MEM_stage_inst_dmem_U3492 ( .A1(MEM_stage_inst_dmem_n3347), .A2(MEM_stage_inst_dmem_n3346), .ZN(MEM_stage_inst_dmem_n3351) );
NAND2_X1 MEM_stage_inst_dmem_U3491 ( .A1(MEM_stage_inst_dmem_ram_2101), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n3346) );
NAND2_X1 MEM_stage_inst_dmem_U3490 ( .A1(MEM_stage_inst_dmem_ram_2325), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n3347) );
NOR2_X1 MEM_stage_inst_dmem_U3489 ( .A1(MEM_stage_inst_dmem_n3345), .A2(MEM_stage_inst_dmem_n3344), .ZN(MEM_stage_inst_dmem_n3353) );
NAND2_X1 MEM_stage_inst_dmem_U3488 ( .A1(MEM_stage_inst_dmem_n3343), .A2(MEM_stage_inst_dmem_n3342), .ZN(MEM_stage_inst_dmem_n3344) );
NAND2_X1 MEM_stage_inst_dmem_U3487 ( .A1(MEM_stage_inst_dmem_ram_2933), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n3342) );
NAND2_X1 MEM_stage_inst_dmem_U3486 ( .A1(MEM_stage_inst_dmem_ram_2069), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n3343) );
NAND2_X1 MEM_stage_inst_dmem_U3485 ( .A1(MEM_stage_inst_dmem_n3341), .A2(MEM_stage_inst_dmem_n3340), .ZN(MEM_stage_inst_dmem_n3345) );
NAND2_X1 MEM_stage_inst_dmem_U3484 ( .A1(MEM_stage_inst_dmem_ram_2549), .A2(MEM_stage_inst_dmem_n8535), .ZN(MEM_stage_inst_dmem_n3340) );
NAND2_X1 MEM_stage_inst_dmem_U3483 ( .A1(MEM_stage_inst_dmem_ram_3045), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n3341) );
NAND2_X1 MEM_stage_inst_dmem_U3482 ( .A1(MEM_stage_inst_dmem_n3339), .A2(MEM_stage_inst_dmem_n3338), .ZN(MEM_stage_inst_dmem_n3355) );
NOR2_X1 MEM_stage_inst_dmem_U3481 ( .A1(MEM_stage_inst_dmem_n3337), .A2(MEM_stage_inst_dmem_n3336), .ZN(MEM_stage_inst_dmem_n3338) );
NAND2_X1 MEM_stage_inst_dmem_U3480 ( .A1(MEM_stage_inst_dmem_n3335), .A2(MEM_stage_inst_dmem_n3334), .ZN(MEM_stage_inst_dmem_n3336) );
NAND2_X1 MEM_stage_inst_dmem_U3479 ( .A1(MEM_stage_inst_dmem_ram_2405), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n3334) );
NAND2_X1 MEM_stage_inst_dmem_U3478 ( .A1(MEM_stage_inst_dmem_ram_3013), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n3335) );
NAND2_X1 MEM_stage_inst_dmem_U3477 ( .A1(MEM_stage_inst_dmem_n3333), .A2(MEM_stage_inst_dmem_n3332), .ZN(MEM_stage_inst_dmem_n3337) );
NAND2_X1 MEM_stage_inst_dmem_U3476 ( .A1(MEM_stage_inst_dmem_ram_2885), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n3332) );
NAND2_X1 MEM_stage_inst_dmem_U3475 ( .A1(MEM_stage_inst_dmem_ram_2453), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n3333) );
NOR2_X1 MEM_stage_inst_dmem_U3474 ( .A1(MEM_stage_inst_dmem_n3331), .A2(MEM_stage_inst_dmem_n3330), .ZN(MEM_stage_inst_dmem_n3339) );
NAND2_X1 MEM_stage_inst_dmem_U3473 ( .A1(MEM_stage_inst_dmem_n3329), .A2(MEM_stage_inst_dmem_n3328), .ZN(MEM_stage_inst_dmem_n3330) );
NAND2_X1 MEM_stage_inst_dmem_U3472 ( .A1(MEM_stage_inst_dmem_ram_2293), .A2(MEM_stage_inst_dmem_n39), .ZN(MEM_stage_inst_dmem_n3328) );
NAND2_X1 MEM_stage_inst_dmem_U3471 ( .A1(MEM_stage_inst_dmem_ram_2869), .A2(MEM_stage_inst_dmem_n46), .ZN(MEM_stage_inst_dmem_n3329) );
NAND2_X1 MEM_stage_inst_dmem_U3470 ( .A1(MEM_stage_inst_dmem_n3327), .A2(MEM_stage_inst_dmem_n3326), .ZN(MEM_stage_inst_dmem_n3331) );
NAND2_X1 MEM_stage_inst_dmem_U3469 ( .A1(MEM_stage_inst_dmem_ram_2901), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n3326) );
NAND2_X1 MEM_stage_inst_dmem_U3468 ( .A1(MEM_stage_inst_dmem_ram_2517), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n3327) );
NOR2_X1 MEM_stage_inst_dmem_U3467 ( .A1(MEM_stage_inst_dmem_n3325), .A2(MEM_stage_inst_dmem_n3324), .ZN(MEM_stage_inst_dmem_n3357) );
NAND2_X1 MEM_stage_inst_dmem_U3466 ( .A1(MEM_stage_inst_dmem_n3323), .A2(MEM_stage_inst_dmem_n3322), .ZN(MEM_stage_inst_dmem_n3324) );
NOR2_X1 MEM_stage_inst_dmem_U3465 ( .A1(MEM_stage_inst_dmem_n3321), .A2(MEM_stage_inst_dmem_n3320), .ZN(MEM_stage_inst_dmem_n3322) );
NAND2_X1 MEM_stage_inst_dmem_U3464 ( .A1(MEM_stage_inst_dmem_n3319), .A2(MEM_stage_inst_dmem_n3318), .ZN(MEM_stage_inst_dmem_n3320) );
NAND2_X1 MEM_stage_inst_dmem_U3463 ( .A1(MEM_stage_inst_dmem_ram_2917), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n3318) );
NAND2_X1 MEM_stage_inst_dmem_U3462 ( .A1(MEM_stage_inst_dmem_ram_2357), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n3319) );
NAND2_X1 MEM_stage_inst_dmem_U3461 ( .A1(MEM_stage_inst_dmem_n3317), .A2(MEM_stage_inst_dmem_n3316), .ZN(MEM_stage_inst_dmem_n3321) );
NAND2_X1 MEM_stage_inst_dmem_U3460 ( .A1(MEM_stage_inst_dmem_ram_2757), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n3316) );
NAND2_X1 MEM_stage_inst_dmem_U3459 ( .A1(MEM_stage_inst_dmem_ram_2085), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n3317) );
NOR2_X1 MEM_stage_inst_dmem_U3458 ( .A1(MEM_stage_inst_dmem_n3315), .A2(MEM_stage_inst_dmem_n3314), .ZN(MEM_stage_inst_dmem_n3323) );
NAND2_X1 MEM_stage_inst_dmem_U3457 ( .A1(MEM_stage_inst_dmem_n3313), .A2(MEM_stage_inst_dmem_n3312), .ZN(MEM_stage_inst_dmem_n3314) );
NAND2_X1 MEM_stage_inst_dmem_U3456 ( .A1(MEM_stage_inst_dmem_ram_3061), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n3312) );
NAND2_X1 MEM_stage_inst_dmem_U3455 ( .A1(MEM_stage_inst_dmem_ram_2341), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n3313) );
NAND2_X1 MEM_stage_inst_dmem_U3454 ( .A1(MEM_stage_inst_dmem_n3311), .A2(MEM_stage_inst_dmem_n3310), .ZN(MEM_stage_inst_dmem_n3315) );
NAND2_X1 MEM_stage_inst_dmem_U3453 ( .A1(MEM_stage_inst_dmem_ram_3029), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n3310) );
NAND2_X1 MEM_stage_inst_dmem_U3452 ( .A1(MEM_stage_inst_dmem_ram_2437), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n3311) );
NAND2_X1 MEM_stage_inst_dmem_U3451 ( .A1(MEM_stage_inst_dmem_n3309), .A2(MEM_stage_inst_dmem_n3308), .ZN(MEM_stage_inst_dmem_n3325) );
NOR2_X1 MEM_stage_inst_dmem_U3450 ( .A1(MEM_stage_inst_dmem_n3307), .A2(MEM_stage_inst_dmem_n3306), .ZN(MEM_stage_inst_dmem_n3308) );
NAND2_X1 MEM_stage_inst_dmem_U3449 ( .A1(MEM_stage_inst_dmem_n3305), .A2(MEM_stage_inst_dmem_n3304), .ZN(MEM_stage_inst_dmem_n3306) );
NAND2_X1 MEM_stage_inst_dmem_U3448 ( .A1(MEM_stage_inst_dmem_ram_2245), .A2(MEM_stage_inst_dmem_n36), .ZN(MEM_stage_inst_dmem_n3304) );
NAND2_X1 MEM_stage_inst_dmem_U3447 ( .A1(MEM_stage_inst_dmem_ram_2501), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n3305) );
NAND2_X1 MEM_stage_inst_dmem_U3446 ( .A1(MEM_stage_inst_dmem_n3303), .A2(MEM_stage_inst_dmem_n3302), .ZN(MEM_stage_inst_dmem_n3307) );
NAND2_X1 MEM_stage_inst_dmem_U3445 ( .A1(MEM_stage_inst_dmem_ram_2821), .A2(MEM_stage_inst_dmem_n37), .ZN(MEM_stage_inst_dmem_n3302) );
NAND2_X1 MEM_stage_inst_dmem_U3444 ( .A1(MEM_stage_inst_dmem_ram_2469), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n3303) );
NOR2_X1 MEM_stage_inst_dmem_U3443 ( .A1(MEM_stage_inst_dmem_n3301), .A2(MEM_stage_inst_dmem_n3300), .ZN(MEM_stage_inst_dmem_n3309) );
NAND2_X1 MEM_stage_inst_dmem_U3442 ( .A1(MEM_stage_inst_dmem_n3299), .A2(MEM_stage_inst_dmem_n3298), .ZN(MEM_stage_inst_dmem_n3300) );
NAND2_X1 MEM_stage_inst_dmem_U3441 ( .A1(MEM_stage_inst_dmem_ram_2805), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n3298) );
NAND2_X1 MEM_stage_inst_dmem_U3440 ( .A1(MEM_stage_inst_dmem_ram_2741), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n3299) );
NAND2_X1 MEM_stage_inst_dmem_U3439 ( .A1(MEM_stage_inst_dmem_n3297), .A2(MEM_stage_inst_dmem_n3296), .ZN(MEM_stage_inst_dmem_n3301) );
NAND2_X1 MEM_stage_inst_dmem_U3438 ( .A1(MEM_stage_inst_dmem_ram_2309), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n3296) );
NAND2_X1 MEM_stage_inst_dmem_U3437 ( .A1(MEM_stage_inst_dmem_ram_2789), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n3297) );
NAND2_X1 MEM_stage_inst_dmem_U3436 ( .A1(MEM_stage_inst_dmem_n3295), .A2(MEM_stage_inst_dmem_n3294), .ZN(MEM_stage_inst_dmem_n3359) );
NOR2_X1 MEM_stage_inst_dmem_U3435 ( .A1(MEM_stage_inst_dmem_n3293), .A2(MEM_stage_inst_dmem_n3292), .ZN(MEM_stage_inst_dmem_n3294) );
NAND2_X1 MEM_stage_inst_dmem_U3434 ( .A1(MEM_stage_inst_dmem_n3291), .A2(MEM_stage_inst_dmem_n3290), .ZN(MEM_stage_inst_dmem_n3292) );
NOR2_X1 MEM_stage_inst_dmem_U3433 ( .A1(MEM_stage_inst_dmem_n3289), .A2(MEM_stage_inst_dmem_n3288), .ZN(MEM_stage_inst_dmem_n3290) );
NAND2_X1 MEM_stage_inst_dmem_U3432 ( .A1(MEM_stage_inst_dmem_n3287), .A2(MEM_stage_inst_dmem_n3286), .ZN(MEM_stage_inst_dmem_n3288) );
NAND2_X1 MEM_stage_inst_dmem_U3431 ( .A1(MEM_stage_inst_dmem_ram_2613), .A2(MEM_stage_inst_dmem_n41), .ZN(MEM_stage_inst_dmem_n3286) );
NAND2_X1 MEM_stage_inst_dmem_U3430 ( .A1(MEM_stage_inst_dmem_ram_2181), .A2(MEM_stage_inst_dmem_n61), .ZN(MEM_stage_inst_dmem_n3287) );
NAND2_X1 MEM_stage_inst_dmem_U3429 ( .A1(MEM_stage_inst_dmem_n3285), .A2(MEM_stage_inst_dmem_n3284), .ZN(MEM_stage_inst_dmem_n3289) );
NAND2_X1 MEM_stage_inst_dmem_U3428 ( .A1(MEM_stage_inst_dmem_ram_2965), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n3284) );
NAND2_X1 MEM_stage_inst_dmem_U3427 ( .A1(MEM_stage_inst_dmem_ram_2565), .A2(MEM_stage_inst_dmem_n71), .ZN(MEM_stage_inst_dmem_n3285) );
NOR2_X1 MEM_stage_inst_dmem_U3426 ( .A1(MEM_stage_inst_dmem_n3283), .A2(MEM_stage_inst_dmem_n3282), .ZN(MEM_stage_inst_dmem_n3291) );
NAND2_X1 MEM_stage_inst_dmem_U3425 ( .A1(MEM_stage_inst_dmem_n3281), .A2(MEM_stage_inst_dmem_n3280), .ZN(MEM_stage_inst_dmem_n3282) );
NAND2_X1 MEM_stage_inst_dmem_U3424 ( .A1(MEM_stage_inst_dmem_ram_2197), .A2(MEM_stage_inst_dmem_n44), .ZN(MEM_stage_inst_dmem_n3280) );
NAND2_X1 MEM_stage_inst_dmem_U3423 ( .A1(MEM_stage_inst_dmem_ram_2213), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n3281) );
NAND2_X1 MEM_stage_inst_dmem_U3422 ( .A1(MEM_stage_inst_dmem_n3279), .A2(MEM_stage_inst_dmem_n3278), .ZN(MEM_stage_inst_dmem_n3283) );
NAND2_X1 MEM_stage_inst_dmem_U3421 ( .A1(MEM_stage_inst_dmem_ram_2533), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n3278) );
NAND2_X1 MEM_stage_inst_dmem_U3420 ( .A1(MEM_stage_inst_dmem_ram_2661), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n3279) );
NAND2_X1 MEM_stage_inst_dmem_U3419 ( .A1(MEM_stage_inst_dmem_n3277), .A2(MEM_stage_inst_dmem_n3276), .ZN(MEM_stage_inst_dmem_n3293) );
NOR2_X1 MEM_stage_inst_dmem_U3418 ( .A1(MEM_stage_inst_dmem_n3275), .A2(MEM_stage_inst_dmem_n3274), .ZN(MEM_stage_inst_dmem_n3276) );
NAND2_X1 MEM_stage_inst_dmem_U3417 ( .A1(MEM_stage_inst_dmem_n3273), .A2(MEM_stage_inst_dmem_n3272), .ZN(MEM_stage_inst_dmem_n3274) );
NAND2_X1 MEM_stage_inst_dmem_U3416 ( .A1(MEM_stage_inst_dmem_ram_2277), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n3272) );
NAND2_X1 MEM_stage_inst_dmem_U3415 ( .A1(MEM_stage_inst_dmem_ram_2421), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n3273) );
NAND2_X1 MEM_stage_inst_dmem_U3414 ( .A1(MEM_stage_inst_dmem_n3271), .A2(MEM_stage_inst_dmem_n3270), .ZN(MEM_stage_inst_dmem_n3275) );
NAND2_X1 MEM_stage_inst_dmem_U3413 ( .A1(MEM_stage_inst_dmem_ram_2853), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n3270) );
NAND2_X1 MEM_stage_inst_dmem_U3412 ( .A1(MEM_stage_inst_dmem_ram_2133), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n3271) );
NOR2_X1 MEM_stage_inst_dmem_U3411 ( .A1(MEM_stage_inst_dmem_n3269), .A2(MEM_stage_inst_dmem_n3268), .ZN(MEM_stage_inst_dmem_n3277) );
NAND2_X1 MEM_stage_inst_dmem_U3410 ( .A1(MEM_stage_inst_dmem_n3267), .A2(MEM_stage_inst_dmem_n3266), .ZN(MEM_stage_inst_dmem_n3268) );
NAND2_X1 MEM_stage_inst_dmem_U3409 ( .A1(MEM_stage_inst_dmem_ram_2117), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n3266) );
NAND2_X1 MEM_stage_inst_dmem_U3408 ( .A1(MEM_stage_inst_dmem_ram_2677), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n3267) );
NAND2_X1 MEM_stage_inst_dmem_U3407 ( .A1(MEM_stage_inst_dmem_n3265), .A2(MEM_stage_inst_dmem_n3264), .ZN(MEM_stage_inst_dmem_n3269) );
NAND2_X1 MEM_stage_inst_dmem_U3406 ( .A1(MEM_stage_inst_dmem_ram_2389), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n3264) );
NAND2_X1 MEM_stage_inst_dmem_U3405 ( .A1(MEM_stage_inst_dmem_ram_2645), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n3265) );
NOR2_X1 MEM_stage_inst_dmem_U3404 ( .A1(MEM_stage_inst_dmem_n3263), .A2(MEM_stage_inst_dmem_n3262), .ZN(MEM_stage_inst_dmem_n3295) );
NAND2_X1 MEM_stage_inst_dmem_U3403 ( .A1(MEM_stage_inst_dmem_n3261), .A2(MEM_stage_inst_dmem_n3260), .ZN(MEM_stage_inst_dmem_n3262) );
NOR2_X1 MEM_stage_inst_dmem_U3402 ( .A1(MEM_stage_inst_dmem_n3259), .A2(MEM_stage_inst_dmem_n3258), .ZN(MEM_stage_inst_dmem_n3260) );
NAND2_X1 MEM_stage_inst_dmem_U3401 ( .A1(MEM_stage_inst_dmem_n3257), .A2(MEM_stage_inst_dmem_n3256), .ZN(MEM_stage_inst_dmem_n3258) );
NAND2_X1 MEM_stage_inst_dmem_U3400 ( .A1(MEM_stage_inst_dmem_ram_2981), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n3256) );
NAND2_X1 MEM_stage_inst_dmem_U3399 ( .A1(MEM_stage_inst_dmem_ram_2709), .A2(MEM_stage_inst_dmem_n3076), .ZN(MEM_stage_inst_dmem_n3257) );
NAND2_X1 MEM_stage_inst_dmem_U3398 ( .A1(MEM_stage_inst_dmem_n3255), .A2(MEM_stage_inst_dmem_n3254), .ZN(MEM_stage_inst_dmem_n3259) );
NAND2_X1 MEM_stage_inst_dmem_U3397 ( .A1(MEM_stage_inst_dmem_ram_2053), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n3254) );
NAND2_X1 MEM_stage_inst_dmem_U3396 ( .A1(MEM_stage_inst_dmem_ram_2773), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n3255) );
NOR2_X1 MEM_stage_inst_dmem_U3395 ( .A1(MEM_stage_inst_dmem_n3253), .A2(MEM_stage_inst_dmem_n3252), .ZN(MEM_stage_inst_dmem_n3261) );
NAND2_X1 MEM_stage_inst_dmem_U3394 ( .A1(MEM_stage_inst_dmem_n3251), .A2(MEM_stage_inst_dmem_n3250), .ZN(MEM_stage_inst_dmem_n3252) );
NAND2_X1 MEM_stage_inst_dmem_U3393 ( .A1(MEM_stage_inst_dmem_ram_2997), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n3250) );
NAND2_X1 MEM_stage_inst_dmem_U3392 ( .A1(MEM_stage_inst_dmem_ram_2261), .A2(MEM_stage_inst_dmem_n51), .ZN(MEM_stage_inst_dmem_n3251) );
NAND2_X1 MEM_stage_inst_dmem_U3391 ( .A1(MEM_stage_inst_dmem_n3249), .A2(MEM_stage_inst_dmem_n3248), .ZN(MEM_stage_inst_dmem_n3253) );
NAND2_X1 MEM_stage_inst_dmem_U3390 ( .A1(MEM_stage_inst_dmem_ram_2485), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n3248) );
NAND2_X1 MEM_stage_inst_dmem_U3389 ( .A1(MEM_stage_inst_dmem_ram_2837), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n3249) );
NAND2_X1 MEM_stage_inst_dmem_U3388 ( .A1(MEM_stage_inst_dmem_n3247), .A2(MEM_stage_inst_dmem_n3246), .ZN(MEM_stage_inst_dmem_n3263) );
NOR2_X1 MEM_stage_inst_dmem_U3387 ( .A1(MEM_stage_inst_dmem_n3245), .A2(MEM_stage_inst_dmem_n3244), .ZN(MEM_stage_inst_dmem_n3246) );
NAND2_X1 MEM_stage_inst_dmem_U3386 ( .A1(MEM_stage_inst_dmem_n3243), .A2(MEM_stage_inst_dmem_n3242), .ZN(MEM_stage_inst_dmem_n3244) );
NAND2_X1 MEM_stage_inst_dmem_U3385 ( .A1(MEM_stage_inst_dmem_ram_2693), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n3242) );
NAND2_X1 MEM_stage_inst_dmem_U3384 ( .A1(MEM_stage_inst_dmem_ram_2581), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n3243) );
NAND2_X1 MEM_stage_inst_dmem_U3383 ( .A1(MEM_stage_inst_dmem_n3241), .A2(MEM_stage_inst_dmem_n3240), .ZN(MEM_stage_inst_dmem_n3245) );
NAND2_X1 MEM_stage_inst_dmem_U3382 ( .A1(MEM_stage_inst_dmem_ram_2725), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n3240) );
NAND2_X1 MEM_stage_inst_dmem_U3381 ( .A1(MEM_stage_inst_dmem_ram_2629), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n3241) );
NOR2_X1 MEM_stage_inst_dmem_U3380 ( .A1(MEM_stage_inst_dmem_n3239), .A2(MEM_stage_inst_dmem_n3238), .ZN(MEM_stage_inst_dmem_n3247) );
NAND2_X1 MEM_stage_inst_dmem_U3379 ( .A1(MEM_stage_inst_dmem_n3237), .A2(MEM_stage_inst_dmem_n3236), .ZN(MEM_stage_inst_dmem_n3238) );
NAND2_X1 MEM_stage_inst_dmem_U3378 ( .A1(MEM_stage_inst_dmem_ram_2373), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n3236) );
NAND2_X1 MEM_stage_inst_dmem_U3377 ( .A1(MEM_stage_inst_dmem_ram_2149), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n3237) );
NAND2_X1 MEM_stage_inst_dmem_U3376 ( .A1(MEM_stage_inst_dmem_n3235), .A2(MEM_stage_inst_dmem_n3234), .ZN(MEM_stage_inst_dmem_n3239) );
NAND2_X1 MEM_stage_inst_dmem_U3375 ( .A1(MEM_stage_inst_dmem_ram_2597), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n3234) );
NAND2_X1 MEM_stage_inst_dmem_U3374 ( .A1(MEM_stage_inst_dmem_ram_2229), .A2(MEM_stage_inst_dmem_n55), .ZN(MEM_stage_inst_dmem_n3235) );
NOR2_X1 MEM_stage_inst_dmem_U3373 ( .A1(MEM_stage_inst_dmem_n3233), .A2(MEM_stage_inst_dmem_n8152), .ZN(MEM_stage_inst_dmem_n3362) );
NOR2_X1 MEM_stage_inst_dmem_U3372 ( .A1(MEM_stage_inst_dmem_n3232), .A2(MEM_stage_inst_dmem_n3231), .ZN(MEM_stage_inst_dmem_n3233) );
NAND2_X1 MEM_stage_inst_dmem_U3371 ( .A1(MEM_stage_inst_dmem_n3230), .A2(MEM_stage_inst_dmem_n3229), .ZN(MEM_stage_inst_dmem_n3231) );
NOR2_X1 MEM_stage_inst_dmem_U3370 ( .A1(MEM_stage_inst_dmem_n3228), .A2(MEM_stage_inst_dmem_n3227), .ZN(MEM_stage_inst_dmem_n3229) );
NAND2_X1 MEM_stage_inst_dmem_U3369 ( .A1(MEM_stage_inst_dmem_n3226), .A2(MEM_stage_inst_dmem_n3225), .ZN(MEM_stage_inst_dmem_n3227) );
NOR2_X1 MEM_stage_inst_dmem_U3368 ( .A1(MEM_stage_inst_dmem_n3224), .A2(MEM_stage_inst_dmem_n3223), .ZN(MEM_stage_inst_dmem_n3225) );
NAND2_X1 MEM_stage_inst_dmem_U3367 ( .A1(MEM_stage_inst_dmem_n3222), .A2(MEM_stage_inst_dmem_n3221), .ZN(MEM_stage_inst_dmem_n3223) );
NAND2_X1 MEM_stage_inst_dmem_U3366 ( .A1(MEM_stage_inst_dmem_ram_1141), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n3221) );
NAND2_X1 MEM_stage_inst_dmem_U3365 ( .A1(MEM_stage_inst_dmem_ram_1237), .A2(MEM_stage_inst_dmem_n51), .ZN(MEM_stage_inst_dmem_n3222) );
NAND2_X1 MEM_stage_inst_dmem_U3364 ( .A1(MEM_stage_inst_dmem_n3219), .A2(MEM_stage_inst_dmem_n3218), .ZN(MEM_stage_inst_dmem_n3224) );
NAND2_X1 MEM_stage_inst_dmem_U3363 ( .A1(MEM_stage_inst_dmem_ram_1381), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n3218) );
NAND2_X1 MEM_stage_inst_dmem_U3362 ( .A1(MEM_stage_inst_dmem_ram_1365), .A2(MEM_stage_inst_dmem_n3216), .ZN(MEM_stage_inst_dmem_n3219) );
NOR2_X1 MEM_stage_inst_dmem_U3361 ( .A1(MEM_stage_inst_dmem_n3215), .A2(MEM_stage_inst_dmem_n3214), .ZN(MEM_stage_inst_dmem_n3226) );
NAND2_X1 MEM_stage_inst_dmem_U3360 ( .A1(MEM_stage_inst_dmem_n3213), .A2(MEM_stage_inst_dmem_n3212), .ZN(MEM_stage_inst_dmem_n3214) );
NAND2_X1 MEM_stage_inst_dmem_U3359 ( .A1(MEM_stage_inst_dmem_ram_1573), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n3212) );
NAND2_X1 MEM_stage_inst_dmem_U3358 ( .A1(MEM_stage_inst_dmem_ram_1109), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n3213) );
NAND2_X1 MEM_stage_inst_dmem_U3357 ( .A1(MEM_stage_inst_dmem_n3211), .A2(MEM_stage_inst_dmem_n3210), .ZN(MEM_stage_inst_dmem_n3215) );
NAND2_X1 MEM_stage_inst_dmem_U3356 ( .A1(MEM_stage_inst_dmem_ram_1269), .A2(MEM_stage_inst_dmem_n39), .ZN(MEM_stage_inst_dmem_n3210) );
NAND2_X1 MEM_stage_inst_dmem_U3355 ( .A1(MEM_stage_inst_dmem_ram_1317), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n3211) );
NAND2_X1 MEM_stage_inst_dmem_U3354 ( .A1(MEM_stage_inst_dmem_n3208), .A2(MEM_stage_inst_dmem_n3207), .ZN(MEM_stage_inst_dmem_n3228) );
NOR2_X1 MEM_stage_inst_dmem_U3353 ( .A1(MEM_stage_inst_dmem_n3206), .A2(MEM_stage_inst_dmem_n3205), .ZN(MEM_stage_inst_dmem_n3207) );
NAND2_X1 MEM_stage_inst_dmem_U3352 ( .A1(MEM_stage_inst_dmem_n3204), .A2(MEM_stage_inst_dmem_n3203), .ZN(MEM_stage_inst_dmem_n3205) );
NAND2_X1 MEM_stage_inst_dmem_U3351 ( .A1(MEM_stage_inst_dmem_ram_1781), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n3203) );
NAND2_X1 MEM_stage_inst_dmem_U3350 ( .A1(MEM_stage_inst_dmem_ram_1605), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n3204) );
NAND2_X1 MEM_stage_inst_dmem_U3349 ( .A1(MEM_stage_inst_dmem_n3201), .A2(MEM_stage_inst_dmem_n3200), .ZN(MEM_stage_inst_dmem_n3206) );
NAND2_X1 MEM_stage_inst_dmem_U3348 ( .A1(MEM_stage_inst_dmem_ram_2037), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n3200) );
NAND2_X1 MEM_stage_inst_dmem_U3347 ( .A1(MEM_stage_inst_dmem_ram_1957), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n3201) );
NOR2_X1 MEM_stage_inst_dmem_U3346 ( .A1(MEM_stage_inst_dmem_n3198), .A2(MEM_stage_inst_dmem_n3197), .ZN(MEM_stage_inst_dmem_n3208) );
NAND2_X1 MEM_stage_inst_dmem_U3345 ( .A1(MEM_stage_inst_dmem_n3196), .A2(MEM_stage_inst_dmem_n3195), .ZN(MEM_stage_inst_dmem_n3197) );
NAND2_X1 MEM_stage_inst_dmem_U3344 ( .A1(MEM_stage_inst_dmem_ram_1797), .A2(MEM_stage_inst_dmem_n37), .ZN(MEM_stage_inst_dmem_n3195) );
NAND2_X1 MEM_stage_inst_dmem_U3343 ( .A1(MEM_stage_inst_dmem_ram_1413), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n3196) );
NAND2_X1 MEM_stage_inst_dmem_U3342 ( .A1(MEM_stage_inst_dmem_n3194), .A2(MEM_stage_inst_dmem_n3193), .ZN(MEM_stage_inst_dmem_n3198) );
NAND2_X1 MEM_stage_inst_dmem_U3341 ( .A1(MEM_stage_inst_dmem_ram_1733), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n3193) );
NAND2_X1 MEM_stage_inst_dmem_U3340 ( .A1(MEM_stage_inst_dmem_ram_1813), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n3194) );
NOR2_X1 MEM_stage_inst_dmem_U3339 ( .A1(MEM_stage_inst_dmem_n3190), .A2(MEM_stage_inst_dmem_n3189), .ZN(MEM_stage_inst_dmem_n3230) );
NAND2_X1 MEM_stage_inst_dmem_U3338 ( .A1(MEM_stage_inst_dmem_n3188), .A2(MEM_stage_inst_dmem_n3187), .ZN(MEM_stage_inst_dmem_n3189) );
NOR2_X1 MEM_stage_inst_dmem_U3337 ( .A1(MEM_stage_inst_dmem_n3186), .A2(MEM_stage_inst_dmem_n3185), .ZN(MEM_stage_inst_dmem_n3187) );
NAND2_X1 MEM_stage_inst_dmem_U3336 ( .A1(MEM_stage_inst_dmem_n3184), .A2(MEM_stage_inst_dmem_n3183), .ZN(MEM_stage_inst_dmem_n3185) );
NAND2_X1 MEM_stage_inst_dmem_U3335 ( .A1(MEM_stage_inst_dmem_ram_1509), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n3183) );
NAND2_X1 MEM_stage_inst_dmem_U3334 ( .A1(MEM_stage_inst_dmem_ram_1541), .A2(MEM_stage_inst_dmem_n71), .ZN(MEM_stage_inst_dmem_n3184) );
NAND2_X1 MEM_stage_inst_dmem_U3333 ( .A1(MEM_stage_inst_dmem_n3181), .A2(MEM_stage_inst_dmem_n3180), .ZN(MEM_stage_inst_dmem_n3186) );
NAND2_X1 MEM_stage_inst_dmem_U3332 ( .A1(MEM_stage_inst_dmem_ram_1173), .A2(MEM_stage_inst_dmem_n44), .ZN(MEM_stage_inst_dmem_n3180) );
NAND2_X1 MEM_stage_inst_dmem_U3331 ( .A1(MEM_stage_inst_dmem_ram_1125), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n3181) );
NOR2_X1 MEM_stage_inst_dmem_U3330 ( .A1(MEM_stage_inst_dmem_n3178), .A2(MEM_stage_inst_dmem_n3177), .ZN(MEM_stage_inst_dmem_n3188) );
NAND2_X1 MEM_stage_inst_dmem_U3329 ( .A1(MEM_stage_inst_dmem_n3176), .A2(MEM_stage_inst_dmem_n3175), .ZN(MEM_stage_inst_dmem_n3177) );
NAND2_X1 MEM_stage_inst_dmem_U3328 ( .A1(MEM_stage_inst_dmem_ram_1493), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n3175) );
NAND2_X1 MEM_stage_inst_dmem_U3327 ( .A1(MEM_stage_inst_dmem_ram_1477), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n3176) );
NAND2_X1 MEM_stage_inst_dmem_U3326 ( .A1(MEM_stage_inst_dmem_n3172), .A2(MEM_stage_inst_dmem_n3171), .ZN(MEM_stage_inst_dmem_n3178) );
NAND2_X1 MEM_stage_inst_dmem_U3325 ( .A1(MEM_stage_inst_dmem_ram_1525), .A2(MEM_stage_inst_dmem_n64), .ZN(MEM_stage_inst_dmem_n3171) );
NAND2_X1 MEM_stage_inst_dmem_U3324 ( .A1(MEM_stage_inst_dmem_ram_1397), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n3172) );
NAND2_X1 MEM_stage_inst_dmem_U3323 ( .A1(MEM_stage_inst_dmem_n3169), .A2(MEM_stage_inst_dmem_n3168), .ZN(MEM_stage_inst_dmem_n3190) );
NOR2_X1 MEM_stage_inst_dmem_U3322 ( .A1(MEM_stage_inst_dmem_n3167), .A2(MEM_stage_inst_dmem_n3166), .ZN(MEM_stage_inst_dmem_n3168) );
NAND2_X1 MEM_stage_inst_dmem_U3321 ( .A1(MEM_stage_inst_dmem_n3165), .A2(MEM_stage_inst_dmem_n3164), .ZN(MEM_stage_inst_dmem_n3166) );
NAND2_X1 MEM_stage_inst_dmem_U3320 ( .A1(MEM_stage_inst_dmem_ram_1973), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n3164) );
NAND2_X1 MEM_stage_inst_dmem_U3319 ( .A1(MEM_stage_inst_dmem_ram_1045), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n3165) );
NAND2_X1 MEM_stage_inst_dmem_U3318 ( .A1(MEM_stage_inst_dmem_n3162), .A2(MEM_stage_inst_dmem_n3161), .ZN(MEM_stage_inst_dmem_n3167) );
NAND2_X1 MEM_stage_inst_dmem_U3317 ( .A1(MEM_stage_inst_dmem_ram_1429), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n3161) );
NAND2_X1 MEM_stage_inst_dmem_U3316 ( .A1(MEM_stage_inst_dmem_ram_1557), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n3162) );
NOR2_X1 MEM_stage_inst_dmem_U3315 ( .A1(MEM_stage_inst_dmem_n3159), .A2(MEM_stage_inst_dmem_n3158), .ZN(MEM_stage_inst_dmem_n3169) );
NAND2_X1 MEM_stage_inst_dmem_U3314 ( .A1(MEM_stage_inst_dmem_n3157), .A2(MEM_stage_inst_dmem_n3156), .ZN(MEM_stage_inst_dmem_n3158) );
NAND2_X1 MEM_stage_inst_dmem_U3313 ( .A1(MEM_stage_inst_dmem_ram_1989), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n3156) );
NAND2_X1 MEM_stage_inst_dmem_U3312 ( .A1(MEM_stage_inst_dmem_ram_1701), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n3157) );
NAND2_X1 MEM_stage_inst_dmem_U3311 ( .A1(MEM_stage_inst_dmem_n3154), .A2(MEM_stage_inst_dmem_n3153), .ZN(MEM_stage_inst_dmem_n3159) );
NAND2_X1 MEM_stage_inst_dmem_U3310 ( .A1(MEM_stage_inst_dmem_ram_1253), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n3153) );
NAND2_X1 MEM_stage_inst_dmem_U3309 ( .A1(MEM_stage_inst_dmem_ram_1717), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n3154) );
NAND2_X1 MEM_stage_inst_dmem_U3308 ( .A1(MEM_stage_inst_dmem_n3151), .A2(MEM_stage_inst_dmem_n3150), .ZN(MEM_stage_inst_dmem_n3232) );
NOR2_X1 MEM_stage_inst_dmem_U3307 ( .A1(MEM_stage_inst_dmem_n3149), .A2(MEM_stage_inst_dmem_n3148), .ZN(MEM_stage_inst_dmem_n3150) );
NAND2_X1 MEM_stage_inst_dmem_U3306 ( .A1(MEM_stage_inst_dmem_n3147), .A2(MEM_stage_inst_dmem_n3146), .ZN(MEM_stage_inst_dmem_n3148) );
NOR2_X1 MEM_stage_inst_dmem_U3305 ( .A1(MEM_stage_inst_dmem_n3145), .A2(MEM_stage_inst_dmem_n3144), .ZN(MEM_stage_inst_dmem_n3146) );
NAND2_X1 MEM_stage_inst_dmem_U3304 ( .A1(MEM_stage_inst_dmem_n3143), .A2(MEM_stage_inst_dmem_n3142), .ZN(MEM_stage_inst_dmem_n3144) );
NAND2_X1 MEM_stage_inst_dmem_U3303 ( .A1(MEM_stage_inst_dmem_ram_1877), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n3142) );
NAND2_X1 MEM_stage_inst_dmem_U3302 ( .A1(MEM_stage_inst_dmem_ram_1621), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n3143) );
NAND2_X1 MEM_stage_inst_dmem_U3301 ( .A1(MEM_stage_inst_dmem_n3139), .A2(MEM_stage_inst_dmem_n3138), .ZN(MEM_stage_inst_dmem_n3145) );
NAND2_X1 MEM_stage_inst_dmem_U3300 ( .A1(MEM_stage_inst_dmem_ram_1349), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n3138) );
NAND2_X1 MEM_stage_inst_dmem_U3299 ( .A1(MEM_stage_inst_dmem_ram_1829), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n3139) );
NOR2_X1 MEM_stage_inst_dmem_U3298 ( .A1(MEM_stage_inst_dmem_n3136), .A2(MEM_stage_inst_dmem_n3135), .ZN(MEM_stage_inst_dmem_n3147) );
NAND2_X1 MEM_stage_inst_dmem_U3297 ( .A1(MEM_stage_inst_dmem_n3134), .A2(MEM_stage_inst_dmem_n3133), .ZN(MEM_stage_inst_dmem_n3135) );
NAND2_X1 MEM_stage_inst_dmem_U3296 ( .A1(MEM_stage_inst_dmem_ram_2005), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n3133) );
NAND2_X1 MEM_stage_inst_dmem_U3295 ( .A1(MEM_stage_inst_dmem_ram_1285), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n3134) );
NAND2_X1 MEM_stage_inst_dmem_U3294 ( .A1(MEM_stage_inst_dmem_n3132), .A2(MEM_stage_inst_dmem_n3131), .ZN(MEM_stage_inst_dmem_n3136) );
NAND2_X1 MEM_stage_inst_dmem_U3293 ( .A1(MEM_stage_inst_dmem_ram_1157), .A2(MEM_stage_inst_dmem_n61), .ZN(MEM_stage_inst_dmem_n3131) );
NAND2_X1 MEM_stage_inst_dmem_U3292 ( .A1(MEM_stage_inst_dmem_ram_1029), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n3132) );
NAND2_X1 MEM_stage_inst_dmem_U3291 ( .A1(MEM_stage_inst_dmem_n3129), .A2(MEM_stage_inst_dmem_n3128), .ZN(MEM_stage_inst_dmem_n3149) );
NOR2_X1 MEM_stage_inst_dmem_U3290 ( .A1(MEM_stage_inst_dmem_n3127), .A2(MEM_stage_inst_dmem_n3126), .ZN(MEM_stage_inst_dmem_n3128) );
NAND2_X1 MEM_stage_inst_dmem_U3289 ( .A1(MEM_stage_inst_dmem_n3125), .A2(MEM_stage_inst_dmem_n3124), .ZN(MEM_stage_inst_dmem_n3126) );
NAND2_X1 MEM_stage_inst_dmem_U3288 ( .A1(MEM_stage_inst_dmem_ram_1669), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n3124) );
NAND2_X1 MEM_stage_inst_dmem_U3287 ( .A1(MEM_stage_inst_dmem_ram_1925), .A2(MEM_stage_inst_dmem_n72), .ZN(MEM_stage_inst_dmem_n3125) );
NAND2_X1 MEM_stage_inst_dmem_U3286 ( .A1(MEM_stage_inst_dmem_n3122), .A2(MEM_stage_inst_dmem_n3121), .ZN(MEM_stage_inst_dmem_n3127) );
NAND2_X1 MEM_stage_inst_dmem_U3285 ( .A1(MEM_stage_inst_dmem_ram_1861), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n3121) );
NAND2_X1 MEM_stage_inst_dmem_U3284 ( .A1(MEM_stage_inst_dmem_ram_1637), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n3122) );
NOR2_X1 MEM_stage_inst_dmem_U3283 ( .A1(MEM_stage_inst_dmem_n3119), .A2(MEM_stage_inst_dmem_n3118), .ZN(MEM_stage_inst_dmem_n3129) );
NAND2_X1 MEM_stage_inst_dmem_U3282 ( .A1(MEM_stage_inst_dmem_n3117), .A2(MEM_stage_inst_dmem_n3116), .ZN(MEM_stage_inst_dmem_n3118) );
NAND2_X1 MEM_stage_inst_dmem_U3281 ( .A1(MEM_stage_inst_dmem_ram_1845), .A2(MEM_stage_inst_dmem_n46), .ZN(MEM_stage_inst_dmem_n3116) );
NAND2_X1 MEM_stage_inst_dmem_U3280 ( .A1(MEM_stage_inst_dmem_ram_1653), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n3117) );
NAND2_X1 MEM_stage_inst_dmem_U3279 ( .A1(MEM_stage_inst_dmem_n3115), .A2(MEM_stage_inst_dmem_n3114), .ZN(MEM_stage_inst_dmem_n3119) );
NAND2_X1 MEM_stage_inst_dmem_U3278 ( .A1(MEM_stage_inst_dmem_ram_2021), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n3114) );
NAND2_X1 MEM_stage_inst_dmem_U3277 ( .A1(MEM_stage_inst_dmem_ram_1749), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n3115) );
NOR2_X1 MEM_stage_inst_dmem_U3276 ( .A1(MEM_stage_inst_dmem_n3111), .A2(MEM_stage_inst_dmem_n3110), .ZN(MEM_stage_inst_dmem_n3151) );
NAND2_X1 MEM_stage_inst_dmem_U3275 ( .A1(MEM_stage_inst_dmem_n3109), .A2(MEM_stage_inst_dmem_n3108), .ZN(MEM_stage_inst_dmem_n3110) );
NOR2_X1 MEM_stage_inst_dmem_U3274 ( .A1(MEM_stage_inst_dmem_n3107), .A2(MEM_stage_inst_dmem_n3106), .ZN(MEM_stage_inst_dmem_n3108) );
NAND2_X1 MEM_stage_inst_dmem_U3273 ( .A1(MEM_stage_inst_dmem_n3105), .A2(MEM_stage_inst_dmem_n3104), .ZN(MEM_stage_inst_dmem_n3106) );
NAND2_X1 MEM_stage_inst_dmem_U3272 ( .A1(MEM_stage_inst_dmem_ram_1077), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n3104) );
NAND2_X1 MEM_stage_inst_dmem_U3271 ( .A1(MEM_stage_inst_dmem_ram_1093), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n3105) );
NAND2_X1 MEM_stage_inst_dmem_U3270 ( .A1(MEM_stage_inst_dmem_n3101), .A2(MEM_stage_inst_dmem_n3100), .ZN(MEM_stage_inst_dmem_n3107) );
NAND2_X1 MEM_stage_inst_dmem_U3269 ( .A1(MEM_stage_inst_dmem_ram_1909), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n3100) );
NAND2_X1 MEM_stage_inst_dmem_U3268 ( .A1(MEM_stage_inst_dmem_ram_1893), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n3101) );
NOR2_X1 MEM_stage_inst_dmem_U3267 ( .A1(MEM_stage_inst_dmem_n3098), .A2(MEM_stage_inst_dmem_n3097), .ZN(MEM_stage_inst_dmem_n3109) );
NAND2_X1 MEM_stage_inst_dmem_U3266 ( .A1(MEM_stage_inst_dmem_n3096), .A2(MEM_stage_inst_dmem_n3095), .ZN(MEM_stage_inst_dmem_n3097) );
NAND2_X1 MEM_stage_inst_dmem_U3265 ( .A1(MEM_stage_inst_dmem_ram_1445), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n3095) );
NAND2_X1 MEM_stage_inst_dmem_U3264 ( .A1(MEM_stage_inst_dmem_ram_1765), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n3096) );
NAND2_X1 MEM_stage_inst_dmem_U3263 ( .A1(MEM_stage_inst_dmem_n3094), .A2(MEM_stage_inst_dmem_n3093), .ZN(MEM_stage_inst_dmem_n3098) );
NAND2_X1 MEM_stage_inst_dmem_U3262 ( .A1(MEM_stage_inst_dmem_ram_1061), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n3093) );
NAND2_X1 MEM_stage_inst_dmem_U3261 ( .A1(MEM_stage_inst_dmem_ram_1301), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n3094) );
NAND2_X1 MEM_stage_inst_dmem_U3260 ( .A1(MEM_stage_inst_dmem_n3091), .A2(MEM_stage_inst_dmem_n3090), .ZN(MEM_stage_inst_dmem_n3111) );
NOR2_X1 MEM_stage_inst_dmem_U3259 ( .A1(MEM_stage_inst_dmem_n3089), .A2(MEM_stage_inst_dmem_n3088), .ZN(MEM_stage_inst_dmem_n3090) );
NAND2_X1 MEM_stage_inst_dmem_U3258 ( .A1(MEM_stage_inst_dmem_n3087), .A2(MEM_stage_inst_dmem_n3086), .ZN(MEM_stage_inst_dmem_n3088) );
NAND2_X1 MEM_stage_inst_dmem_U3257 ( .A1(MEM_stage_inst_dmem_ram_1461), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n3086) );
NAND2_X1 MEM_stage_inst_dmem_U3256 ( .A1(MEM_stage_inst_dmem_ram_1589), .A2(MEM_stage_inst_dmem_n41), .ZN(MEM_stage_inst_dmem_n3087) );
NAND2_X1 MEM_stage_inst_dmem_U3255 ( .A1(MEM_stage_inst_dmem_n3084), .A2(MEM_stage_inst_dmem_n3083), .ZN(MEM_stage_inst_dmem_n3089) );
NAND2_X1 MEM_stage_inst_dmem_U3254 ( .A1(MEM_stage_inst_dmem_ram_1221), .A2(MEM_stage_inst_dmem_n36), .ZN(MEM_stage_inst_dmem_n3083) );
NAND2_X1 MEM_stage_inst_dmem_U3253 ( .A1(MEM_stage_inst_dmem_ram_1189), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n3084) );
NOR2_X1 MEM_stage_inst_dmem_U3252 ( .A1(MEM_stage_inst_dmem_n3080), .A2(MEM_stage_inst_dmem_n3079), .ZN(MEM_stage_inst_dmem_n3091) );
NAND2_X1 MEM_stage_inst_dmem_U3251 ( .A1(MEM_stage_inst_dmem_n3078), .A2(MEM_stage_inst_dmem_n3077), .ZN(MEM_stage_inst_dmem_n3079) );
NAND2_X1 MEM_stage_inst_dmem_U3250 ( .A1(MEM_stage_inst_dmem_ram_1205), .A2(MEM_stage_inst_dmem_n55), .ZN(MEM_stage_inst_dmem_n3077) );
NAND2_X1 MEM_stage_inst_dmem_U3249 ( .A1(MEM_stage_inst_dmem_ram_1685), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n3078) );
NAND2_X1 MEM_stage_inst_dmem_U3248 ( .A1(MEM_stage_inst_dmem_n3075), .A2(MEM_stage_inst_dmem_n3074), .ZN(MEM_stage_inst_dmem_n3080) );
NAND2_X1 MEM_stage_inst_dmem_U3247 ( .A1(MEM_stage_inst_dmem_ram_1333), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n3074) );
NAND2_X1 MEM_stage_inst_dmem_U3246 ( .A1(MEM_stage_inst_dmem_ram_1941), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n3075) );
NOR2_X1 MEM_stage_inst_dmem_U3245 ( .A1(MEM_stage_inst_dmem_n3072), .A2(MEM_stage_inst_dmem_n3071), .ZN(MEM_stage_inst_dmem_n3364) );
NOR2_X1 MEM_stage_inst_dmem_U3244 ( .A1(MEM_stage_inst_dmem_n3070), .A2(MEM_stage_inst_dmem_n8417), .ZN(MEM_stage_inst_dmem_n3071) );
NOR2_X1 MEM_stage_inst_dmem_U3243 ( .A1(MEM_stage_inst_dmem_n3069), .A2(MEM_stage_inst_dmem_n3068), .ZN(MEM_stage_inst_dmem_n3070) );
NAND2_X1 MEM_stage_inst_dmem_U3242 ( .A1(MEM_stage_inst_dmem_n3067), .A2(MEM_stage_inst_dmem_n3066), .ZN(MEM_stage_inst_dmem_n3068) );
NOR2_X1 MEM_stage_inst_dmem_U3241 ( .A1(MEM_stage_inst_dmem_n3065), .A2(MEM_stage_inst_dmem_n3064), .ZN(MEM_stage_inst_dmem_n3066) );
NAND2_X1 MEM_stage_inst_dmem_U3240 ( .A1(MEM_stage_inst_dmem_n3063), .A2(MEM_stage_inst_dmem_n3062), .ZN(MEM_stage_inst_dmem_n3064) );
NOR2_X1 MEM_stage_inst_dmem_U3239 ( .A1(MEM_stage_inst_dmem_n3061), .A2(MEM_stage_inst_dmem_n3060), .ZN(MEM_stage_inst_dmem_n3062) );
NAND2_X1 MEM_stage_inst_dmem_U3238 ( .A1(MEM_stage_inst_dmem_n3059), .A2(MEM_stage_inst_dmem_n3058), .ZN(MEM_stage_inst_dmem_n3060) );
NAND2_X1 MEM_stage_inst_dmem_U3237 ( .A1(MEM_stage_inst_dmem_ram_3941), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n3058) );
NAND2_X1 MEM_stage_inst_dmem_U3236 ( .A1(MEM_stage_inst_dmem_ram_3381), .A2(MEM_stage_inst_dmem_n4731), .ZN(MEM_stage_inst_dmem_n3059) );
NAND2_X1 MEM_stage_inst_dmem_U3235 ( .A1(MEM_stage_inst_dmem_n3057), .A2(MEM_stage_inst_dmem_n3056), .ZN(MEM_stage_inst_dmem_n3061) );
NAND2_X1 MEM_stage_inst_dmem_U3234 ( .A1(MEM_stage_inst_dmem_ram_3685), .A2(MEM_stage_inst_dmem_n4701), .ZN(MEM_stage_inst_dmem_n3056) );
NAND2_X1 MEM_stage_inst_dmem_U3233 ( .A1(MEM_stage_inst_dmem_ram_3813), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n3057) );
NOR2_X1 MEM_stage_inst_dmem_U3232 ( .A1(MEM_stage_inst_dmem_n3055), .A2(MEM_stage_inst_dmem_n3054), .ZN(MEM_stage_inst_dmem_n3063) );
NAND2_X1 MEM_stage_inst_dmem_U3231 ( .A1(MEM_stage_inst_dmem_n3053), .A2(MEM_stage_inst_dmem_n3052), .ZN(MEM_stage_inst_dmem_n3054) );
NAND2_X1 MEM_stage_inst_dmem_U3230 ( .A1(MEM_stage_inst_dmem_ram_4037), .A2(MEM_stage_inst_dmem_n4728), .ZN(MEM_stage_inst_dmem_n3052) );
NAND2_X1 MEM_stage_inst_dmem_U3229 ( .A1(MEM_stage_inst_dmem_ram_4053), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n3053) );
NAND2_X1 MEM_stage_inst_dmem_U3228 ( .A1(MEM_stage_inst_dmem_n3051), .A2(MEM_stage_inst_dmem_n3050), .ZN(MEM_stage_inst_dmem_n3055) );
NAND2_X1 MEM_stage_inst_dmem_U3227 ( .A1(MEM_stage_inst_dmem_ram_3237), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n3050) );
NAND2_X1 MEM_stage_inst_dmem_U3226 ( .A1(MEM_stage_inst_dmem_ram_3589), .A2(MEM_stage_inst_dmem_n8225), .ZN(MEM_stage_inst_dmem_n3051) );
BUF_X1 MEM_stage_inst_dmem_U3225 ( .A(MEM_stage_inst_dmem_n3182), .Z(MEM_stage_inst_dmem_n8225) );
NAND2_X1 MEM_stage_inst_dmem_U3224 ( .A1(MEM_stage_inst_dmem_n3049), .A2(MEM_stage_inst_dmem_n3048), .ZN(MEM_stage_inst_dmem_n3065) );
NOR2_X1 MEM_stage_inst_dmem_U3223 ( .A1(MEM_stage_inst_dmem_n3047), .A2(MEM_stage_inst_dmem_n3046), .ZN(MEM_stage_inst_dmem_n3048) );
NAND2_X1 MEM_stage_inst_dmem_U3222 ( .A1(MEM_stage_inst_dmem_n3045), .A2(MEM_stage_inst_dmem_n3044), .ZN(MEM_stage_inst_dmem_n3046) );
NAND2_X1 MEM_stage_inst_dmem_U3221 ( .A1(MEM_stage_inst_dmem_ram_3829), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n3044) );
NAND2_X1 MEM_stage_inst_dmem_U3220 ( .A1(MEM_stage_inst_dmem_ram_3205), .A2(MEM_stage_inst_dmem_n8174), .ZN(MEM_stage_inst_dmem_n3045) );
BUF_X1 MEM_stage_inst_dmem_U3219 ( .A(MEM_stage_inst_dmem_n3130), .Z(MEM_stage_inst_dmem_n8174) );
NAND2_X1 MEM_stage_inst_dmem_U3218 ( .A1(MEM_stage_inst_dmem_n3043), .A2(MEM_stage_inst_dmem_n3042), .ZN(MEM_stage_inst_dmem_n3047) );
NAND2_X1 MEM_stage_inst_dmem_U3217 ( .A1(MEM_stage_inst_dmem_ram_3349), .A2(MEM_stage_inst_dmem_n4672), .ZN(MEM_stage_inst_dmem_n3042) );
NAND2_X1 MEM_stage_inst_dmem_U3216 ( .A1(MEM_stage_inst_dmem_ram_3765), .A2(MEM_stage_inst_dmem_n4709), .ZN(MEM_stage_inst_dmem_n3043) );
NOR2_X1 MEM_stage_inst_dmem_U3215 ( .A1(MEM_stage_inst_dmem_n3041), .A2(MEM_stage_inst_dmem_n3040), .ZN(MEM_stage_inst_dmem_n3049) );
NAND2_X1 MEM_stage_inst_dmem_U3214 ( .A1(MEM_stage_inst_dmem_n3039), .A2(MEM_stage_inst_dmem_n3038), .ZN(MEM_stage_inst_dmem_n3040) );
NAND2_X1 MEM_stage_inst_dmem_U3213 ( .A1(MEM_stage_inst_dmem_ram_4069), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n3038) );
NAND2_X1 MEM_stage_inst_dmem_U3212 ( .A1(MEM_stage_inst_dmem_ram_3461), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n3039) );
NAND2_X1 MEM_stage_inst_dmem_U3211 ( .A1(MEM_stage_inst_dmem_n3037), .A2(MEM_stage_inst_dmem_n3036), .ZN(MEM_stage_inst_dmem_n3041) );
NAND2_X1 MEM_stage_inst_dmem_U3210 ( .A1(MEM_stage_inst_dmem_ram_3717), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n3036) );
NAND2_X1 MEM_stage_inst_dmem_U3209 ( .A1(MEM_stage_inst_dmem_ram_3109), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n3037) );
NOR2_X1 MEM_stage_inst_dmem_U3208 ( .A1(MEM_stage_inst_dmem_n3035), .A2(MEM_stage_inst_dmem_n3034), .ZN(MEM_stage_inst_dmem_n3067) );
NAND2_X1 MEM_stage_inst_dmem_U3207 ( .A1(MEM_stage_inst_dmem_n3033), .A2(MEM_stage_inst_dmem_n3032), .ZN(MEM_stage_inst_dmem_n3034) );
NOR2_X1 MEM_stage_inst_dmem_U3206 ( .A1(MEM_stage_inst_dmem_n3031), .A2(MEM_stage_inst_dmem_n3030), .ZN(MEM_stage_inst_dmem_n3032) );
NAND2_X1 MEM_stage_inst_dmem_U3205 ( .A1(MEM_stage_inst_dmem_n3029), .A2(MEM_stage_inst_dmem_n3028), .ZN(MEM_stage_inst_dmem_n3030) );
NAND2_X1 MEM_stage_inst_dmem_U3204 ( .A1(MEM_stage_inst_dmem_ram_3557), .A2(MEM_stage_inst_dmem_n4667), .ZN(MEM_stage_inst_dmem_n3028) );
NAND2_X1 MEM_stage_inst_dmem_U3203 ( .A1(MEM_stage_inst_dmem_ram_3749), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n3029) );
NAND2_X1 MEM_stage_inst_dmem_U3202 ( .A1(MEM_stage_inst_dmem_n3027), .A2(MEM_stage_inst_dmem_n3026), .ZN(MEM_stage_inst_dmem_n3031) );
NAND2_X1 MEM_stage_inst_dmem_U3201 ( .A1(MEM_stage_inst_dmem_ram_3317), .A2(MEM_stage_inst_dmem_n4649), .ZN(MEM_stage_inst_dmem_n3026) );
NAND2_X1 MEM_stage_inst_dmem_U3200 ( .A1(MEM_stage_inst_dmem_ram_3861), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n3027) );
NOR2_X1 MEM_stage_inst_dmem_U3199 ( .A1(MEM_stage_inst_dmem_n3025), .A2(MEM_stage_inst_dmem_n3024), .ZN(MEM_stage_inst_dmem_n3033) );
NAND2_X1 MEM_stage_inst_dmem_U3198 ( .A1(MEM_stage_inst_dmem_n3023), .A2(MEM_stage_inst_dmem_n3022), .ZN(MEM_stage_inst_dmem_n3024) );
NAND2_X1 MEM_stage_inst_dmem_U3197 ( .A1(MEM_stage_inst_dmem_ram_3189), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n3022) );
NAND2_X1 MEM_stage_inst_dmem_U3196 ( .A1(MEM_stage_inst_dmem_ram_4085), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n3023) );
NAND2_X1 MEM_stage_inst_dmem_U3195 ( .A1(MEM_stage_inst_dmem_n3021), .A2(MEM_stage_inst_dmem_n3020), .ZN(MEM_stage_inst_dmem_n3025) );
NAND2_X1 MEM_stage_inst_dmem_U3194 ( .A1(MEM_stage_inst_dmem_ram_3845), .A2(MEM_stage_inst_dmem_n37), .ZN(MEM_stage_inst_dmem_n3020) );
NAND2_X1 MEM_stage_inst_dmem_U3193 ( .A1(MEM_stage_inst_dmem_ram_3541), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n3021) );
NAND2_X1 MEM_stage_inst_dmem_U3192 ( .A1(MEM_stage_inst_dmem_n3019), .A2(MEM_stage_inst_dmem_n3018), .ZN(MEM_stage_inst_dmem_n3035) );
NOR2_X1 MEM_stage_inst_dmem_U3191 ( .A1(MEM_stage_inst_dmem_n3017), .A2(MEM_stage_inst_dmem_n3016), .ZN(MEM_stage_inst_dmem_n3018) );
NAND2_X1 MEM_stage_inst_dmem_U3190 ( .A1(MEM_stage_inst_dmem_n3015), .A2(MEM_stage_inst_dmem_n3014), .ZN(MEM_stage_inst_dmem_n3016) );
NAND2_X1 MEM_stage_inst_dmem_U3189 ( .A1(MEM_stage_inst_dmem_ram_3301), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n3014) );
NAND2_X1 MEM_stage_inst_dmem_U3188 ( .A1(MEM_stage_inst_dmem_ram_3781), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n3015) );
NAND2_X1 MEM_stage_inst_dmem_U3187 ( .A1(MEM_stage_inst_dmem_n3013), .A2(MEM_stage_inst_dmem_n3012), .ZN(MEM_stage_inst_dmem_n3017) );
NAND2_X1 MEM_stage_inst_dmem_U3186 ( .A1(MEM_stage_inst_dmem_ram_3509), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n3012) );
NAND2_X1 MEM_stage_inst_dmem_U3185 ( .A1(MEM_stage_inst_dmem_ram_3653), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n3013) );
NOR2_X1 MEM_stage_inst_dmem_U3184 ( .A1(MEM_stage_inst_dmem_n3011), .A2(MEM_stage_inst_dmem_n3010), .ZN(MEM_stage_inst_dmem_n3019) );
NAND2_X1 MEM_stage_inst_dmem_U3183 ( .A1(MEM_stage_inst_dmem_n3009), .A2(MEM_stage_inst_dmem_n3008), .ZN(MEM_stage_inst_dmem_n3010) );
NAND2_X1 MEM_stage_inst_dmem_U3182 ( .A1(MEM_stage_inst_dmem_ram_3701), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n3008) );
NAND2_X1 MEM_stage_inst_dmem_U3181 ( .A1(MEM_stage_inst_dmem_ram_3333), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n3009) );
NAND2_X1 MEM_stage_inst_dmem_U3180 ( .A1(MEM_stage_inst_dmem_n3007), .A2(MEM_stage_inst_dmem_n3006), .ZN(MEM_stage_inst_dmem_n3011) );
NAND2_X1 MEM_stage_inst_dmem_U3179 ( .A1(MEM_stage_inst_dmem_ram_3877), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n3006) );
NAND2_X1 MEM_stage_inst_dmem_U3178 ( .A1(MEM_stage_inst_dmem_ram_3733), .A2(MEM_stage_inst_dmem_n3076), .ZN(MEM_stage_inst_dmem_n3007) );
NAND2_X1 MEM_stage_inst_dmem_U3177 ( .A1(MEM_stage_inst_dmem_n3005), .A2(MEM_stage_inst_dmem_n3004), .ZN(MEM_stage_inst_dmem_n3069) );
NOR2_X1 MEM_stage_inst_dmem_U3176 ( .A1(MEM_stage_inst_dmem_n3003), .A2(MEM_stage_inst_dmem_n3002), .ZN(MEM_stage_inst_dmem_n3004) );
NAND2_X1 MEM_stage_inst_dmem_U3175 ( .A1(MEM_stage_inst_dmem_n3001), .A2(MEM_stage_inst_dmem_n3000), .ZN(MEM_stage_inst_dmem_n3002) );
NOR2_X1 MEM_stage_inst_dmem_U3174 ( .A1(MEM_stage_inst_dmem_n2999), .A2(MEM_stage_inst_dmem_n2998), .ZN(MEM_stage_inst_dmem_n3000) );
NAND2_X1 MEM_stage_inst_dmem_U3173 ( .A1(MEM_stage_inst_dmem_n2997), .A2(MEM_stage_inst_dmem_n2996), .ZN(MEM_stage_inst_dmem_n2998) );
NAND2_X1 MEM_stage_inst_dmem_U3172 ( .A1(MEM_stage_inst_dmem_ram_3269), .A2(MEM_stage_inst_dmem_n8256), .ZN(MEM_stage_inst_dmem_n2996) );
BUF_X1 MEM_stage_inst_dmem_U3171 ( .A(MEM_stage_inst_dmem_n3082), .Z(MEM_stage_inst_dmem_n8256) );
NAND2_X1 MEM_stage_inst_dmem_U3170 ( .A1(MEM_stage_inst_dmem_ram_3173), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n2997) );
NAND2_X1 MEM_stage_inst_dmem_U3169 ( .A1(MEM_stage_inst_dmem_n2995), .A2(MEM_stage_inst_dmem_n2994), .ZN(MEM_stage_inst_dmem_n2999) );
NAND2_X1 MEM_stage_inst_dmem_U3168 ( .A1(MEM_stage_inst_dmem_ram_4021), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n2994) );
NAND2_X1 MEM_stage_inst_dmem_U3167 ( .A1(MEM_stage_inst_dmem_ram_3365), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n2995) );
NOR2_X1 MEM_stage_inst_dmem_U3166 ( .A1(MEM_stage_inst_dmem_n2993), .A2(MEM_stage_inst_dmem_n2992), .ZN(MEM_stage_inst_dmem_n3001) );
NAND2_X1 MEM_stage_inst_dmem_U3165 ( .A1(MEM_stage_inst_dmem_n2991), .A2(MEM_stage_inst_dmem_n2990), .ZN(MEM_stage_inst_dmem_n2992) );
NAND2_X1 MEM_stage_inst_dmem_U3164 ( .A1(MEM_stage_inst_dmem_ram_3477), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n2990) );
NAND2_X1 MEM_stage_inst_dmem_U3163 ( .A1(MEM_stage_inst_dmem_ram_3893), .A2(MEM_stage_inst_dmem_n4740), .ZN(MEM_stage_inst_dmem_n2991) );
NAND2_X1 MEM_stage_inst_dmem_U3162 ( .A1(MEM_stage_inst_dmem_n2989), .A2(MEM_stage_inst_dmem_n2988), .ZN(MEM_stage_inst_dmem_n2993) );
NAND2_X1 MEM_stage_inst_dmem_U3161 ( .A1(MEM_stage_inst_dmem_ram_3957), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n2988) );
NAND2_X1 MEM_stage_inst_dmem_U3160 ( .A1(MEM_stage_inst_dmem_ram_3413), .A2(MEM_stage_inst_dmem_n3216), .ZN(MEM_stage_inst_dmem_n2989) );
NAND2_X1 MEM_stage_inst_dmem_U3159 ( .A1(MEM_stage_inst_dmem_n2987), .A2(MEM_stage_inst_dmem_n2986), .ZN(MEM_stage_inst_dmem_n3003) );
NOR2_X1 MEM_stage_inst_dmem_U3158 ( .A1(MEM_stage_inst_dmem_n2985), .A2(MEM_stage_inst_dmem_n2984), .ZN(MEM_stage_inst_dmem_n2986) );
NAND2_X1 MEM_stage_inst_dmem_U3157 ( .A1(MEM_stage_inst_dmem_n2983), .A2(MEM_stage_inst_dmem_n2982), .ZN(MEM_stage_inst_dmem_n2984) );
NAND2_X1 MEM_stage_inst_dmem_U3156 ( .A1(MEM_stage_inst_dmem_ram_3493), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n2982) );
NAND2_X1 MEM_stage_inst_dmem_U3155 ( .A1(MEM_stage_inst_dmem_ram_3157), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n2983) );
NAND2_X1 MEM_stage_inst_dmem_U3154 ( .A1(MEM_stage_inst_dmem_n2981), .A2(MEM_stage_inst_dmem_n2980), .ZN(MEM_stage_inst_dmem_n2985) );
NAND2_X1 MEM_stage_inst_dmem_U3153 ( .A1(MEM_stage_inst_dmem_ram_3989), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n2980) );
NAND2_X1 MEM_stage_inst_dmem_U3152 ( .A1(MEM_stage_inst_dmem_ram_3973), .A2(MEM_stage_inst_dmem_n8193), .ZN(MEM_stage_inst_dmem_n2981) );
BUF_X1 MEM_stage_inst_dmem_U3151 ( .A(MEM_stage_inst_dmem_n3123), .Z(MEM_stage_inst_dmem_n8193) );
NOR2_X1 MEM_stage_inst_dmem_U3150 ( .A1(MEM_stage_inst_dmem_n2979), .A2(MEM_stage_inst_dmem_n2978), .ZN(MEM_stage_inst_dmem_n2987) );
NAND2_X1 MEM_stage_inst_dmem_U3149 ( .A1(MEM_stage_inst_dmem_n2977), .A2(MEM_stage_inst_dmem_n2976), .ZN(MEM_stage_inst_dmem_n2978) );
NAND2_X1 MEM_stage_inst_dmem_U3148 ( .A1(MEM_stage_inst_dmem_ram_3397), .A2(MEM_stage_inst_dmem_n4706), .ZN(MEM_stage_inst_dmem_n2976) );
NAND2_X1 MEM_stage_inst_dmem_U3147 ( .A1(MEM_stage_inst_dmem_ram_3221), .A2(MEM_stage_inst_dmem_n44), .ZN(MEM_stage_inst_dmem_n2977) );
NAND2_X1 MEM_stage_inst_dmem_U3146 ( .A1(MEM_stage_inst_dmem_n2975), .A2(MEM_stage_inst_dmem_n2974), .ZN(MEM_stage_inst_dmem_n2979) );
NAND2_X1 MEM_stage_inst_dmem_U3145 ( .A1(MEM_stage_inst_dmem_ram_3909), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n2974) );
NAND2_X1 MEM_stage_inst_dmem_U3144 ( .A1(MEM_stage_inst_dmem_ram_3093), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n2975) );
NOR2_X1 MEM_stage_inst_dmem_U3143 ( .A1(MEM_stage_inst_dmem_n2973), .A2(MEM_stage_inst_dmem_n2972), .ZN(MEM_stage_inst_dmem_n3005) );
NAND2_X1 MEM_stage_inst_dmem_U3142 ( .A1(MEM_stage_inst_dmem_n2971), .A2(MEM_stage_inst_dmem_n2970), .ZN(MEM_stage_inst_dmem_n2972) );
NOR2_X1 MEM_stage_inst_dmem_U3141 ( .A1(MEM_stage_inst_dmem_n2969), .A2(MEM_stage_inst_dmem_n2968), .ZN(MEM_stage_inst_dmem_n2970) );
NAND2_X1 MEM_stage_inst_dmem_U3140 ( .A1(MEM_stage_inst_dmem_n2967), .A2(MEM_stage_inst_dmem_n2966), .ZN(MEM_stage_inst_dmem_n2968) );
NAND2_X1 MEM_stage_inst_dmem_U3139 ( .A1(MEM_stage_inst_dmem_ram_3621), .A2(MEM_stage_inst_dmem_n4692), .ZN(MEM_stage_inst_dmem_n2966) );
NAND2_X1 MEM_stage_inst_dmem_U3138 ( .A1(MEM_stage_inst_dmem_ram_3445), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n2967) );
NAND2_X1 MEM_stage_inst_dmem_U3137 ( .A1(MEM_stage_inst_dmem_n2965), .A2(MEM_stage_inst_dmem_n2964), .ZN(MEM_stage_inst_dmem_n2969) );
NAND2_X1 MEM_stage_inst_dmem_U3136 ( .A1(MEM_stage_inst_dmem_ram_3525), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n2964) );
NAND2_X1 MEM_stage_inst_dmem_U3135 ( .A1(MEM_stage_inst_dmem_ram_3797), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n2965) );
NOR2_X1 MEM_stage_inst_dmem_U3134 ( .A1(MEM_stage_inst_dmem_n2963), .A2(MEM_stage_inst_dmem_n2962), .ZN(MEM_stage_inst_dmem_n2971) );
NAND2_X1 MEM_stage_inst_dmem_U3133 ( .A1(MEM_stage_inst_dmem_n2961), .A2(MEM_stage_inst_dmem_n2960), .ZN(MEM_stage_inst_dmem_n2962) );
NAND2_X1 MEM_stage_inst_dmem_U3132 ( .A1(MEM_stage_inst_dmem_ram_3925), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n2960) );
NAND2_X1 MEM_stage_inst_dmem_U3131 ( .A1(MEM_stage_inst_dmem_ram_3253), .A2(MEM_stage_inst_dmem_n55), .ZN(MEM_stage_inst_dmem_n2961) );
NAND2_X1 MEM_stage_inst_dmem_U3130 ( .A1(MEM_stage_inst_dmem_n2959), .A2(MEM_stage_inst_dmem_n2958), .ZN(MEM_stage_inst_dmem_n2963) );
NAND2_X1 MEM_stage_inst_dmem_U3129 ( .A1(MEM_stage_inst_dmem_ram_3429), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n2958) );
NAND2_X1 MEM_stage_inst_dmem_U3128 ( .A1(MEM_stage_inst_dmem_ram_3077), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n2959) );
NAND2_X1 MEM_stage_inst_dmem_U3127 ( .A1(MEM_stage_inst_dmem_n2957), .A2(MEM_stage_inst_dmem_n2956), .ZN(MEM_stage_inst_dmem_n2973) );
NOR2_X1 MEM_stage_inst_dmem_U3126 ( .A1(MEM_stage_inst_dmem_n2955), .A2(MEM_stage_inst_dmem_n2954), .ZN(MEM_stage_inst_dmem_n2956) );
NAND2_X1 MEM_stage_inst_dmem_U3125 ( .A1(MEM_stage_inst_dmem_n2953), .A2(MEM_stage_inst_dmem_n2952), .ZN(MEM_stage_inst_dmem_n2954) );
NAND2_X1 MEM_stage_inst_dmem_U3124 ( .A1(MEM_stage_inst_dmem_ram_4005), .A2(MEM_stage_inst_dmem_n4675), .ZN(MEM_stage_inst_dmem_n2952) );
NAND2_X1 MEM_stage_inst_dmem_U3123 ( .A1(MEM_stage_inst_dmem_ram_3605), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n2953) );
NAND2_X1 MEM_stage_inst_dmem_U3122 ( .A1(MEM_stage_inst_dmem_n2951), .A2(MEM_stage_inst_dmem_n2950), .ZN(MEM_stage_inst_dmem_n2955) );
NAND2_X1 MEM_stage_inst_dmem_U3121 ( .A1(MEM_stage_inst_dmem_ram_3573), .A2(MEM_stage_inst_dmem_n64), .ZN(MEM_stage_inst_dmem_n2950) );
NAND2_X1 MEM_stage_inst_dmem_U3120 ( .A1(MEM_stage_inst_dmem_ram_3669), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n2951) );
NOR2_X1 MEM_stage_inst_dmem_U3119 ( .A1(MEM_stage_inst_dmem_n2949), .A2(MEM_stage_inst_dmem_n2948), .ZN(MEM_stage_inst_dmem_n2957) );
NAND2_X1 MEM_stage_inst_dmem_U3118 ( .A1(MEM_stage_inst_dmem_n2947), .A2(MEM_stage_inst_dmem_n2946), .ZN(MEM_stage_inst_dmem_n2948) );
NAND2_X1 MEM_stage_inst_dmem_U3117 ( .A1(MEM_stage_inst_dmem_ram_3637), .A2(MEM_stage_inst_dmem_n8169), .ZN(MEM_stage_inst_dmem_n2946) );
BUF_X1 MEM_stage_inst_dmem_U3116 ( .A(MEM_stage_inst_dmem_n3085), .Z(MEM_stage_inst_dmem_n8169) );
NAND2_X1 MEM_stage_inst_dmem_U3115 ( .A1(MEM_stage_inst_dmem_ram_3125), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n2947) );
NAND2_X1 MEM_stage_inst_dmem_U3114 ( .A1(MEM_stage_inst_dmem_n2945), .A2(MEM_stage_inst_dmem_n2944), .ZN(MEM_stage_inst_dmem_n2949) );
NAND2_X1 MEM_stage_inst_dmem_U3113 ( .A1(MEM_stage_inst_dmem_ram_3141), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n2944) );
NAND2_X1 MEM_stage_inst_dmem_U3112 ( .A1(MEM_stage_inst_dmem_ram_3285), .A2(MEM_stage_inst_dmem_n8206), .ZN(MEM_stage_inst_dmem_n2945) );
BUF_X1 MEM_stage_inst_dmem_U3111 ( .A(MEM_stage_inst_dmem_n3220), .Z(MEM_stage_inst_dmem_n8206) );
NOR2_X1 MEM_stage_inst_dmem_U3110 ( .A1(MEM_stage_inst_dmem_n2943), .A2(MEM_stage_inst_dmem_n8551), .ZN(MEM_stage_inst_dmem_n3072) );
NOR2_X1 MEM_stage_inst_dmem_U3109 ( .A1(MEM_stage_inst_dmem_n2942), .A2(MEM_stage_inst_dmem_n2941), .ZN(MEM_stage_inst_dmem_n2943) );
NAND2_X1 MEM_stage_inst_dmem_U3108 ( .A1(MEM_stage_inst_dmem_n2940), .A2(MEM_stage_inst_dmem_n2939), .ZN(MEM_stage_inst_dmem_n2941) );
NOR2_X1 MEM_stage_inst_dmem_U3107 ( .A1(MEM_stage_inst_dmem_n2938), .A2(MEM_stage_inst_dmem_n2937), .ZN(MEM_stage_inst_dmem_n2939) );
NAND2_X1 MEM_stage_inst_dmem_U3106 ( .A1(MEM_stage_inst_dmem_n2936), .A2(MEM_stage_inst_dmem_n2935), .ZN(MEM_stage_inst_dmem_n2937) );
NOR2_X1 MEM_stage_inst_dmem_U3105 ( .A1(MEM_stage_inst_dmem_n2934), .A2(MEM_stage_inst_dmem_n2933), .ZN(MEM_stage_inst_dmem_n2935) );
NAND2_X1 MEM_stage_inst_dmem_U3104 ( .A1(MEM_stage_inst_dmem_n2932), .A2(MEM_stage_inst_dmem_n2931), .ZN(MEM_stage_inst_dmem_n2933) );
NAND2_X1 MEM_stage_inst_dmem_U3103 ( .A1(MEM_stage_inst_dmem_ram_245), .A2(MEM_stage_inst_dmem_n4649), .ZN(MEM_stage_inst_dmem_n2931) );
NAND2_X1 MEM_stage_inst_dmem_U3102 ( .A1(MEM_stage_inst_dmem_ram_1013), .A2(MEM_stage_inst_dmem_n3199), .ZN(MEM_stage_inst_dmem_n2932) );
NAND2_X1 MEM_stage_inst_dmem_U3101 ( .A1(MEM_stage_inst_dmem_n2930), .A2(MEM_stage_inst_dmem_n2929), .ZN(MEM_stage_inst_dmem_n2934) );
NAND2_X1 MEM_stage_inst_dmem_U3100 ( .A1(MEM_stage_inst_dmem_ram_533), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n2929) );
NAND2_X1 MEM_stage_inst_dmem_U3099 ( .A1(MEM_stage_inst_dmem_ram_597), .A2(MEM_stage_inst_dmem_n3140), .ZN(MEM_stage_inst_dmem_n2930) );
NOR2_X1 MEM_stage_inst_dmem_U3098 ( .A1(MEM_stage_inst_dmem_n2928), .A2(MEM_stage_inst_dmem_n2927), .ZN(MEM_stage_inst_dmem_n2936) );
NAND2_X1 MEM_stage_inst_dmem_U3097 ( .A1(MEM_stage_inst_dmem_n2926), .A2(MEM_stage_inst_dmem_n2925), .ZN(MEM_stage_inst_dmem_n2927) );
NAND2_X1 MEM_stage_inst_dmem_U3096 ( .A1(MEM_stage_inst_dmem_ram_997), .A2(MEM_stage_inst_dmem_n3113), .ZN(MEM_stage_inst_dmem_n2925) );
NAND2_X1 MEM_stage_inst_dmem_U3095 ( .A1(MEM_stage_inst_dmem_ram_725), .A2(MEM_stage_inst_dmem_n3112), .ZN(MEM_stage_inst_dmem_n2926) );
NAND2_X1 MEM_stage_inst_dmem_U3094 ( .A1(MEM_stage_inst_dmem_n2924), .A2(MEM_stage_inst_dmem_n2923), .ZN(MEM_stage_inst_dmem_n2928) );
NAND2_X1 MEM_stage_inst_dmem_U3093 ( .A1(MEM_stage_inst_dmem_ram_405), .A2(MEM_stage_inst_dmem_n3160), .ZN(MEM_stage_inst_dmem_n2923) );
NAND2_X1 MEM_stage_inst_dmem_U3092 ( .A1(MEM_stage_inst_dmem_ram_389), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n2924) );
NAND2_X1 MEM_stage_inst_dmem_U3091 ( .A1(MEM_stage_inst_dmem_n2922), .A2(MEM_stage_inst_dmem_n2921), .ZN(MEM_stage_inst_dmem_n2938) );
NOR2_X1 MEM_stage_inst_dmem_U3090 ( .A1(MEM_stage_inst_dmem_n2920), .A2(MEM_stage_inst_dmem_n2919), .ZN(MEM_stage_inst_dmem_n2921) );
NAND2_X1 MEM_stage_inst_dmem_U3089 ( .A1(MEM_stage_inst_dmem_n2918), .A2(MEM_stage_inst_dmem_n2917), .ZN(MEM_stage_inst_dmem_n2919) );
NAND2_X1 MEM_stage_inst_dmem_U3088 ( .A1(MEM_stage_inst_dmem_ram_485), .A2(MEM_stage_inst_dmem_n4667), .ZN(MEM_stage_inst_dmem_n2917) );
NAND2_X1 MEM_stage_inst_dmem_U3087 ( .A1(MEM_stage_inst_dmem_ram_181), .A2(MEM_stage_inst_dmem_n55), .ZN(MEM_stage_inst_dmem_n2918) );
NAND2_X1 MEM_stage_inst_dmem_U3086 ( .A1(MEM_stage_inst_dmem_n2916), .A2(MEM_stage_inst_dmem_n2915), .ZN(MEM_stage_inst_dmem_n2920) );
NAND2_X1 MEM_stage_inst_dmem_U3085 ( .A1(MEM_stage_inst_dmem_ram_549), .A2(MEM_stage_inst_dmem_n4692), .ZN(MEM_stage_inst_dmem_n2915) );
NAND2_X1 MEM_stage_inst_dmem_U3084 ( .A1(MEM_stage_inst_dmem_ram_677), .A2(MEM_stage_inst_dmem_n3155), .ZN(MEM_stage_inst_dmem_n2916) );
NOR2_X1 MEM_stage_inst_dmem_U3083 ( .A1(MEM_stage_inst_dmem_n2914), .A2(MEM_stage_inst_dmem_n2913), .ZN(MEM_stage_inst_dmem_n2922) );
NAND2_X1 MEM_stage_inst_dmem_U3082 ( .A1(MEM_stage_inst_dmem_n2912), .A2(MEM_stage_inst_dmem_n2911), .ZN(MEM_stage_inst_dmem_n2913) );
NAND2_X1 MEM_stage_inst_dmem_U3081 ( .A1(MEM_stage_inst_dmem_ram_213), .A2(MEM_stage_inst_dmem_n3220), .ZN(MEM_stage_inst_dmem_n2911) );
NAND2_X1 MEM_stage_inst_dmem_U3080 ( .A1(MEM_stage_inst_dmem_ram_373), .A2(MEM_stage_inst_dmem_n4721), .ZN(MEM_stage_inst_dmem_n2912) );
NAND2_X1 MEM_stage_inst_dmem_U3079 ( .A1(MEM_stage_inst_dmem_n2910), .A2(MEM_stage_inst_dmem_n2909), .ZN(MEM_stage_inst_dmem_n2914) );
NAND2_X1 MEM_stage_inst_dmem_U3078 ( .A1(MEM_stage_inst_dmem_ram_37), .A2(MEM_stage_inst_dmem_n3092), .ZN(MEM_stage_inst_dmem_n2909) );
NAND2_X1 MEM_stage_inst_dmem_U3077 ( .A1(MEM_stage_inst_dmem_ram_261), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n2910) );
NOR2_X1 MEM_stage_inst_dmem_U3076 ( .A1(MEM_stage_inst_dmem_n2908), .A2(MEM_stage_inst_dmem_n2907), .ZN(MEM_stage_inst_dmem_n2940) );
NAND2_X1 MEM_stage_inst_dmem_U3075 ( .A1(MEM_stage_inst_dmem_n2906), .A2(MEM_stage_inst_dmem_n2905), .ZN(MEM_stage_inst_dmem_n2907) );
NOR2_X1 MEM_stage_inst_dmem_U3074 ( .A1(MEM_stage_inst_dmem_n2904), .A2(MEM_stage_inst_dmem_n2903), .ZN(MEM_stage_inst_dmem_n2905) );
NAND2_X1 MEM_stage_inst_dmem_U3073 ( .A1(MEM_stage_inst_dmem_n2902), .A2(MEM_stage_inst_dmem_n2901), .ZN(MEM_stage_inst_dmem_n2903) );
NAND2_X1 MEM_stage_inst_dmem_U3072 ( .A1(MEM_stage_inst_dmem_ram_901), .A2(MEM_stage_inst_dmem_n3123), .ZN(MEM_stage_inst_dmem_n2901) );
NAND2_X1 MEM_stage_inst_dmem_U3071 ( .A1(MEM_stage_inst_dmem_ram_629), .A2(MEM_stage_inst_dmem_n4652), .ZN(MEM_stage_inst_dmem_n2902) );
NAND2_X1 MEM_stage_inst_dmem_U3070 ( .A1(MEM_stage_inst_dmem_n2900), .A2(MEM_stage_inst_dmem_n2899), .ZN(MEM_stage_inst_dmem_n2904) );
NAND2_X1 MEM_stage_inst_dmem_U3069 ( .A1(MEM_stage_inst_dmem_ram_357), .A2(MEM_stage_inst_dmem_n3217), .ZN(MEM_stage_inst_dmem_n2899) );
NAND2_X1 MEM_stage_inst_dmem_U3068 ( .A1(MEM_stage_inst_dmem_ram_165), .A2(MEM_stage_inst_dmem_n3081), .ZN(MEM_stage_inst_dmem_n2900) );
NOR2_X1 MEM_stage_inst_dmem_U3067 ( .A1(MEM_stage_inst_dmem_n2898), .A2(MEM_stage_inst_dmem_n2897), .ZN(MEM_stage_inst_dmem_n2906) );
NAND2_X1 MEM_stage_inst_dmem_U3066 ( .A1(MEM_stage_inst_dmem_n2896), .A2(MEM_stage_inst_dmem_n2895), .ZN(MEM_stage_inst_dmem_n2897) );
NAND2_X1 MEM_stage_inst_dmem_U3065 ( .A1(MEM_stage_inst_dmem_ram_229), .A2(MEM_stage_inst_dmem_n3152), .ZN(MEM_stage_inst_dmem_n2895) );
NAND2_X1 MEM_stage_inst_dmem_U3064 ( .A1(MEM_stage_inst_dmem_ram_277), .A2(MEM_stage_inst_dmem_n4672), .ZN(MEM_stage_inst_dmem_n2896) );
NAND2_X1 MEM_stage_inst_dmem_U3063 ( .A1(MEM_stage_inst_dmem_n2894), .A2(MEM_stage_inst_dmem_n2893), .ZN(MEM_stage_inst_dmem_n2898) );
NAND2_X1 MEM_stage_inst_dmem_U3062 ( .A1(MEM_stage_inst_dmem_ram_565), .A2(MEM_stage_inst_dmem_n3085), .ZN(MEM_stage_inst_dmem_n2893) );
NAND2_X1 MEM_stage_inst_dmem_U3061 ( .A1(MEM_stage_inst_dmem_ram_709), .A2(MEM_stage_inst_dmem_n3192), .ZN(MEM_stage_inst_dmem_n2894) );
NAND2_X1 MEM_stage_inst_dmem_U3060 ( .A1(MEM_stage_inst_dmem_n2892), .A2(MEM_stage_inst_dmem_n2891), .ZN(MEM_stage_inst_dmem_n2908) );
NOR2_X1 MEM_stage_inst_dmem_U3059 ( .A1(MEM_stage_inst_dmem_n2890), .A2(MEM_stage_inst_dmem_n2889), .ZN(MEM_stage_inst_dmem_n2891) );
NAND2_X1 MEM_stage_inst_dmem_U3058 ( .A1(MEM_stage_inst_dmem_n2888), .A2(MEM_stage_inst_dmem_n2887), .ZN(MEM_stage_inst_dmem_n2889) );
NAND2_X1 MEM_stage_inst_dmem_U3057 ( .A1(MEM_stage_inst_dmem_ram_421), .A2(MEM_stage_inst_dmem_n4772), .ZN(MEM_stage_inst_dmem_n2887) );
NAND2_X1 MEM_stage_inst_dmem_U3056 ( .A1(MEM_stage_inst_dmem_ram_149), .A2(MEM_stage_inst_dmem_n44), .ZN(MEM_stage_inst_dmem_n2888) );
NAND2_X1 MEM_stage_inst_dmem_U3055 ( .A1(MEM_stage_inst_dmem_n2886), .A2(MEM_stage_inst_dmem_n2885), .ZN(MEM_stage_inst_dmem_n2890) );
NAND2_X1 MEM_stage_inst_dmem_U3054 ( .A1(MEM_stage_inst_dmem_ram_917), .A2(MEM_stage_inst_dmem_n3073), .ZN(MEM_stage_inst_dmem_n2885) );
NAND2_X1 MEM_stage_inst_dmem_U3053 ( .A1(MEM_stage_inst_dmem_ram_21), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n2886) );
NOR2_X1 MEM_stage_inst_dmem_U3052 ( .A1(MEM_stage_inst_dmem_n2884), .A2(MEM_stage_inst_dmem_n2883), .ZN(MEM_stage_inst_dmem_n2892) );
NAND2_X1 MEM_stage_inst_dmem_U3051 ( .A1(MEM_stage_inst_dmem_n2882), .A2(MEM_stage_inst_dmem_n2881), .ZN(MEM_stage_inst_dmem_n2883) );
NAND2_X1 MEM_stage_inst_dmem_U3050 ( .A1(MEM_stage_inst_dmem_ram_837), .A2(MEM_stage_inst_dmem_n3120), .ZN(MEM_stage_inst_dmem_n2881) );
NAND2_X1 MEM_stage_inst_dmem_U3049 ( .A1(MEM_stage_inst_dmem_ram_293), .A2(MEM_stage_inst_dmem_n3209), .ZN(MEM_stage_inst_dmem_n2882) );
NAND2_X1 MEM_stage_inst_dmem_U3048 ( .A1(MEM_stage_inst_dmem_n2880), .A2(MEM_stage_inst_dmem_n2879), .ZN(MEM_stage_inst_dmem_n2884) );
NAND2_X1 MEM_stage_inst_dmem_U3047 ( .A1(MEM_stage_inst_dmem_ram_53), .A2(MEM_stage_inst_dmem_n3103), .ZN(MEM_stage_inst_dmem_n2879) );
NAND2_X1 MEM_stage_inst_dmem_U3046 ( .A1(MEM_stage_inst_dmem_ram_981), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n2880) );
NAND2_X1 MEM_stage_inst_dmem_U3045 ( .A1(MEM_stage_inst_dmem_n2878), .A2(MEM_stage_inst_dmem_n2877), .ZN(MEM_stage_inst_dmem_n2942) );
NOR2_X1 MEM_stage_inst_dmem_U3044 ( .A1(MEM_stage_inst_dmem_n2876), .A2(MEM_stage_inst_dmem_n2875), .ZN(MEM_stage_inst_dmem_n2877) );
NAND2_X1 MEM_stage_inst_dmem_U3043 ( .A1(MEM_stage_inst_dmem_n2874), .A2(MEM_stage_inst_dmem_n2873), .ZN(MEM_stage_inst_dmem_n2875) );
NOR2_X1 MEM_stage_inst_dmem_U3042 ( .A1(MEM_stage_inst_dmem_n2872), .A2(MEM_stage_inst_dmem_n2871), .ZN(MEM_stage_inst_dmem_n2873) );
NAND2_X1 MEM_stage_inst_dmem_U3041 ( .A1(MEM_stage_inst_dmem_n2870), .A2(MEM_stage_inst_dmem_n2869), .ZN(MEM_stage_inst_dmem_n2871) );
NAND2_X1 MEM_stage_inst_dmem_U3040 ( .A1(MEM_stage_inst_dmem_ram_773), .A2(MEM_stage_inst_dmem_n37), .ZN(MEM_stage_inst_dmem_n2869) );
NAND2_X1 MEM_stage_inst_dmem_U3039 ( .A1(MEM_stage_inst_dmem_ram_613), .A2(MEM_stage_inst_dmem_n4701), .ZN(MEM_stage_inst_dmem_n2870) );
NAND2_X1 MEM_stage_inst_dmem_U3038 ( .A1(MEM_stage_inst_dmem_n2868), .A2(MEM_stage_inst_dmem_n2867), .ZN(MEM_stage_inst_dmem_n2872) );
NAND2_X1 MEM_stage_inst_dmem_U3037 ( .A1(MEM_stage_inst_dmem_ram_197), .A2(MEM_stage_inst_dmem_n3082), .ZN(MEM_stage_inst_dmem_n2867) );
NAND2_X1 MEM_stage_inst_dmem_U3036 ( .A1(MEM_stage_inst_dmem_ram_661), .A2(MEM_stage_inst_dmem_n3076), .ZN(MEM_stage_inst_dmem_n2868) );
NOR2_X1 MEM_stage_inst_dmem_U3035 ( .A1(MEM_stage_inst_dmem_n2866), .A2(MEM_stage_inst_dmem_n2865), .ZN(MEM_stage_inst_dmem_n2874) );
NAND2_X1 MEM_stage_inst_dmem_U3034 ( .A1(MEM_stage_inst_dmem_n2864), .A2(MEM_stage_inst_dmem_n2863), .ZN(MEM_stage_inst_dmem_n2865) );
NAND2_X1 MEM_stage_inst_dmem_U3033 ( .A1(MEM_stage_inst_dmem_ram_69), .A2(MEM_stage_inst_dmem_n3102), .ZN(MEM_stage_inst_dmem_n2863) );
NAND2_X1 MEM_stage_inst_dmem_U3032 ( .A1(MEM_stage_inst_dmem_ram_469), .A2(MEM_stage_inst_dmem_n3174), .ZN(MEM_stage_inst_dmem_n2864) );
NAND2_X1 MEM_stage_inst_dmem_U3031 ( .A1(MEM_stage_inst_dmem_n2862), .A2(MEM_stage_inst_dmem_n2861), .ZN(MEM_stage_inst_dmem_n2866) );
NAND2_X1 MEM_stage_inst_dmem_U3030 ( .A1(MEM_stage_inst_dmem_ram_949), .A2(MEM_stage_inst_dmem_n3163), .ZN(MEM_stage_inst_dmem_n2861) );
NAND2_X1 MEM_stage_inst_dmem_U3029 ( .A1(MEM_stage_inst_dmem_ram_821), .A2(MEM_stage_inst_dmem_n4740), .ZN(MEM_stage_inst_dmem_n2862) );
NAND2_X1 MEM_stage_inst_dmem_U3028 ( .A1(MEM_stage_inst_dmem_n2860), .A2(MEM_stage_inst_dmem_n2859), .ZN(MEM_stage_inst_dmem_n2876) );
NOR2_X1 MEM_stage_inst_dmem_U3027 ( .A1(MEM_stage_inst_dmem_n2858), .A2(MEM_stage_inst_dmem_n2857), .ZN(MEM_stage_inst_dmem_n2859) );
NAND2_X1 MEM_stage_inst_dmem_U3026 ( .A1(MEM_stage_inst_dmem_n2856), .A2(MEM_stage_inst_dmem_n2855), .ZN(MEM_stage_inst_dmem_n2857) );
NAND2_X1 MEM_stage_inst_dmem_U3025 ( .A1(MEM_stage_inst_dmem_ram_309), .A2(MEM_stage_inst_dmem_n4731), .ZN(MEM_stage_inst_dmem_n2855) );
NAND2_X1 MEM_stage_inst_dmem_U3024 ( .A1(MEM_stage_inst_dmem_ram_85), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n2856) );
NAND2_X1 MEM_stage_inst_dmem_U3023 ( .A1(MEM_stage_inst_dmem_n2854), .A2(MEM_stage_inst_dmem_n2853), .ZN(MEM_stage_inst_dmem_n2858) );
NAND2_X1 MEM_stage_inst_dmem_U3022 ( .A1(MEM_stage_inst_dmem_ram_805), .A2(MEM_stage_inst_dmem_n3137), .ZN(MEM_stage_inst_dmem_n2853) );
NAND2_X1 MEM_stage_inst_dmem_U3021 ( .A1(MEM_stage_inst_dmem_ram_101), .A2(MEM_stage_inst_dmem_n3179), .ZN(MEM_stage_inst_dmem_n2854) );
NOR2_X1 MEM_stage_inst_dmem_U3020 ( .A1(MEM_stage_inst_dmem_n2852), .A2(MEM_stage_inst_dmem_n2851), .ZN(MEM_stage_inst_dmem_n2860) );
NAND2_X1 MEM_stage_inst_dmem_U3019 ( .A1(MEM_stage_inst_dmem_n2850), .A2(MEM_stage_inst_dmem_n2849), .ZN(MEM_stage_inst_dmem_n2851) );
NAND2_X1 MEM_stage_inst_dmem_U3018 ( .A1(MEM_stage_inst_dmem_ram_133), .A2(MEM_stage_inst_dmem_n3130), .ZN(MEM_stage_inst_dmem_n2849) );
NAND2_X1 MEM_stage_inst_dmem_U3017 ( .A1(MEM_stage_inst_dmem_ram_741), .A2(MEM_stage_inst_dmem_n4769), .ZN(MEM_stage_inst_dmem_n2850) );
NAND2_X1 MEM_stage_inst_dmem_U3016 ( .A1(MEM_stage_inst_dmem_n2848), .A2(MEM_stage_inst_dmem_n2847), .ZN(MEM_stage_inst_dmem_n2852) );
NAND2_X1 MEM_stage_inst_dmem_U3015 ( .A1(MEM_stage_inst_dmem_ram_517), .A2(MEM_stage_inst_dmem_n3182), .ZN(MEM_stage_inst_dmem_n2847) );
NAND2_X1 MEM_stage_inst_dmem_U3014 ( .A1(MEM_stage_inst_dmem_ram_581), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n2848) );
NOR2_X1 MEM_stage_inst_dmem_U3013 ( .A1(MEM_stage_inst_dmem_n2846), .A2(MEM_stage_inst_dmem_n2845), .ZN(MEM_stage_inst_dmem_n2878) );
NAND2_X1 MEM_stage_inst_dmem_U3012 ( .A1(MEM_stage_inst_dmem_n2844), .A2(MEM_stage_inst_dmem_n2843), .ZN(MEM_stage_inst_dmem_n2845) );
NOR2_X1 MEM_stage_inst_dmem_U3011 ( .A1(MEM_stage_inst_dmem_n2842), .A2(MEM_stage_inst_dmem_n2841), .ZN(MEM_stage_inst_dmem_n2843) );
NAND2_X1 MEM_stage_inst_dmem_U3010 ( .A1(MEM_stage_inst_dmem_n2840), .A2(MEM_stage_inst_dmem_n2839), .ZN(MEM_stage_inst_dmem_n2841) );
NAND2_X1 MEM_stage_inst_dmem_U3009 ( .A1(MEM_stage_inst_dmem_ram_325), .A2(MEM_stage_inst_dmem_n4706), .ZN(MEM_stage_inst_dmem_n2839) );
NAND2_X1 MEM_stage_inst_dmem_U3008 ( .A1(MEM_stage_inst_dmem_ram_645), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n2840) );
NAND2_X1 MEM_stage_inst_dmem_U3007 ( .A1(MEM_stage_inst_dmem_n2838), .A2(MEM_stage_inst_dmem_n2837), .ZN(MEM_stage_inst_dmem_n2842) );
NAND2_X1 MEM_stage_inst_dmem_U3006 ( .A1(MEM_stage_inst_dmem_ram_117), .A2(MEM_stage_inst_dmem_n4710), .ZN(MEM_stage_inst_dmem_n2837) );
NAND2_X1 MEM_stage_inst_dmem_U3005 ( .A1(MEM_stage_inst_dmem_ram_341), .A2(MEM_stage_inst_dmem_n3216), .ZN(MEM_stage_inst_dmem_n2838) );
NOR2_X1 MEM_stage_inst_dmem_U3004 ( .A1(MEM_stage_inst_dmem_n2836), .A2(MEM_stage_inst_dmem_n2835), .ZN(MEM_stage_inst_dmem_n2844) );
NAND2_X1 MEM_stage_inst_dmem_U3003 ( .A1(MEM_stage_inst_dmem_n2834), .A2(MEM_stage_inst_dmem_n2833), .ZN(MEM_stage_inst_dmem_n2835) );
NAND2_X1 MEM_stage_inst_dmem_U3002 ( .A1(MEM_stage_inst_dmem_ram_437), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n2833) );
NAND2_X1 MEM_stage_inst_dmem_U3001 ( .A1(MEM_stage_inst_dmem_ram_453), .A2(MEM_stage_inst_dmem_n3173), .ZN(MEM_stage_inst_dmem_n2834) );
NAND2_X1 MEM_stage_inst_dmem_U3000 ( .A1(MEM_stage_inst_dmem_n2832), .A2(MEM_stage_inst_dmem_n2831), .ZN(MEM_stage_inst_dmem_n2836) );
NAND2_X1 MEM_stage_inst_dmem_U2999 ( .A1(MEM_stage_inst_dmem_ram_869), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n2831) );
NAND2_X1 MEM_stage_inst_dmem_U2998 ( .A1(MEM_stage_inst_dmem_ram_853), .A2(MEM_stage_inst_dmem_n3141), .ZN(MEM_stage_inst_dmem_n2832) );
NAND2_X1 MEM_stage_inst_dmem_U2997 ( .A1(MEM_stage_inst_dmem_n2830), .A2(MEM_stage_inst_dmem_n2829), .ZN(MEM_stage_inst_dmem_n2846) );
NOR2_X1 MEM_stage_inst_dmem_U2996 ( .A1(MEM_stage_inst_dmem_n2828), .A2(MEM_stage_inst_dmem_n2827), .ZN(MEM_stage_inst_dmem_n2829) );
NAND2_X1 MEM_stage_inst_dmem_U2995 ( .A1(MEM_stage_inst_dmem_n2826), .A2(MEM_stage_inst_dmem_n2825), .ZN(MEM_stage_inst_dmem_n2827) );
NAND2_X1 MEM_stage_inst_dmem_U2994 ( .A1(MEM_stage_inst_dmem_ram_501), .A2(MEM_stage_inst_dmem_n3170), .ZN(MEM_stage_inst_dmem_n2825) );
NAND2_X1 MEM_stage_inst_dmem_U2993 ( .A1(MEM_stage_inst_dmem_ram_789), .A2(MEM_stage_inst_dmem_n3191), .ZN(MEM_stage_inst_dmem_n2826) );
NAND2_X1 MEM_stage_inst_dmem_U2992 ( .A1(MEM_stage_inst_dmem_n2824), .A2(MEM_stage_inst_dmem_n2823), .ZN(MEM_stage_inst_dmem_n2828) );
NAND2_X1 MEM_stage_inst_dmem_U2991 ( .A1(MEM_stage_inst_dmem_ram_933), .A2(MEM_stage_inst_dmem_n4675), .ZN(MEM_stage_inst_dmem_n2823) );
NAND2_X1 MEM_stage_inst_dmem_U2990 ( .A1(MEM_stage_inst_dmem_ram_5), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n2824) );
NOR2_X1 MEM_stage_inst_dmem_U2989 ( .A1(MEM_stage_inst_dmem_n2822), .A2(MEM_stage_inst_dmem_n2821), .ZN(MEM_stage_inst_dmem_n2830) );
NAND2_X1 MEM_stage_inst_dmem_U2988 ( .A1(MEM_stage_inst_dmem_n2820), .A2(MEM_stage_inst_dmem_n2819), .ZN(MEM_stage_inst_dmem_n2821) );
NAND2_X1 MEM_stage_inst_dmem_U2987 ( .A1(MEM_stage_inst_dmem_ram_965), .A2(MEM_stage_inst_dmem_n4728), .ZN(MEM_stage_inst_dmem_n2819) );
NAND2_X1 MEM_stage_inst_dmem_U2986 ( .A1(MEM_stage_inst_dmem_ram_693), .A2(MEM_stage_inst_dmem_n4709), .ZN(MEM_stage_inst_dmem_n2820) );
NAND2_X1 MEM_stage_inst_dmem_U2985 ( .A1(MEM_stage_inst_dmem_n2818), .A2(MEM_stage_inst_dmem_n2817), .ZN(MEM_stage_inst_dmem_n2822) );
NAND2_X1 MEM_stage_inst_dmem_U2984 ( .A1(MEM_stage_inst_dmem_ram_885), .A2(MEM_stage_inst_dmem_n3099), .ZN(MEM_stage_inst_dmem_n2817) );
NAND2_X1 MEM_stage_inst_dmem_U2983 ( .A1(MEM_stage_inst_dmem_ram_757), .A2(MEM_stage_inst_dmem_n3202), .ZN(MEM_stage_inst_dmem_n2818) );
NAND2_X1 MEM_stage_inst_dmem_U2982 ( .A1(MEM_stage_inst_dmem_n2816), .A2(MEM_stage_inst_dmem_n2815), .ZN(MEM_stage_inst_mem_read_data_4) );
NOR2_X1 MEM_stage_inst_dmem_U2981 ( .A1(MEM_stage_inst_dmem_n2814), .A2(MEM_stage_inst_dmem_n2813), .ZN(MEM_stage_inst_dmem_n2815) );
NOR2_X1 MEM_stage_inst_dmem_U2980 ( .A1(MEM_stage_inst_dmem_n2812), .A2(MEM_stage_inst_dmem_n8417), .ZN(MEM_stage_inst_dmem_n2813) );
NOR2_X1 MEM_stage_inst_dmem_U2979 ( .A1(MEM_stage_inst_dmem_n2811), .A2(MEM_stage_inst_dmem_n2810), .ZN(MEM_stage_inst_dmem_n2812) );
NAND2_X1 MEM_stage_inst_dmem_U2978 ( .A1(MEM_stage_inst_dmem_n2809), .A2(MEM_stage_inst_dmem_n2808), .ZN(MEM_stage_inst_dmem_n2810) );
NOR2_X1 MEM_stage_inst_dmem_U2977 ( .A1(MEM_stage_inst_dmem_n2807), .A2(MEM_stage_inst_dmem_n2806), .ZN(MEM_stage_inst_dmem_n2808) );
NAND2_X1 MEM_stage_inst_dmem_U2976 ( .A1(MEM_stage_inst_dmem_n2805), .A2(MEM_stage_inst_dmem_n2804), .ZN(MEM_stage_inst_dmem_n2806) );
NOR2_X1 MEM_stage_inst_dmem_U2975 ( .A1(MEM_stage_inst_dmem_n2803), .A2(MEM_stage_inst_dmem_n2802), .ZN(MEM_stage_inst_dmem_n2804) );
NAND2_X1 MEM_stage_inst_dmem_U2974 ( .A1(MEM_stage_inst_dmem_n2801), .A2(MEM_stage_inst_dmem_n2800), .ZN(MEM_stage_inst_dmem_n2802) );
NAND2_X1 MEM_stage_inst_dmem_U2973 ( .A1(MEM_stage_inst_dmem_ram_3428), .A2(MEM_stage_inst_dmem_n3217), .ZN(MEM_stage_inst_dmem_n2800) );
NAND2_X1 MEM_stage_inst_dmem_U2972 ( .A1(MEM_stage_inst_dmem_ram_3300), .A2(MEM_stage_inst_dmem_n3152), .ZN(MEM_stage_inst_dmem_n2801) );
NAND2_X1 MEM_stage_inst_dmem_U2971 ( .A1(MEM_stage_inst_dmem_n2799), .A2(MEM_stage_inst_dmem_n2798), .ZN(MEM_stage_inst_dmem_n2803) );
NAND2_X1 MEM_stage_inst_dmem_U2970 ( .A1(MEM_stage_inst_dmem_ram_3780), .A2(MEM_stage_inst_dmem_n3192), .ZN(MEM_stage_inst_dmem_n2798) );
NAND2_X1 MEM_stage_inst_dmem_U2969 ( .A1(MEM_stage_inst_dmem_ram_3492), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n2799) );
NOR2_X1 MEM_stage_inst_dmem_U2968 ( .A1(MEM_stage_inst_dmem_n2797), .A2(MEM_stage_inst_dmem_n2796), .ZN(MEM_stage_inst_dmem_n2805) );
NAND2_X1 MEM_stage_inst_dmem_U2967 ( .A1(MEM_stage_inst_dmem_n2795), .A2(MEM_stage_inst_dmem_n2794), .ZN(MEM_stage_inst_dmem_n2796) );
NAND2_X1 MEM_stage_inst_dmem_U2966 ( .A1(MEM_stage_inst_dmem_ram_3108), .A2(MEM_stage_inst_dmem_n3092), .ZN(MEM_stage_inst_dmem_n2794) );
NAND2_X1 MEM_stage_inst_dmem_U2965 ( .A1(MEM_stage_inst_dmem_ram_4084), .A2(MEM_stage_inst_dmem_n3199), .ZN(MEM_stage_inst_dmem_n2795) );
NAND2_X1 MEM_stage_inst_dmem_U2964 ( .A1(MEM_stage_inst_dmem_n2793), .A2(MEM_stage_inst_dmem_n2792), .ZN(MEM_stage_inst_dmem_n2797) );
NAND2_X1 MEM_stage_inst_dmem_U2963 ( .A1(MEM_stage_inst_dmem_ram_3204), .A2(MEM_stage_inst_dmem_n3130), .ZN(MEM_stage_inst_dmem_n2792) );
NAND2_X1 MEM_stage_inst_dmem_U2962 ( .A1(MEM_stage_inst_dmem_ram_3620), .A2(MEM_stage_inst_dmem_n4692), .ZN(MEM_stage_inst_dmem_n2793) );
NAND2_X1 MEM_stage_inst_dmem_U2961 ( .A1(MEM_stage_inst_dmem_n2791), .A2(MEM_stage_inst_dmem_n2790), .ZN(MEM_stage_inst_dmem_n2807) );
NOR2_X1 MEM_stage_inst_dmem_U2960 ( .A1(MEM_stage_inst_dmem_n2789), .A2(MEM_stage_inst_dmem_n2788), .ZN(MEM_stage_inst_dmem_n2790) );
NAND2_X1 MEM_stage_inst_dmem_U2959 ( .A1(MEM_stage_inst_dmem_n2787), .A2(MEM_stage_inst_dmem_n2786), .ZN(MEM_stage_inst_dmem_n2788) );
NAND2_X1 MEM_stage_inst_dmem_U2958 ( .A1(MEM_stage_inst_dmem_ram_3988), .A2(MEM_stage_inst_dmem_n3073), .ZN(MEM_stage_inst_dmem_n2786) );
NAND2_X1 MEM_stage_inst_dmem_U2957 ( .A1(MEM_stage_inst_dmem_ram_3796), .A2(MEM_stage_inst_dmem_n3112), .ZN(MEM_stage_inst_dmem_n2787) );
NAND2_X1 MEM_stage_inst_dmem_U2956 ( .A1(MEM_stage_inst_dmem_n2785), .A2(MEM_stage_inst_dmem_n2784), .ZN(MEM_stage_inst_dmem_n2789) );
NAND2_X1 MEM_stage_inst_dmem_U2955 ( .A1(MEM_stage_inst_dmem_ram_3348), .A2(MEM_stage_inst_dmem_n4672), .ZN(MEM_stage_inst_dmem_n2784) );
NAND2_X1 MEM_stage_inst_dmem_U2954 ( .A1(MEM_stage_inst_dmem_ram_3460), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n2785) );
NOR2_X1 MEM_stage_inst_dmem_U2953 ( .A1(MEM_stage_inst_dmem_n2783), .A2(MEM_stage_inst_dmem_n2782), .ZN(MEM_stage_inst_dmem_n2791) );
NAND2_X1 MEM_stage_inst_dmem_U2952 ( .A1(MEM_stage_inst_dmem_n2781), .A2(MEM_stage_inst_dmem_n2780), .ZN(MEM_stage_inst_dmem_n2782) );
NAND2_X1 MEM_stage_inst_dmem_U2951 ( .A1(MEM_stage_inst_dmem_ram_3956), .A2(MEM_stage_inst_dmem_n3099), .ZN(MEM_stage_inst_dmem_n2780) );
NAND2_X1 MEM_stage_inst_dmem_U2950 ( .A1(MEM_stage_inst_dmem_ram_3892), .A2(MEM_stage_inst_dmem_n4740), .ZN(MEM_stage_inst_dmem_n2781) );
NAND2_X1 MEM_stage_inst_dmem_U2949 ( .A1(MEM_stage_inst_dmem_n2779), .A2(MEM_stage_inst_dmem_n2778), .ZN(MEM_stage_inst_dmem_n2783) );
NAND2_X1 MEM_stage_inst_dmem_U2948 ( .A1(MEM_stage_inst_dmem_ram_3860), .A2(MEM_stage_inst_dmem_n3191), .ZN(MEM_stage_inst_dmem_n2778) );
NAND2_X1 MEM_stage_inst_dmem_U2947 ( .A1(MEM_stage_inst_dmem_ram_3588), .A2(MEM_stage_inst_dmem_n3182), .ZN(MEM_stage_inst_dmem_n2779) );
NOR2_X1 MEM_stage_inst_dmem_U2946 ( .A1(MEM_stage_inst_dmem_n2777), .A2(MEM_stage_inst_dmem_n2776), .ZN(MEM_stage_inst_dmem_n2809) );
NAND2_X1 MEM_stage_inst_dmem_U2945 ( .A1(MEM_stage_inst_dmem_n2775), .A2(MEM_stage_inst_dmem_n2774), .ZN(MEM_stage_inst_dmem_n2776) );
NOR2_X1 MEM_stage_inst_dmem_U2944 ( .A1(MEM_stage_inst_dmem_n2773), .A2(MEM_stage_inst_dmem_n2772), .ZN(MEM_stage_inst_dmem_n2774) );
NAND2_X1 MEM_stage_inst_dmem_U2943 ( .A1(MEM_stage_inst_dmem_n2771), .A2(MEM_stage_inst_dmem_n2770), .ZN(MEM_stage_inst_dmem_n2772) );
NAND2_X1 MEM_stage_inst_dmem_U2942 ( .A1(MEM_stage_inst_dmem_ram_3508), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n2770) );
NAND2_X1 MEM_stage_inst_dmem_U2941 ( .A1(MEM_stage_inst_dmem_ram_3284), .A2(MEM_stage_inst_dmem_n3220), .ZN(MEM_stage_inst_dmem_n2771) );
NAND2_X1 MEM_stage_inst_dmem_U2940 ( .A1(MEM_stage_inst_dmem_n2769), .A2(MEM_stage_inst_dmem_n2768), .ZN(MEM_stage_inst_dmem_n2773) );
NAND2_X1 MEM_stage_inst_dmem_U2939 ( .A1(MEM_stage_inst_dmem_ram_4020), .A2(MEM_stage_inst_dmem_n3163), .ZN(MEM_stage_inst_dmem_n2768) );
NAND2_X1 MEM_stage_inst_dmem_U2938 ( .A1(MEM_stage_inst_dmem_ram_3700), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n2769) );
NOR2_X1 MEM_stage_inst_dmem_U2937 ( .A1(MEM_stage_inst_dmem_n2767), .A2(MEM_stage_inst_dmem_n2766), .ZN(MEM_stage_inst_dmem_n2775) );
NAND2_X1 MEM_stage_inst_dmem_U2936 ( .A1(MEM_stage_inst_dmem_n2765), .A2(MEM_stage_inst_dmem_n2764), .ZN(MEM_stage_inst_dmem_n2766) );
NAND2_X1 MEM_stage_inst_dmem_U2935 ( .A1(MEM_stage_inst_dmem_ram_3636), .A2(MEM_stage_inst_dmem_n3085), .ZN(MEM_stage_inst_dmem_n2764) );
NAND2_X1 MEM_stage_inst_dmem_U2934 ( .A1(MEM_stage_inst_dmem_ram_3076), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n2765) );
NAND2_X1 MEM_stage_inst_dmem_U2933 ( .A1(MEM_stage_inst_dmem_n2763), .A2(MEM_stage_inst_dmem_n2762), .ZN(MEM_stage_inst_dmem_n2767) );
NAND2_X1 MEM_stage_inst_dmem_U2932 ( .A1(MEM_stage_inst_dmem_ram_3908), .A2(MEM_stage_inst_dmem_n3120), .ZN(MEM_stage_inst_dmem_n2762) );
NAND2_X1 MEM_stage_inst_dmem_U2931 ( .A1(MEM_stage_inst_dmem_ram_3316), .A2(MEM_stage_inst_dmem_n4649), .ZN(MEM_stage_inst_dmem_n2763) );
NAND2_X1 MEM_stage_inst_dmem_U2930 ( .A1(MEM_stage_inst_dmem_n2761), .A2(MEM_stage_inst_dmem_n2760), .ZN(MEM_stage_inst_dmem_n2777) );
NOR2_X1 MEM_stage_inst_dmem_U2929 ( .A1(MEM_stage_inst_dmem_n2759), .A2(MEM_stage_inst_dmem_n2758), .ZN(MEM_stage_inst_dmem_n2760) );
NAND2_X1 MEM_stage_inst_dmem_U2928 ( .A1(MEM_stage_inst_dmem_n2757), .A2(MEM_stage_inst_dmem_n2756), .ZN(MEM_stage_inst_dmem_n2758) );
NAND2_X1 MEM_stage_inst_dmem_U2927 ( .A1(MEM_stage_inst_dmem_ram_3092), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n2756) );
NAND2_X1 MEM_stage_inst_dmem_U2926 ( .A1(MEM_stage_inst_dmem_ram_3412), .A2(MEM_stage_inst_dmem_n3216), .ZN(MEM_stage_inst_dmem_n2757) );
NAND2_X1 MEM_stage_inst_dmem_U2925 ( .A1(MEM_stage_inst_dmem_n2755), .A2(MEM_stage_inst_dmem_n2754), .ZN(MEM_stage_inst_dmem_n2759) );
NAND2_X1 MEM_stage_inst_dmem_U2924 ( .A1(MEM_stage_inst_dmem_ram_3876), .A2(MEM_stage_inst_dmem_n3137), .ZN(MEM_stage_inst_dmem_n2754) );
NAND2_X1 MEM_stage_inst_dmem_U2923 ( .A1(MEM_stage_inst_dmem_ram_3172), .A2(MEM_stage_inst_dmem_n3179), .ZN(MEM_stage_inst_dmem_n2755) );
NOR2_X1 MEM_stage_inst_dmem_U2922 ( .A1(MEM_stage_inst_dmem_n2753), .A2(MEM_stage_inst_dmem_n2752), .ZN(MEM_stage_inst_dmem_n2761) );
NAND2_X1 MEM_stage_inst_dmem_U2921 ( .A1(MEM_stage_inst_dmem_n2751), .A2(MEM_stage_inst_dmem_n2750), .ZN(MEM_stage_inst_dmem_n2752) );
NAND2_X1 MEM_stage_inst_dmem_U2920 ( .A1(MEM_stage_inst_dmem_ram_3572), .A2(MEM_stage_inst_dmem_n3170), .ZN(MEM_stage_inst_dmem_n2750) );
NAND2_X1 MEM_stage_inst_dmem_U2919 ( .A1(MEM_stage_inst_dmem_ram_3540), .A2(MEM_stage_inst_dmem_n3174), .ZN(MEM_stage_inst_dmem_n2751) );
NAND2_X1 MEM_stage_inst_dmem_U2918 ( .A1(MEM_stage_inst_dmem_n2749), .A2(MEM_stage_inst_dmem_n2748), .ZN(MEM_stage_inst_dmem_n2753) );
NAND2_X1 MEM_stage_inst_dmem_U2917 ( .A1(MEM_stage_inst_dmem_ram_3124), .A2(MEM_stage_inst_dmem_n3103), .ZN(MEM_stage_inst_dmem_n2748) );
NAND2_X1 MEM_stage_inst_dmem_U2916 ( .A1(MEM_stage_inst_dmem_ram_3236), .A2(MEM_stage_inst_dmem_n3081), .ZN(MEM_stage_inst_dmem_n2749) );
NAND2_X1 MEM_stage_inst_dmem_U2915 ( .A1(MEM_stage_inst_dmem_n2747), .A2(MEM_stage_inst_dmem_n2746), .ZN(MEM_stage_inst_dmem_n2811) );
NOR2_X1 MEM_stage_inst_dmem_U2914 ( .A1(MEM_stage_inst_dmem_n2745), .A2(MEM_stage_inst_dmem_n2744), .ZN(MEM_stage_inst_dmem_n2746) );
NAND2_X1 MEM_stage_inst_dmem_U2913 ( .A1(MEM_stage_inst_dmem_n2743), .A2(MEM_stage_inst_dmem_n2742), .ZN(MEM_stage_inst_dmem_n2744) );
NOR2_X1 MEM_stage_inst_dmem_U2912 ( .A1(MEM_stage_inst_dmem_n2741), .A2(MEM_stage_inst_dmem_n2740), .ZN(MEM_stage_inst_dmem_n2742) );
NAND2_X1 MEM_stage_inst_dmem_U2911 ( .A1(MEM_stage_inst_dmem_n2739), .A2(MEM_stage_inst_dmem_n2738), .ZN(MEM_stage_inst_dmem_n2740) );
NAND2_X1 MEM_stage_inst_dmem_U2910 ( .A1(MEM_stage_inst_dmem_ram_3764), .A2(MEM_stage_inst_dmem_n4709), .ZN(MEM_stage_inst_dmem_n2738) );
NAND2_X1 MEM_stage_inst_dmem_U2909 ( .A1(MEM_stage_inst_dmem_ram_3524), .A2(MEM_stage_inst_dmem_n3173), .ZN(MEM_stage_inst_dmem_n2739) );
NAND2_X1 MEM_stage_inst_dmem_U2908 ( .A1(MEM_stage_inst_dmem_n2737), .A2(MEM_stage_inst_dmem_n2736), .ZN(MEM_stage_inst_dmem_n2741) );
NAND2_X1 MEM_stage_inst_dmem_U2907 ( .A1(MEM_stage_inst_dmem_ram_3940), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n2736) );
NAND2_X1 MEM_stage_inst_dmem_U2906 ( .A1(MEM_stage_inst_dmem_ram_3140), .A2(MEM_stage_inst_dmem_n3102), .ZN(MEM_stage_inst_dmem_n2737) );
NOR2_X1 MEM_stage_inst_dmem_U2905 ( .A1(MEM_stage_inst_dmem_n2735), .A2(MEM_stage_inst_dmem_n2734), .ZN(MEM_stage_inst_dmem_n2743) );
NAND2_X1 MEM_stage_inst_dmem_U2904 ( .A1(MEM_stage_inst_dmem_n2733), .A2(MEM_stage_inst_dmem_n2732), .ZN(MEM_stage_inst_dmem_n2734) );
NAND2_X1 MEM_stage_inst_dmem_U2903 ( .A1(MEM_stage_inst_dmem_ram_3972), .A2(MEM_stage_inst_dmem_n3123), .ZN(MEM_stage_inst_dmem_n2732) );
NAND2_X1 MEM_stage_inst_dmem_U2902 ( .A1(MEM_stage_inst_dmem_ram_3732), .A2(MEM_stage_inst_dmem_n3076), .ZN(MEM_stage_inst_dmem_n2733) );
NAND2_X1 MEM_stage_inst_dmem_U2901 ( .A1(MEM_stage_inst_dmem_n2731), .A2(MEM_stage_inst_dmem_n2730), .ZN(MEM_stage_inst_dmem_n2735) );
NAND2_X1 MEM_stage_inst_dmem_U2900 ( .A1(MEM_stage_inst_dmem_ram_4036), .A2(MEM_stage_inst_dmem_n4728), .ZN(MEM_stage_inst_dmem_n2730) );
NAND2_X1 MEM_stage_inst_dmem_U2899 ( .A1(MEM_stage_inst_dmem_ram_3652), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n2731) );
NAND2_X1 MEM_stage_inst_dmem_U2898 ( .A1(MEM_stage_inst_dmem_n2729), .A2(MEM_stage_inst_dmem_n2728), .ZN(MEM_stage_inst_dmem_n2745) );
NOR2_X1 MEM_stage_inst_dmem_U2897 ( .A1(MEM_stage_inst_dmem_n2727), .A2(MEM_stage_inst_dmem_n2726), .ZN(MEM_stage_inst_dmem_n2728) );
NAND2_X1 MEM_stage_inst_dmem_U2896 ( .A1(MEM_stage_inst_dmem_n2725), .A2(MEM_stage_inst_dmem_n2724), .ZN(MEM_stage_inst_dmem_n2726) );
NAND2_X1 MEM_stage_inst_dmem_U2895 ( .A1(MEM_stage_inst_dmem_ram_3844), .A2(MEM_stage_inst_dmem_n37), .ZN(MEM_stage_inst_dmem_n2724) );
NAND2_X1 MEM_stage_inst_dmem_U2894 ( .A1(MEM_stage_inst_dmem_ram_3220), .A2(MEM_stage_inst_dmem_n44), .ZN(MEM_stage_inst_dmem_n2725) );
NAND2_X1 MEM_stage_inst_dmem_U2893 ( .A1(MEM_stage_inst_dmem_n2723), .A2(MEM_stage_inst_dmem_n2722), .ZN(MEM_stage_inst_dmem_n2727) );
NAND2_X1 MEM_stage_inst_dmem_U2892 ( .A1(MEM_stage_inst_dmem_ram_3476), .A2(MEM_stage_inst_dmem_n3160), .ZN(MEM_stage_inst_dmem_n2722) );
NAND2_X1 MEM_stage_inst_dmem_U2891 ( .A1(MEM_stage_inst_dmem_ram_3748), .A2(MEM_stage_inst_dmem_n3155), .ZN(MEM_stage_inst_dmem_n2723) );
NOR2_X1 MEM_stage_inst_dmem_U2890 ( .A1(MEM_stage_inst_dmem_n2721), .A2(MEM_stage_inst_dmem_n2720), .ZN(MEM_stage_inst_dmem_n2729) );
NAND2_X1 MEM_stage_inst_dmem_U2889 ( .A1(MEM_stage_inst_dmem_n2719), .A2(MEM_stage_inst_dmem_n2718), .ZN(MEM_stage_inst_dmem_n2720) );
NAND2_X1 MEM_stage_inst_dmem_U2888 ( .A1(MEM_stage_inst_dmem_ram_3364), .A2(MEM_stage_inst_dmem_n3209), .ZN(MEM_stage_inst_dmem_n2718) );
NAND2_X1 MEM_stage_inst_dmem_U2887 ( .A1(MEM_stage_inst_dmem_ram_3668), .A2(MEM_stage_inst_dmem_n3140), .ZN(MEM_stage_inst_dmem_n2719) );
NAND2_X1 MEM_stage_inst_dmem_U2886 ( .A1(MEM_stage_inst_dmem_n2717), .A2(MEM_stage_inst_dmem_n2716), .ZN(MEM_stage_inst_dmem_n2721) );
NAND2_X1 MEM_stage_inst_dmem_U2885 ( .A1(MEM_stage_inst_dmem_ram_3924), .A2(MEM_stage_inst_dmem_n3141), .ZN(MEM_stage_inst_dmem_n2716) );
NAND2_X1 MEM_stage_inst_dmem_U2884 ( .A1(MEM_stage_inst_dmem_ram_3828), .A2(MEM_stage_inst_dmem_n3202), .ZN(MEM_stage_inst_dmem_n2717) );
NOR2_X1 MEM_stage_inst_dmem_U2883 ( .A1(MEM_stage_inst_dmem_n2715), .A2(MEM_stage_inst_dmem_n2714), .ZN(MEM_stage_inst_dmem_n2747) );
NAND2_X1 MEM_stage_inst_dmem_U2882 ( .A1(MEM_stage_inst_dmem_n2713), .A2(MEM_stage_inst_dmem_n2712), .ZN(MEM_stage_inst_dmem_n2714) );
NOR2_X1 MEM_stage_inst_dmem_U2881 ( .A1(MEM_stage_inst_dmem_n2711), .A2(MEM_stage_inst_dmem_n2710), .ZN(MEM_stage_inst_dmem_n2712) );
NAND2_X1 MEM_stage_inst_dmem_U2880 ( .A1(MEM_stage_inst_dmem_n2709), .A2(MEM_stage_inst_dmem_n2708), .ZN(MEM_stage_inst_dmem_n2710) );
NAND2_X1 MEM_stage_inst_dmem_U2879 ( .A1(MEM_stage_inst_dmem_ram_3268), .A2(MEM_stage_inst_dmem_n3082), .ZN(MEM_stage_inst_dmem_n2708) );
NAND2_X1 MEM_stage_inst_dmem_U2878 ( .A1(MEM_stage_inst_dmem_ram_3812), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n2709) );
NAND2_X1 MEM_stage_inst_dmem_U2877 ( .A1(MEM_stage_inst_dmem_n2707), .A2(MEM_stage_inst_dmem_n2706), .ZN(MEM_stage_inst_dmem_n2711) );
NAND2_X1 MEM_stage_inst_dmem_U2876 ( .A1(MEM_stage_inst_dmem_ram_4068), .A2(MEM_stage_inst_dmem_n3113), .ZN(MEM_stage_inst_dmem_n2706) );
NAND2_X1 MEM_stage_inst_dmem_U2875 ( .A1(MEM_stage_inst_dmem_ram_4004), .A2(MEM_stage_inst_dmem_n4675), .ZN(MEM_stage_inst_dmem_n2707) );
NOR2_X1 MEM_stage_inst_dmem_U2874 ( .A1(MEM_stage_inst_dmem_n2705), .A2(MEM_stage_inst_dmem_n2704), .ZN(MEM_stage_inst_dmem_n2713) );
NAND2_X1 MEM_stage_inst_dmem_U2873 ( .A1(MEM_stage_inst_dmem_n2703), .A2(MEM_stage_inst_dmem_n2702), .ZN(MEM_stage_inst_dmem_n2704) );
NAND2_X1 MEM_stage_inst_dmem_U2872 ( .A1(MEM_stage_inst_dmem_ram_3380), .A2(MEM_stage_inst_dmem_n4731), .ZN(MEM_stage_inst_dmem_n2702) );
NAND2_X1 MEM_stage_inst_dmem_U2871 ( .A1(MEM_stage_inst_dmem_ram_3604), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n2703) );
NAND2_X1 MEM_stage_inst_dmem_U2870 ( .A1(MEM_stage_inst_dmem_n2701), .A2(MEM_stage_inst_dmem_n2700), .ZN(MEM_stage_inst_dmem_n2705) );
NAND2_X1 MEM_stage_inst_dmem_U2869 ( .A1(MEM_stage_inst_dmem_ram_3156), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n2700) );
NAND2_X1 MEM_stage_inst_dmem_U2868 ( .A1(MEM_stage_inst_dmem_ram_3332), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n2701) );
NAND2_X1 MEM_stage_inst_dmem_U2867 ( .A1(MEM_stage_inst_dmem_n2699), .A2(MEM_stage_inst_dmem_n2698), .ZN(MEM_stage_inst_dmem_n2715) );
NOR2_X1 MEM_stage_inst_dmem_U2866 ( .A1(MEM_stage_inst_dmem_n2697), .A2(MEM_stage_inst_dmem_n2696), .ZN(MEM_stage_inst_dmem_n2698) );
NAND2_X1 MEM_stage_inst_dmem_U2865 ( .A1(MEM_stage_inst_dmem_n2695), .A2(MEM_stage_inst_dmem_n2694), .ZN(MEM_stage_inst_dmem_n2696) );
NAND2_X1 MEM_stage_inst_dmem_U2864 ( .A1(MEM_stage_inst_dmem_ram_4052), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n2694) );
NAND2_X1 MEM_stage_inst_dmem_U2863 ( .A1(MEM_stage_inst_dmem_ram_3252), .A2(MEM_stage_inst_dmem_n55), .ZN(MEM_stage_inst_dmem_n2695) );
NAND2_X1 MEM_stage_inst_dmem_U2862 ( .A1(MEM_stage_inst_dmem_n2693), .A2(MEM_stage_inst_dmem_n2692), .ZN(MEM_stage_inst_dmem_n2697) );
NAND2_X1 MEM_stage_inst_dmem_U2861 ( .A1(MEM_stage_inst_dmem_ram_3684), .A2(MEM_stage_inst_dmem_n4701), .ZN(MEM_stage_inst_dmem_n2692) );
NAND2_X1 MEM_stage_inst_dmem_U2860 ( .A1(MEM_stage_inst_dmem_ram_3444), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n2693) );
NOR2_X1 MEM_stage_inst_dmem_U2859 ( .A1(MEM_stage_inst_dmem_n2691), .A2(MEM_stage_inst_dmem_n2690), .ZN(MEM_stage_inst_dmem_n2699) );
NAND2_X1 MEM_stage_inst_dmem_U2858 ( .A1(MEM_stage_inst_dmem_n2689), .A2(MEM_stage_inst_dmem_n2688), .ZN(MEM_stage_inst_dmem_n2690) );
NAND2_X1 MEM_stage_inst_dmem_U2857 ( .A1(MEM_stage_inst_dmem_ram_3716), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n2688) );
NAND2_X1 MEM_stage_inst_dmem_U2856 ( .A1(MEM_stage_inst_dmem_ram_3188), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n2689) );
NAND2_X1 MEM_stage_inst_dmem_U2855 ( .A1(MEM_stage_inst_dmem_n2687), .A2(MEM_stage_inst_dmem_n2686), .ZN(MEM_stage_inst_dmem_n2691) );
NAND2_X1 MEM_stage_inst_dmem_U2854 ( .A1(MEM_stage_inst_dmem_ram_3396), .A2(MEM_stage_inst_dmem_n4706), .ZN(MEM_stage_inst_dmem_n2686) );
NAND2_X1 MEM_stage_inst_dmem_U2853 ( .A1(MEM_stage_inst_dmem_ram_3556), .A2(MEM_stage_inst_dmem_n4667), .ZN(MEM_stage_inst_dmem_n2687) );
NOR2_X1 MEM_stage_inst_dmem_U2852 ( .A1(MEM_stage_inst_dmem_n2685), .A2(MEM_stage_inst_dmem_n8152), .ZN(MEM_stage_inst_dmem_n2814) );
NOR2_X1 MEM_stage_inst_dmem_U2851 ( .A1(MEM_stage_inst_dmem_n2684), .A2(MEM_stage_inst_dmem_n2683), .ZN(MEM_stage_inst_dmem_n2685) );
NAND2_X1 MEM_stage_inst_dmem_U2850 ( .A1(MEM_stage_inst_dmem_n2682), .A2(MEM_stage_inst_dmem_n2681), .ZN(MEM_stage_inst_dmem_n2683) );
NOR2_X1 MEM_stage_inst_dmem_U2849 ( .A1(MEM_stage_inst_dmem_n2680), .A2(MEM_stage_inst_dmem_n2679), .ZN(MEM_stage_inst_dmem_n2681) );
NAND2_X1 MEM_stage_inst_dmem_U2848 ( .A1(MEM_stage_inst_dmem_n2678), .A2(MEM_stage_inst_dmem_n2677), .ZN(MEM_stage_inst_dmem_n2679) );
NOR2_X1 MEM_stage_inst_dmem_U2847 ( .A1(MEM_stage_inst_dmem_n2676), .A2(MEM_stage_inst_dmem_n2675), .ZN(MEM_stage_inst_dmem_n2677) );
NAND2_X1 MEM_stage_inst_dmem_U2846 ( .A1(MEM_stage_inst_dmem_n2674), .A2(MEM_stage_inst_dmem_n2673), .ZN(MEM_stage_inst_dmem_n2675) );
NAND2_X1 MEM_stage_inst_dmem_U2845 ( .A1(MEM_stage_inst_dmem_ram_1524), .A2(MEM_stage_inst_dmem_n3170), .ZN(MEM_stage_inst_dmem_n2673) );
NAND2_X1 MEM_stage_inst_dmem_U2844 ( .A1(MEM_stage_inst_dmem_ram_1140), .A2(MEM_stage_inst_dmem_n4710), .ZN(MEM_stage_inst_dmem_n2674) );
NAND2_X1 MEM_stage_inst_dmem_U2843 ( .A1(MEM_stage_inst_dmem_n2672), .A2(MEM_stage_inst_dmem_n2671), .ZN(MEM_stage_inst_dmem_n2676) );
NAND2_X1 MEM_stage_inst_dmem_U2842 ( .A1(MEM_stage_inst_dmem_ram_1156), .A2(MEM_stage_inst_dmem_n3130), .ZN(MEM_stage_inst_dmem_n2671) );
NAND2_X1 MEM_stage_inst_dmem_U2841 ( .A1(MEM_stage_inst_dmem_ram_1060), .A2(MEM_stage_inst_dmem_n3092), .ZN(MEM_stage_inst_dmem_n2672) );
NOR2_X1 MEM_stage_inst_dmem_U2840 ( .A1(MEM_stage_inst_dmem_n2670), .A2(MEM_stage_inst_dmem_n2669), .ZN(MEM_stage_inst_dmem_n2678) );
NAND2_X1 MEM_stage_inst_dmem_U2839 ( .A1(MEM_stage_inst_dmem_n2668), .A2(MEM_stage_inst_dmem_n2667), .ZN(MEM_stage_inst_dmem_n2669) );
NAND2_X1 MEM_stage_inst_dmem_U2838 ( .A1(MEM_stage_inst_dmem_ram_1348), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n2667) );
NAND2_X1 MEM_stage_inst_dmem_U2837 ( .A1(MEM_stage_inst_dmem_ram_1924), .A2(MEM_stage_inst_dmem_n3123), .ZN(MEM_stage_inst_dmem_n2668) );
NAND2_X1 MEM_stage_inst_dmem_U2836 ( .A1(MEM_stage_inst_dmem_n2666), .A2(MEM_stage_inst_dmem_n2665), .ZN(MEM_stage_inst_dmem_n2670) );
NAND2_X1 MEM_stage_inst_dmem_U2835 ( .A1(MEM_stage_inst_dmem_ram_1908), .A2(MEM_stage_inst_dmem_n3099), .ZN(MEM_stage_inst_dmem_n2665) );
NAND2_X1 MEM_stage_inst_dmem_U2834 ( .A1(MEM_stage_inst_dmem_ram_1956), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n2666) );
NAND2_X1 MEM_stage_inst_dmem_U2833 ( .A1(MEM_stage_inst_dmem_n2664), .A2(MEM_stage_inst_dmem_n2663), .ZN(MEM_stage_inst_dmem_n2680) );
NOR2_X1 MEM_stage_inst_dmem_U2832 ( .A1(MEM_stage_inst_dmem_n2662), .A2(MEM_stage_inst_dmem_n2661), .ZN(MEM_stage_inst_dmem_n2663) );
NAND2_X1 MEM_stage_inst_dmem_U2831 ( .A1(MEM_stage_inst_dmem_n2660), .A2(MEM_stage_inst_dmem_n2659), .ZN(MEM_stage_inst_dmem_n2661) );
NAND2_X1 MEM_stage_inst_dmem_U2830 ( .A1(MEM_stage_inst_dmem_ram_1236), .A2(MEM_stage_inst_dmem_n3220), .ZN(MEM_stage_inst_dmem_n2659) );
NAND2_X1 MEM_stage_inst_dmem_U2829 ( .A1(MEM_stage_inst_dmem_ram_1204), .A2(MEM_stage_inst_dmem_n55), .ZN(MEM_stage_inst_dmem_n2660) );
NAND2_X1 MEM_stage_inst_dmem_U2828 ( .A1(MEM_stage_inst_dmem_n2658), .A2(MEM_stage_inst_dmem_n2657), .ZN(MEM_stage_inst_dmem_n2662) );
NAND2_X1 MEM_stage_inst_dmem_U2827 ( .A1(MEM_stage_inst_dmem_ram_1636), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n2657) );
NAND2_X1 MEM_stage_inst_dmem_U2826 ( .A1(MEM_stage_inst_dmem_ram_1812), .A2(MEM_stage_inst_dmem_n3191), .ZN(MEM_stage_inst_dmem_n2658) );
NOR2_X1 MEM_stage_inst_dmem_U2825 ( .A1(MEM_stage_inst_dmem_n2656), .A2(MEM_stage_inst_dmem_n2655), .ZN(MEM_stage_inst_dmem_n2664) );
NAND2_X1 MEM_stage_inst_dmem_U2824 ( .A1(MEM_stage_inst_dmem_n2654), .A2(MEM_stage_inst_dmem_n2653), .ZN(MEM_stage_inst_dmem_n2655) );
NAND2_X1 MEM_stage_inst_dmem_U2823 ( .A1(MEM_stage_inst_dmem_ram_1860), .A2(MEM_stage_inst_dmem_n3120), .ZN(MEM_stage_inst_dmem_n2653) );
NAND2_X1 MEM_stage_inst_dmem_U2822 ( .A1(MEM_stage_inst_dmem_ram_1300), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n2654) );
NAND2_X1 MEM_stage_inst_dmem_U2821 ( .A1(MEM_stage_inst_dmem_n2652), .A2(MEM_stage_inst_dmem_n2651), .ZN(MEM_stage_inst_dmem_n2656) );
NAND2_X1 MEM_stage_inst_dmem_U2820 ( .A1(MEM_stage_inst_dmem_ram_1620), .A2(MEM_stage_inst_dmem_n3140), .ZN(MEM_stage_inst_dmem_n2651) );
NAND2_X1 MEM_stage_inst_dmem_U2819 ( .A1(MEM_stage_inst_dmem_ram_1748), .A2(MEM_stage_inst_dmem_n3112), .ZN(MEM_stage_inst_dmem_n2652) );
NOR2_X1 MEM_stage_inst_dmem_U2818 ( .A1(MEM_stage_inst_dmem_n2650), .A2(MEM_stage_inst_dmem_n2649), .ZN(MEM_stage_inst_dmem_n2682) );
NAND2_X1 MEM_stage_inst_dmem_U2817 ( .A1(MEM_stage_inst_dmem_n2648), .A2(MEM_stage_inst_dmem_n2647), .ZN(MEM_stage_inst_dmem_n2649) );
NOR2_X1 MEM_stage_inst_dmem_U2816 ( .A1(MEM_stage_inst_dmem_n2646), .A2(MEM_stage_inst_dmem_n2645), .ZN(MEM_stage_inst_dmem_n2647) );
NAND2_X1 MEM_stage_inst_dmem_U2815 ( .A1(MEM_stage_inst_dmem_n2644), .A2(MEM_stage_inst_dmem_n2643), .ZN(MEM_stage_inst_dmem_n2645) );
NAND2_X1 MEM_stage_inst_dmem_U2814 ( .A1(MEM_stage_inst_dmem_ram_1668), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n2643) );
NAND2_X1 MEM_stage_inst_dmem_U2813 ( .A1(MEM_stage_inst_dmem_ram_1316), .A2(MEM_stage_inst_dmem_n3209), .ZN(MEM_stage_inst_dmem_n2644) );
NAND2_X1 MEM_stage_inst_dmem_U2812 ( .A1(MEM_stage_inst_dmem_n2642), .A2(MEM_stage_inst_dmem_n2641), .ZN(MEM_stage_inst_dmem_n2646) );
NAND2_X1 MEM_stage_inst_dmem_U2811 ( .A1(MEM_stage_inst_dmem_ram_1220), .A2(MEM_stage_inst_dmem_n3082), .ZN(MEM_stage_inst_dmem_n2641) );
NAND2_X1 MEM_stage_inst_dmem_U2810 ( .A1(MEM_stage_inst_dmem_ram_1332), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n2642) );
NOR2_X1 MEM_stage_inst_dmem_U2809 ( .A1(MEM_stage_inst_dmem_n2640), .A2(MEM_stage_inst_dmem_n2639), .ZN(MEM_stage_inst_dmem_n2648) );
NAND2_X1 MEM_stage_inst_dmem_U2808 ( .A1(MEM_stage_inst_dmem_n2638), .A2(MEM_stage_inst_dmem_n2637), .ZN(MEM_stage_inst_dmem_n2639) );
NAND2_X1 MEM_stage_inst_dmem_U2807 ( .A1(MEM_stage_inst_dmem_ram_1428), .A2(MEM_stage_inst_dmem_n3160), .ZN(MEM_stage_inst_dmem_n2637) );
NAND2_X1 MEM_stage_inst_dmem_U2806 ( .A1(MEM_stage_inst_dmem_ram_2036), .A2(MEM_stage_inst_dmem_n3199), .ZN(MEM_stage_inst_dmem_n2638) );
NAND2_X1 MEM_stage_inst_dmem_U2805 ( .A1(MEM_stage_inst_dmem_n2636), .A2(MEM_stage_inst_dmem_n2635), .ZN(MEM_stage_inst_dmem_n2640) );
NAND2_X1 MEM_stage_inst_dmem_U2804 ( .A1(MEM_stage_inst_dmem_ram_1892), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n2635) );
NAND2_X1 MEM_stage_inst_dmem_U2803 ( .A1(MEM_stage_inst_dmem_ram_1844), .A2(MEM_stage_inst_dmem_n46), .ZN(MEM_stage_inst_dmem_n2636) );
NAND2_X1 MEM_stage_inst_dmem_U2802 ( .A1(MEM_stage_inst_dmem_n2634), .A2(MEM_stage_inst_dmem_n2633), .ZN(MEM_stage_inst_dmem_n2650) );
NOR2_X1 MEM_stage_inst_dmem_U2801 ( .A1(MEM_stage_inst_dmem_n2632), .A2(MEM_stage_inst_dmem_n2631), .ZN(MEM_stage_inst_dmem_n2633) );
NAND2_X1 MEM_stage_inst_dmem_U2800 ( .A1(MEM_stage_inst_dmem_n2630), .A2(MEM_stage_inst_dmem_n2629), .ZN(MEM_stage_inst_dmem_n2631) );
NAND2_X1 MEM_stage_inst_dmem_U2799 ( .A1(MEM_stage_inst_dmem_ram_1076), .A2(MEM_stage_inst_dmem_n3103), .ZN(MEM_stage_inst_dmem_n2629) );
NAND2_X1 MEM_stage_inst_dmem_U2798 ( .A1(MEM_stage_inst_dmem_ram_1972), .A2(MEM_stage_inst_dmem_n3163), .ZN(MEM_stage_inst_dmem_n2630) );
NAND2_X1 MEM_stage_inst_dmem_U2797 ( .A1(MEM_stage_inst_dmem_n2628), .A2(MEM_stage_inst_dmem_n2627), .ZN(MEM_stage_inst_dmem_n2632) );
NAND2_X1 MEM_stage_inst_dmem_U2796 ( .A1(MEM_stage_inst_dmem_ram_1092), .A2(MEM_stage_inst_dmem_n3102), .ZN(MEM_stage_inst_dmem_n2627) );
NAND2_X1 MEM_stage_inst_dmem_U2795 ( .A1(MEM_stage_inst_dmem_ram_1828), .A2(MEM_stage_inst_dmem_n3137), .ZN(MEM_stage_inst_dmem_n2628) );
NOR2_X1 MEM_stage_inst_dmem_U2794 ( .A1(MEM_stage_inst_dmem_n2626), .A2(MEM_stage_inst_dmem_n2625), .ZN(MEM_stage_inst_dmem_n2634) );
NAND2_X1 MEM_stage_inst_dmem_U2793 ( .A1(MEM_stage_inst_dmem_n2624), .A2(MEM_stage_inst_dmem_n2623), .ZN(MEM_stage_inst_dmem_n2625) );
NAND2_X1 MEM_stage_inst_dmem_U2792 ( .A1(MEM_stage_inst_dmem_ram_1876), .A2(MEM_stage_inst_dmem_n3141), .ZN(MEM_stage_inst_dmem_n2623) );
NAND2_X1 MEM_stage_inst_dmem_U2791 ( .A1(MEM_stage_inst_dmem_ram_1940), .A2(MEM_stage_inst_dmem_n3073), .ZN(MEM_stage_inst_dmem_n2624) );
NAND2_X1 MEM_stage_inst_dmem_U2790 ( .A1(MEM_stage_inst_dmem_n2622), .A2(MEM_stage_inst_dmem_n2621), .ZN(MEM_stage_inst_dmem_n2626) );
NAND2_X1 MEM_stage_inst_dmem_U2789 ( .A1(MEM_stage_inst_dmem_ram_2004), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n2621) );
NAND2_X1 MEM_stage_inst_dmem_U2788 ( .A1(MEM_stage_inst_dmem_ram_1764), .A2(MEM_stage_inst_dmem_n4769), .ZN(MEM_stage_inst_dmem_n2622) );
NAND2_X1 MEM_stage_inst_dmem_U2787 ( .A1(MEM_stage_inst_dmem_n2620), .A2(MEM_stage_inst_dmem_n2619), .ZN(MEM_stage_inst_dmem_n2684) );
NOR2_X1 MEM_stage_inst_dmem_U2786 ( .A1(MEM_stage_inst_dmem_n2618), .A2(MEM_stage_inst_dmem_n2617), .ZN(MEM_stage_inst_dmem_n2619) );
NAND2_X1 MEM_stage_inst_dmem_U2785 ( .A1(MEM_stage_inst_dmem_n2616), .A2(MEM_stage_inst_dmem_n2615), .ZN(MEM_stage_inst_dmem_n2617) );
NOR2_X1 MEM_stage_inst_dmem_U2784 ( .A1(MEM_stage_inst_dmem_n2614), .A2(MEM_stage_inst_dmem_n2613), .ZN(MEM_stage_inst_dmem_n2615) );
NAND2_X1 MEM_stage_inst_dmem_U2783 ( .A1(MEM_stage_inst_dmem_n2612), .A2(MEM_stage_inst_dmem_n2611), .ZN(MEM_stage_inst_dmem_n2613) );
NAND2_X1 MEM_stage_inst_dmem_U2782 ( .A1(MEM_stage_inst_dmem_ram_1444), .A2(MEM_stage_inst_dmem_n4772), .ZN(MEM_stage_inst_dmem_n2611) );
NAND2_X1 MEM_stage_inst_dmem_U2781 ( .A1(MEM_stage_inst_dmem_ram_1540), .A2(MEM_stage_inst_dmem_n3182), .ZN(MEM_stage_inst_dmem_n2612) );
NAND2_X1 MEM_stage_inst_dmem_U2780 ( .A1(MEM_stage_inst_dmem_n2610), .A2(MEM_stage_inst_dmem_n2609), .ZN(MEM_stage_inst_dmem_n2614) );
NAND2_X1 MEM_stage_inst_dmem_U2779 ( .A1(MEM_stage_inst_dmem_ram_1732), .A2(MEM_stage_inst_dmem_n3192), .ZN(MEM_stage_inst_dmem_n2609) );
NAND2_X1 MEM_stage_inst_dmem_U2778 ( .A1(MEM_stage_inst_dmem_ram_1716), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n2610) );
NOR2_X1 MEM_stage_inst_dmem_U2777 ( .A1(MEM_stage_inst_dmem_n2608), .A2(MEM_stage_inst_dmem_n2607), .ZN(MEM_stage_inst_dmem_n2616) );
NAND2_X1 MEM_stage_inst_dmem_U2776 ( .A1(MEM_stage_inst_dmem_n2606), .A2(MEM_stage_inst_dmem_n2605), .ZN(MEM_stage_inst_dmem_n2607) );
NAND2_X1 MEM_stage_inst_dmem_U2775 ( .A1(MEM_stage_inst_dmem_ram_1588), .A2(MEM_stage_inst_dmem_n3085), .ZN(MEM_stage_inst_dmem_n2605) );
NAND2_X1 MEM_stage_inst_dmem_U2774 ( .A1(MEM_stage_inst_dmem_ram_1028), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n2606) );
NAND2_X1 MEM_stage_inst_dmem_U2773 ( .A1(MEM_stage_inst_dmem_n2604), .A2(MEM_stage_inst_dmem_n2603), .ZN(MEM_stage_inst_dmem_n2608) );
NAND2_X1 MEM_stage_inst_dmem_U2772 ( .A1(MEM_stage_inst_dmem_ram_1380), .A2(MEM_stage_inst_dmem_n3217), .ZN(MEM_stage_inst_dmem_n2603) );
NAND2_X1 MEM_stage_inst_dmem_U2771 ( .A1(MEM_stage_inst_dmem_ram_1364), .A2(MEM_stage_inst_dmem_n3216), .ZN(MEM_stage_inst_dmem_n2604) );
NAND2_X1 MEM_stage_inst_dmem_U2770 ( .A1(MEM_stage_inst_dmem_n2602), .A2(MEM_stage_inst_dmem_n2601), .ZN(MEM_stage_inst_dmem_n2618) );
NOR2_X1 MEM_stage_inst_dmem_U2769 ( .A1(MEM_stage_inst_dmem_n2600), .A2(MEM_stage_inst_dmem_n2599), .ZN(MEM_stage_inst_dmem_n2601) );
NAND2_X1 MEM_stage_inst_dmem_U2768 ( .A1(MEM_stage_inst_dmem_n2598), .A2(MEM_stage_inst_dmem_n2597), .ZN(MEM_stage_inst_dmem_n2599) );
NAND2_X1 MEM_stage_inst_dmem_U2767 ( .A1(MEM_stage_inst_dmem_ram_2020), .A2(MEM_stage_inst_dmem_n3113), .ZN(MEM_stage_inst_dmem_n2597) );
NAND2_X1 MEM_stage_inst_dmem_U2766 ( .A1(MEM_stage_inst_dmem_ram_1572), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n2598) );
NAND2_X1 MEM_stage_inst_dmem_U2765 ( .A1(MEM_stage_inst_dmem_n2596), .A2(MEM_stage_inst_dmem_n2595), .ZN(MEM_stage_inst_dmem_n2600) );
NAND2_X1 MEM_stage_inst_dmem_U2764 ( .A1(MEM_stage_inst_dmem_ram_1460), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n2595) );
NAND2_X1 MEM_stage_inst_dmem_U2763 ( .A1(MEM_stage_inst_dmem_ram_1044), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n2596) );
NOR2_X1 MEM_stage_inst_dmem_U2762 ( .A1(MEM_stage_inst_dmem_n2594), .A2(MEM_stage_inst_dmem_n2593), .ZN(MEM_stage_inst_dmem_n2602) );
NAND2_X1 MEM_stage_inst_dmem_U2761 ( .A1(MEM_stage_inst_dmem_n2592), .A2(MEM_stage_inst_dmem_n2591), .ZN(MEM_stage_inst_dmem_n2593) );
NAND2_X1 MEM_stage_inst_dmem_U2760 ( .A1(MEM_stage_inst_dmem_ram_1796), .A2(MEM_stage_inst_dmem_n37), .ZN(MEM_stage_inst_dmem_n2591) );
NAND2_X1 MEM_stage_inst_dmem_U2759 ( .A1(MEM_stage_inst_dmem_ram_1396), .A2(MEM_stage_inst_dmem_n4721), .ZN(MEM_stage_inst_dmem_n2592) );
NAND2_X1 MEM_stage_inst_dmem_U2758 ( .A1(MEM_stage_inst_dmem_n2590), .A2(MEM_stage_inst_dmem_n2589), .ZN(MEM_stage_inst_dmem_n2594) );
NAND2_X1 MEM_stage_inst_dmem_U2757 ( .A1(MEM_stage_inst_dmem_ram_1780), .A2(MEM_stage_inst_dmem_n3202), .ZN(MEM_stage_inst_dmem_n2589) );
NAND2_X1 MEM_stage_inst_dmem_U2756 ( .A1(MEM_stage_inst_dmem_ram_1652), .A2(MEM_stage_inst_dmem_n4652), .ZN(MEM_stage_inst_dmem_n2590) );
NOR2_X1 MEM_stage_inst_dmem_U2755 ( .A1(MEM_stage_inst_dmem_n2588), .A2(MEM_stage_inst_dmem_n2587), .ZN(MEM_stage_inst_dmem_n2620) );
NAND2_X1 MEM_stage_inst_dmem_U2754 ( .A1(MEM_stage_inst_dmem_n2586), .A2(MEM_stage_inst_dmem_n2585), .ZN(MEM_stage_inst_dmem_n2587) );
NOR2_X1 MEM_stage_inst_dmem_U2753 ( .A1(MEM_stage_inst_dmem_n2584), .A2(MEM_stage_inst_dmem_n2583), .ZN(MEM_stage_inst_dmem_n2585) );
NAND2_X1 MEM_stage_inst_dmem_U2752 ( .A1(MEM_stage_inst_dmem_n2582), .A2(MEM_stage_inst_dmem_n2581), .ZN(MEM_stage_inst_dmem_n2583) );
NAND2_X1 MEM_stage_inst_dmem_U2751 ( .A1(MEM_stage_inst_dmem_ram_1412), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n2581) );
NAND2_X1 MEM_stage_inst_dmem_U2750 ( .A1(MEM_stage_inst_dmem_ram_1188), .A2(MEM_stage_inst_dmem_n3081), .ZN(MEM_stage_inst_dmem_n2582) );
NAND2_X1 MEM_stage_inst_dmem_U2749 ( .A1(MEM_stage_inst_dmem_n2580), .A2(MEM_stage_inst_dmem_n2579), .ZN(MEM_stage_inst_dmem_n2584) );
NAND2_X1 MEM_stage_inst_dmem_U2748 ( .A1(MEM_stage_inst_dmem_ram_1476), .A2(MEM_stage_inst_dmem_n3173), .ZN(MEM_stage_inst_dmem_n2579) );
NAND2_X1 MEM_stage_inst_dmem_U2747 ( .A1(MEM_stage_inst_dmem_ram_1172), .A2(MEM_stage_inst_dmem_n44), .ZN(MEM_stage_inst_dmem_n2580) );
NOR2_X1 MEM_stage_inst_dmem_U2746 ( .A1(MEM_stage_inst_dmem_n2578), .A2(MEM_stage_inst_dmem_n2577), .ZN(MEM_stage_inst_dmem_n2586) );
NAND2_X1 MEM_stage_inst_dmem_U2745 ( .A1(MEM_stage_inst_dmem_n2576), .A2(MEM_stage_inst_dmem_n2575), .ZN(MEM_stage_inst_dmem_n2577) );
NAND2_X1 MEM_stage_inst_dmem_U2744 ( .A1(MEM_stage_inst_dmem_ram_1988), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n2575) );
NAND2_X1 MEM_stage_inst_dmem_U2743 ( .A1(MEM_stage_inst_dmem_ram_1684), .A2(MEM_stage_inst_dmem_n3076), .ZN(MEM_stage_inst_dmem_n2576) );
NAND2_X1 MEM_stage_inst_dmem_U2742 ( .A1(MEM_stage_inst_dmem_n2574), .A2(MEM_stage_inst_dmem_n2573), .ZN(MEM_stage_inst_dmem_n2578) );
NAND2_X1 MEM_stage_inst_dmem_U2741 ( .A1(MEM_stage_inst_dmem_ram_1108), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n2573) );
NAND2_X1 MEM_stage_inst_dmem_U2740 ( .A1(MEM_stage_inst_dmem_ram_1604), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n2574) );
NAND2_X1 MEM_stage_inst_dmem_U2739 ( .A1(MEM_stage_inst_dmem_n2572), .A2(MEM_stage_inst_dmem_n2571), .ZN(MEM_stage_inst_dmem_n2588) );
NOR2_X1 MEM_stage_inst_dmem_U2738 ( .A1(MEM_stage_inst_dmem_n2570), .A2(MEM_stage_inst_dmem_n2569), .ZN(MEM_stage_inst_dmem_n2571) );
NAND2_X1 MEM_stage_inst_dmem_U2737 ( .A1(MEM_stage_inst_dmem_n2568), .A2(MEM_stage_inst_dmem_n2567), .ZN(MEM_stage_inst_dmem_n2569) );
NAND2_X1 MEM_stage_inst_dmem_U2736 ( .A1(MEM_stage_inst_dmem_ram_1508), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n2567) );
NAND2_X1 MEM_stage_inst_dmem_U2735 ( .A1(MEM_stage_inst_dmem_ram_1268), .A2(MEM_stage_inst_dmem_n39), .ZN(MEM_stage_inst_dmem_n2568) );
NAND2_X1 MEM_stage_inst_dmem_U2734 ( .A1(MEM_stage_inst_dmem_n2566), .A2(MEM_stage_inst_dmem_n2565), .ZN(MEM_stage_inst_dmem_n2570) );
NAND2_X1 MEM_stage_inst_dmem_U2733 ( .A1(MEM_stage_inst_dmem_ram_1492), .A2(MEM_stage_inst_dmem_n3174), .ZN(MEM_stage_inst_dmem_n2565) );
NAND2_X1 MEM_stage_inst_dmem_U2732 ( .A1(MEM_stage_inst_dmem_ram_1284), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n2566) );
NOR2_X1 MEM_stage_inst_dmem_U2731 ( .A1(MEM_stage_inst_dmem_n2564), .A2(MEM_stage_inst_dmem_n2563), .ZN(MEM_stage_inst_dmem_n2572) );
NAND2_X1 MEM_stage_inst_dmem_U2730 ( .A1(MEM_stage_inst_dmem_n2562), .A2(MEM_stage_inst_dmem_n2561), .ZN(MEM_stage_inst_dmem_n2563) );
NAND2_X1 MEM_stage_inst_dmem_U2729 ( .A1(MEM_stage_inst_dmem_ram_1252), .A2(MEM_stage_inst_dmem_n3152), .ZN(MEM_stage_inst_dmem_n2561) );
NAND2_X1 MEM_stage_inst_dmem_U2728 ( .A1(MEM_stage_inst_dmem_ram_1700), .A2(MEM_stage_inst_dmem_n3155), .ZN(MEM_stage_inst_dmem_n2562) );
NAND2_X1 MEM_stage_inst_dmem_U2727 ( .A1(MEM_stage_inst_dmem_n2560), .A2(MEM_stage_inst_dmem_n2559), .ZN(MEM_stage_inst_dmem_n2564) );
NAND2_X1 MEM_stage_inst_dmem_U2726 ( .A1(MEM_stage_inst_dmem_ram_1556), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n2559) );
NAND2_X1 MEM_stage_inst_dmem_U2725 ( .A1(MEM_stage_inst_dmem_ram_1124), .A2(MEM_stage_inst_dmem_n3179), .ZN(MEM_stage_inst_dmem_n2560) );
NOR2_X1 MEM_stage_inst_dmem_U2724 ( .A1(MEM_stage_inst_dmem_n2558), .A2(MEM_stage_inst_dmem_n2557), .ZN(MEM_stage_inst_dmem_n2816) );
NOR2_X1 MEM_stage_inst_dmem_U2723 ( .A1(MEM_stage_inst_dmem_n2556), .A2(MEM_stage_inst_dmem_n8286), .ZN(MEM_stage_inst_dmem_n2557) );
NOR2_X1 MEM_stage_inst_dmem_U2722 ( .A1(MEM_stage_inst_dmem_n2555), .A2(MEM_stage_inst_dmem_n2554), .ZN(MEM_stage_inst_dmem_n2556) );
NAND2_X1 MEM_stage_inst_dmem_U2721 ( .A1(MEM_stage_inst_dmem_n2553), .A2(MEM_stage_inst_dmem_n2552), .ZN(MEM_stage_inst_dmem_n2554) );
NOR2_X1 MEM_stage_inst_dmem_U2720 ( .A1(MEM_stage_inst_dmem_n2551), .A2(MEM_stage_inst_dmem_n2550), .ZN(MEM_stage_inst_dmem_n2552) );
NAND2_X1 MEM_stage_inst_dmem_U2719 ( .A1(MEM_stage_inst_dmem_n2549), .A2(MEM_stage_inst_dmem_n2548), .ZN(MEM_stage_inst_dmem_n2550) );
NOR2_X1 MEM_stage_inst_dmem_U2718 ( .A1(MEM_stage_inst_dmem_n2547), .A2(MEM_stage_inst_dmem_n2546), .ZN(MEM_stage_inst_dmem_n2548) );
NAND2_X1 MEM_stage_inst_dmem_U2717 ( .A1(MEM_stage_inst_dmem_n2545), .A2(MEM_stage_inst_dmem_n2544), .ZN(MEM_stage_inst_dmem_n2546) );
NAND2_X1 MEM_stage_inst_dmem_U2716 ( .A1(MEM_stage_inst_dmem_ram_2660), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n2544) );
NAND2_X1 MEM_stage_inst_dmem_U2715 ( .A1(MEM_stage_inst_dmem_ram_2388), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n2545) );
NAND2_X1 MEM_stage_inst_dmem_U2714 ( .A1(MEM_stage_inst_dmem_n2543), .A2(MEM_stage_inst_dmem_n2542), .ZN(MEM_stage_inst_dmem_n2547) );
NAND2_X1 MEM_stage_inst_dmem_U2713 ( .A1(MEM_stage_inst_dmem_ram_2452), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n2542) );
NAND2_X1 MEM_stage_inst_dmem_U2712 ( .A1(MEM_stage_inst_dmem_ram_2436), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n2543) );
NOR2_X1 MEM_stage_inst_dmem_U2711 ( .A1(MEM_stage_inst_dmem_n2541), .A2(MEM_stage_inst_dmem_n2540), .ZN(MEM_stage_inst_dmem_n2549) );
NAND2_X1 MEM_stage_inst_dmem_U2710 ( .A1(MEM_stage_inst_dmem_n2539), .A2(MEM_stage_inst_dmem_n2538), .ZN(MEM_stage_inst_dmem_n2540) );
NAND2_X1 MEM_stage_inst_dmem_U2709 ( .A1(MEM_stage_inst_dmem_ram_2052), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n2538) );
NAND2_X1 MEM_stage_inst_dmem_U2708 ( .A1(MEM_stage_inst_dmem_ram_2708), .A2(MEM_stage_inst_dmem_n3076), .ZN(MEM_stage_inst_dmem_n2539) );
NAND2_X1 MEM_stage_inst_dmem_U2707 ( .A1(MEM_stage_inst_dmem_n2537), .A2(MEM_stage_inst_dmem_n2536), .ZN(MEM_stage_inst_dmem_n2541) );
NAND2_X1 MEM_stage_inst_dmem_U2706 ( .A1(MEM_stage_inst_dmem_ram_2164), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n2536) );
NAND2_X1 MEM_stage_inst_dmem_U2705 ( .A1(MEM_stage_inst_dmem_ram_2228), .A2(MEM_stage_inst_dmem_n55), .ZN(MEM_stage_inst_dmem_n2537) );
NAND2_X1 MEM_stage_inst_dmem_U2704 ( .A1(MEM_stage_inst_dmem_n2535), .A2(MEM_stage_inst_dmem_n2534), .ZN(MEM_stage_inst_dmem_n2551) );
NOR2_X1 MEM_stage_inst_dmem_U2703 ( .A1(MEM_stage_inst_dmem_n2533), .A2(MEM_stage_inst_dmem_n2532), .ZN(MEM_stage_inst_dmem_n2534) );
NAND2_X1 MEM_stage_inst_dmem_U2702 ( .A1(MEM_stage_inst_dmem_n2531), .A2(MEM_stage_inst_dmem_n2530), .ZN(MEM_stage_inst_dmem_n2532) );
NAND2_X1 MEM_stage_inst_dmem_U2701 ( .A1(MEM_stage_inst_dmem_ram_2468), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n2530) );
NAND2_X1 MEM_stage_inst_dmem_U2700 ( .A1(MEM_stage_inst_dmem_ram_3060), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n2531) );
NAND2_X1 MEM_stage_inst_dmem_U2699 ( .A1(MEM_stage_inst_dmem_n2529), .A2(MEM_stage_inst_dmem_n2528), .ZN(MEM_stage_inst_dmem_n2533) );
NAND2_X1 MEM_stage_inst_dmem_U2698 ( .A1(MEM_stage_inst_dmem_ram_2372), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n2528) );
NAND2_X1 MEM_stage_inst_dmem_U2697 ( .A1(MEM_stage_inst_dmem_ram_2068), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n2529) );
NOR2_X1 MEM_stage_inst_dmem_U2696 ( .A1(MEM_stage_inst_dmem_n2527), .A2(MEM_stage_inst_dmem_n2526), .ZN(MEM_stage_inst_dmem_n2535) );
NAND2_X1 MEM_stage_inst_dmem_U2695 ( .A1(MEM_stage_inst_dmem_n2525), .A2(MEM_stage_inst_dmem_n2524), .ZN(MEM_stage_inst_dmem_n2526) );
NAND2_X1 MEM_stage_inst_dmem_U2694 ( .A1(MEM_stage_inst_dmem_ram_2484), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n2524) );
NAND2_X1 MEM_stage_inst_dmem_U2693 ( .A1(MEM_stage_inst_dmem_ram_2676), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n2525) );
NAND2_X1 MEM_stage_inst_dmem_U2692 ( .A1(MEM_stage_inst_dmem_n2523), .A2(MEM_stage_inst_dmem_n2522), .ZN(MEM_stage_inst_dmem_n2527) );
NAND2_X1 MEM_stage_inst_dmem_U2691 ( .A1(MEM_stage_inst_dmem_ram_2916), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n2522) );
NAND2_X1 MEM_stage_inst_dmem_U2690 ( .A1(MEM_stage_inst_dmem_ram_2340), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n2523) );
NOR2_X1 MEM_stage_inst_dmem_U2689 ( .A1(MEM_stage_inst_dmem_n2521), .A2(MEM_stage_inst_dmem_n2520), .ZN(MEM_stage_inst_dmem_n2553) );
NAND2_X1 MEM_stage_inst_dmem_U2688 ( .A1(MEM_stage_inst_dmem_n2519), .A2(MEM_stage_inst_dmem_n2518), .ZN(MEM_stage_inst_dmem_n2520) );
NOR2_X1 MEM_stage_inst_dmem_U2687 ( .A1(MEM_stage_inst_dmem_n2517), .A2(MEM_stage_inst_dmem_n2516), .ZN(MEM_stage_inst_dmem_n2518) );
NAND2_X1 MEM_stage_inst_dmem_U2686 ( .A1(MEM_stage_inst_dmem_n2515), .A2(MEM_stage_inst_dmem_n2514), .ZN(MEM_stage_inst_dmem_n2516) );
NAND2_X1 MEM_stage_inst_dmem_U2685 ( .A1(MEM_stage_inst_dmem_ram_2820), .A2(MEM_stage_inst_dmem_n37), .ZN(MEM_stage_inst_dmem_n2514) );
NAND2_X1 MEM_stage_inst_dmem_U2684 ( .A1(MEM_stage_inst_dmem_ram_2772), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n2515) );
NAND2_X1 MEM_stage_inst_dmem_U2683 ( .A1(MEM_stage_inst_dmem_n2513), .A2(MEM_stage_inst_dmem_n2512), .ZN(MEM_stage_inst_dmem_n2517) );
NAND2_X1 MEM_stage_inst_dmem_U2682 ( .A1(MEM_stage_inst_dmem_ram_2964), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n2512) );
NAND2_X1 MEM_stage_inst_dmem_U2681 ( .A1(MEM_stage_inst_dmem_ram_2260), .A2(MEM_stage_inst_dmem_n51), .ZN(MEM_stage_inst_dmem_n2513) );
NOR2_X1 MEM_stage_inst_dmem_U2680 ( .A1(MEM_stage_inst_dmem_n2511), .A2(MEM_stage_inst_dmem_n2510), .ZN(MEM_stage_inst_dmem_n2519) );
NAND2_X1 MEM_stage_inst_dmem_U2679 ( .A1(MEM_stage_inst_dmem_n2509), .A2(MEM_stage_inst_dmem_n2508), .ZN(MEM_stage_inst_dmem_n2510) );
NAND2_X1 MEM_stage_inst_dmem_U2678 ( .A1(MEM_stage_inst_dmem_ram_2244), .A2(MEM_stage_inst_dmem_n36), .ZN(MEM_stage_inst_dmem_n2508) );
NAND2_X1 MEM_stage_inst_dmem_U2677 ( .A1(MEM_stage_inst_dmem_ram_2788), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n2509) );
NAND2_X1 MEM_stage_inst_dmem_U2676 ( .A1(MEM_stage_inst_dmem_n2507), .A2(MEM_stage_inst_dmem_n2506), .ZN(MEM_stage_inst_dmem_n2511) );
NAND2_X1 MEM_stage_inst_dmem_U2675 ( .A1(MEM_stage_inst_dmem_ram_2948), .A2(MEM_stage_inst_dmem_n72), .ZN(MEM_stage_inst_dmem_n2506) );
NAND2_X1 MEM_stage_inst_dmem_U2674 ( .A1(MEM_stage_inst_dmem_ram_2324), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n2507) );
NAND2_X1 MEM_stage_inst_dmem_U2673 ( .A1(MEM_stage_inst_dmem_n2505), .A2(MEM_stage_inst_dmem_n2504), .ZN(MEM_stage_inst_dmem_n2521) );
NOR2_X1 MEM_stage_inst_dmem_U2672 ( .A1(MEM_stage_inst_dmem_n2503), .A2(MEM_stage_inst_dmem_n2502), .ZN(MEM_stage_inst_dmem_n2504) );
NAND2_X1 MEM_stage_inst_dmem_U2671 ( .A1(MEM_stage_inst_dmem_n2501), .A2(MEM_stage_inst_dmem_n2500), .ZN(MEM_stage_inst_dmem_n2502) );
NAND2_X1 MEM_stage_inst_dmem_U2670 ( .A1(MEM_stage_inst_dmem_ram_2356), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n2500) );
NAND2_X1 MEM_stage_inst_dmem_U2669 ( .A1(MEM_stage_inst_dmem_ram_2308), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n2501) );
NAND2_X1 MEM_stage_inst_dmem_U2668 ( .A1(MEM_stage_inst_dmem_n2499), .A2(MEM_stage_inst_dmem_n2498), .ZN(MEM_stage_inst_dmem_n2503) );
NAND2_X1 MEM_stage_inst_dmem_U2667 ( .A1(MEM_stage_inst_dmem_ram_2996), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n2498) );
NAND2_X1 MEM_stage_inst_dmem_U2666 ( .A1(MEM_stage_inst_dmem_ram_2116), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n2499) );
NOR2_X1 MEM_stage_inst_dmem_U2665 ( .A1(MEM_stage_inst_dmem_n2497), .A2(MEM_stage_inst_dmem_n2496), .ZN(MEM_stage_inst_dmem_n2505) );
NAND2_X1 MEM_stage_inst_dmem_U2664 ( .A1(MEM_stage_inst_dmem_n2495), .A2(MEM_stage_inst_dmem_n2494), .ZN(MEM_stage_inst_dmem_n2496) );
NAND2_X1 MEM_stage_inst_dmem_U2663 ( .A1(MEM_stage_inst_dmem_ram_3012), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n2494) );
NAND2_X1 MEM_stage_inst_dmem_U2662 ( .A1(MEM_stage_inst_dmem_ram_2516), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n2495) );
NAND2_X1 MEM_stage_inst_dmem_U2661 ( .A1(MEM_stage_inst_dmem_n2493), .A2(MEM_stage_inst_dmem_n2492), .ZN(MEM_stage_inst_dmem_n2497) );
NAND2_X1 MEM_stage_inst_dmem_U2660 ( .A1(MEM_stage_inst_dmem_ram_3044), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n2492) );
NAND2_X1 MEM_stage_inst_dmem_U2659 ( .A1(MEM_stage_inst_dmem_ram_2596), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n2493) );
NAND2_X1 MEM_stage_inst_dmem_U2658 ( .A1(MEM_stage_inst_dmem_n2491), .A2(MEM_stage_inst_dmem_n2490), .ZN(MEM_stage_inst_dmem_n2555) );
NOR2_X1 MEM_stage_inst_dmem_U2657 ( .A1(MEM_stage_inst_dmem_n2489), .A2(MEM_stage_inst_dmem_n2488), .ZN(MEM_stage_inst_dmem_n2490) );
NAND2_X1 MEM_stage_inst_dmem_U2656 ( .A1(MEM_stage_inst_dmem_n2487), .A2(MEM_stage_inst_dmem_n2486), .ZN(MEM_stage_inst_dmem_n2488) );
NOR2_X1 MEM_stage_inst_dmem_U2655 ( .A1(MEM_stage_inst_dmem_n2485), .A2(MEM_stage_inst_dmem_n2484), .ZN(MEM_stage_inst_dmem_n2486) );
NAND2_X1 MEM_stage_inst_dmem_U2654 ( .A1(MEM_stage_inst_dmem_n2483), .A2(MEM_stage_inst_dmem_n2482), .ZN(MEM_stage_inst_dmem_n2484) );
NAND2_X1 MEM_stage_inst_dmem_U2653 ( .A1(MEM_stage_inst_dmem_ram_2532), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n2482) );
NAND2_X1 MEM_stage_inst_dmem_U2652 ( .A1(MEM_stage_inst_dmem_ram_2500), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n2483) );
NAND2_X1 MEM_stage_inst_dmem_U2651 ( .A1(MEM_stage_inst_dmem_n2481), .A2(MEM_stage_inst_dmem_n2480), .ZN(MEM_stage_inst_dmem_n2485) );
NAND2_X1 MEM_stage_inst_dmem_U2650 ( .A1(MEM_stage_inst_dmem_ram_2276), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n2480) );
NAND2_X1 MEM_stage_inst_dmem_U2649 ( .A1(MEM_stage_inst_dmem_ram_2180), .A2(MEM_stage_inst_dmem_n61), .ZN(MEM_stage_inst_dmem_n2481) );
NOR2_X1 MEM_stage_inst_dmem_U2648 ( .A1(MEM_stage_inst_dmem_n2479), .A2(MEM_stage_inst_dmem_n2478), .ZN(MEM_stage_inst_dmem_n2487) );
NAND2_X1 MEM_stage_inst_dmem_U2647 ( .A1(MEM_stage_inst_dmem_n2477), .A2(MEM_stage_inst_dmem_n2476), .ZN(MEM_stage_inst_dmem_n2478) );
NAND2_X1 MEM_stage_inst_dmem_U2646 ( .A1(MEM_stage_inst_dmem_ram_2692), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n2476) );
NAND2_X1 MEM_stage_inst_dmem_U2645 ( .A1(MEM_stage_inst_dmem_ram_2580), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n2477) );
NAND2_X1 MEM_stage_inst_dmem_U2644 ( .A1(MEM_stage_inst_dmem_n2475), .A2(MEM_stage_inst_dmem_n2474), .ZN(MEM_stage_inst_dmem_n2479) );
NAND2_X1 MEM_stage_inst_dmem_U2643 ( .A1(MEM_stage_inst_dmem_ram_2884), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n2474) );
NAND2_X1 MEM_stage_inst_dmem_U2642 ( .A1(MEM_stage_inst_dmem_ram_2868), .A2(MEM_stage_inst_dmem_n8005), .ZN(MEM_stage_inst_dmem_n2475) );
NAND2_X1 MEM_stage_inst_dmem_U2641 ( .A1(MEM_stage_inst_dmem_n2473), .A2(MEM_stage_inst_dmem_n2472), .ZN(MEM_stage_inst_dmem_n2489) );
NOR2_X1 MEM_stage_inst_dmem_U2640 ( .A1(MEM_stage_inst_dmem_n2471), .A2(MEM_stage_inst_dmem_n2470), .ZN(MEM_stage_inst_dmem_n2472) );
NAND2_X1 MEM_stage_inst_dmem_U2639 ( .A1(MEM_stage_inst_dmem_n2469), .A2(MEM_stage_inst_dmem_n2468), .ZN(MEM_stage_inst_dmem_n2470) );
NAND2_X1 MEM_stage_inst_dmem_U2638 ( .A1(MEM_stage_inst_dmem_ram_2292), .A2(MEM_stage_inst_dmem_n7914), .ZN(MEM_stage_inst_dmem_n2468) );
NAND2_X1 MEM_stage_inst_dmem_U2637 ( .A1(MEM_stage_inst_dmem_ram_2212), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n2469) );
NAND2_X1 MEM_stage_inst_dmem_U2636 ( .A1(MEM_stage_inst_dmem_n2467), .A2(MEM_stage_inst_dmem_n2466), .ZN(MEM_stage_inst_dmem_n2471) );
NAND2_X1 MEM_stage_inst_dmem_U2635 ( .A1(MEM_stage_inst_dmem_ram_2980), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n2466) );
NAND2_X1 MEM_stage_inst_dmem_U2634 ( .A1(MEM_stage_inst_dmem_ram_2420), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n2467) );
NOR2_X1 MEM_stage_inst_dmem_U2633 ( .A1(MEM_stage_inst_dmem_n2465), .A2(MEM_stage_inst_dmem_n2464), .ZN(MEM_stage_inst_dmem_n2473) );
NAND2_X1 MEM_stage_inst_dmem_U2632 ( .A1(MEM_stage_inst_dmem_n2463), .A2(MEM_stage_inst_dmem_n2462), .ZN(MEM_stage_inst_dmem_n2464) );
NAND2_X1 MEM_stage_inst_dmem_U2631 ( .A1(MEM_stage_inst_dmem_ram_2852), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n2462) );
NAND2_X1 MEM_stage_inst_dmem_U2630 ( .A1(MEM_stage_inst_dmem_ram_2740), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n2463) );
NAND2_X1 MEM_stage_inst_dmem_U2629 ( .A1(MEM_stage_inst_dmem_n2461), .A2(MEM_stage_inst_dmem_n2460), .ZN(MEM_stage_inst_dmem_n2465) );
NAND2_X1 MEM_stage_inst_dmem_U2628 ( .A1(MEM_stage_inst_dmem_ram_2612), .A2(MEM_stage_inst_dmem_n41), .ZN(MEM_stage_inst_dmem_n2460) );
NAND2_X1 MEM_stage_inst_dmem_U2627 ( .A1(MEM_stage_inst_dmem_ram_2132), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n2461) );
NOR2_X1 MEM_stage_inst_dmem_U2626 ( .A1(MEM_stage_inst_dmem_n2459), .A2(MEM_stage_inst_dmem_n2458), .ZN(MEM_stage_inst_dmem_n2491) );
NAND2_X1 MEM_stage_inst_dmem_U2625 ( .A1(MEM_stage_inst_dmem_n2457), .A2(MEM_stage_inst_dmem_n2456), .ZN(MEM_stage_inst_dmem_n2458) );
NOR2_X1 MEM_stage_inst_dmem_U2624 ( .A1(MEM_stage_inst_dmem_n2455), .A2(MEM_stage_inst_dmem_n2454), .ZN(MEM_stage_inst_dmem_n2456) );
NAND2_X1 MEM_stage_inst_dmem_U2623 ( .A1(MEM_stage_inst_dmem_n2453), .A2(MEM_stage_inst_dmem_n2452), .ZN(MEM_stage_inst_dmem_n2454) );
NAND2_X1 MEM_stage_inst_dmem_U2622 ( .A1(MEM_stage_inst_dmem_ram_2100), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n2452) );
NAND2_X1 MEM_stage_inst_dmem_U2621 ( .A1(MEM_stage_inst_dmem_ram_2084), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n2453) );
NAND2_X1 MEM_stage_inst_dmem_U2620 ( .A1(MEM_stage_inst_dmem_n2451), .A2(MEM_stage_inst_dmem_n2450), .ZN(MEM_stage_inst_dmem_n2455) );
NAND2_X1 MEM_stage_inst_dmem_U2619 ( .A1(MEM_stage_inst_dmem_ram_2804), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n2450) );
NAND2_X1 MEM_stage_inst_dmem_U2618 ( .A1(MEM_stage_inst_dmem_ram_2836), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n2451) );
NOR2_X1 MEM_stage_inst_dmem_U2617 ( .A1(MEM_stage_inst_dmem_n2449), .A2(MEM_stage_inst_dmem_n2448), .ZN(MEM_stage_inst_dmem_n2457) );
NAND2_X1 MEM_stage_inst_dmem_U2616 ( .A1(MEM_stage_inst_dmem_n2447), .A2(MEM_stage_inst_dmem_n2446), .ZN(MEM_stage_inst_dmem_n2448) );
NAND2_X1 MEM_stage_inst_dmem_U2615 ( .A1(MEM_stage_inst_dmem_ram_2932), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n2446) );
NAND2_X1 MEM_stage_inst_dmem_U2614 ( .A1(MEM_stage_inst_dmem_ram_2196), .A2(MEM_stage_inst_dmem_n44), .ZN(MEM_stage_inst_dmem_n2447) );
NAND2_X1 MEM_stage_inst_dmem_U2613 ( .A1(MEM_stage_inst_dmem_n2445), .A2(MEM_stage_inst_dmem_n2444), .ZN(MEM_stage_inst_dmem_n2449) );
NAND2_X1 MEM_stage_inst_dmem_U2612 ( .A1(MEM_stage_inst_dmem_ram_2148), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n2444) );
NAND2_X1 MEM_stage_inst_dmem_U2611 ( .A1(MEM_stage_inst_dmem_ram_2628), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n2445) );
NAND2_X1 MEM_stage_inst_dmem_U2610 ( .A1(MEM_stage_inst_dmem_n2443), .A2(MEM_stage_inst_dmem_n2442), .ZN(MEM_stage_inst_dmem_n2459) );
NOR2_X1 MEM_stage_inst_dmem_U2609 ( .A1(MEM_stage_inst_dmem_n2441), .A2(MEM_stage_inst_dmem_n2440), .ZN(MEM_stage_inst_dmem_n2442) );
NAND2_X1 MEM_stage_inst_dmem_U2608 ( .A1(MEM_stage_inst_dmem_n2439), .A2(MEM_stage_inst_dmem_n2438), .ZN(MEM_stage_inst_dmem_n2440) );
NAND2_X1 MEM_stage_inst_dmem_U2607 ( .A1(MEM_stage_inst_dmem_ram_2756), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n2438) );
NAND2_X1 MEM_stage_inst_dmem_U2606 ( .A1(MEM_stage_inst_dmem_ram_2644), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n2439) );
NAND2_X1 MEM_stage_inst_dmem_U2605 ( .A1(MEM_stage_inst_dmem_n2437), .A2(MEM_stage_inst_dmem_n2436), .ZN(MEM_stage_inst_dmem_n2441) );
NAND2_X1 MEM_stage_inst_dmem_U2604 ( .A1(MEM_stage_inst_dmem_ram_2548), .A2(MEM_stage_inst_dmem_n8535), .ZN(MEM_stage_inst_dmem_n2436) );
NAND2_X1 MEM_stage_inst_dmem_U2603 ( .A1(MEM_stage_inst_dmem_ram_3028), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n2437) );
NOR2_X1 MEM_stage_inst_dmem_U2602 ( .A1(MEM_stage_inst_dmem_n2435), .A2(MEM_stage_inst_dmem_n2434), .ZN(MEM_stage_inst_dmem_n2443) );
NAND2_X1 MEM_stage_inst_dmem_U2601 ( .A1(MEM_stage_inst_dmem_n2433), .A2(MEM_stage_inst_dmem_n2432), .ZN(MEM_stage_inst_dmem_n2434) );
NAND2_X1 MEM_stage_inst_dmem_U2600 ( .A1(MEM_stage_inst_dmem_ram_2900), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n2432) );
NAND2_X1 MEM_stage_inst_dmem_U2599 ( .A1(MEM_stage_inst_dmem_ram_2564), .A2(MEM_stage_inst_dmem_n71), .ZN(MEM_stage_inst_dmem_n2433) );
NAND2_X1 MEM_stage_inst_dmem_U2598 ( .A1(MEM_stage_inst_dmem_n2431), .A2(MEM_stage_inst_dmem_n2430), .ZN(MEM_stage_inst_dmem_n2435) );
NAND2_X1 MEM_stage_inst_dmem_U2597 ( .A1(MEM_stage_inst_dmem_ram_2404), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n2430) );
NAND2_X1 MEM_stage_inst_dmem_U2596 ( .A1(MEM_stage_inst_dmem_ram_2724), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n2431) );
NOR2_X1 MEM_stage_inst_dmem_U2595 ( .A1(MEM_stage_inst_dmem_n2429), .A2(MEM_stage_inst_dmem_n8551), .ZN(MEM_stage_inst_dmem_n2558) );
NOR2_X1 MEM_stage_inst_dmem_U2594 ( .A1(MEM_stage_inst_dmem_n2428), .A2(MEM_stage_inst_dmem_n2427), .ZN(MEM_stage_inst_dmem_n2429) );
NAND2_X1 MEM_stage_inst_dmem_U2593 ( .A1(MEM_stage_inst_dmem_n2426), .A2(MEM_stage_inst_dmem_n2425), .ZN(MEM_stage_inst_dmem_n2427) );
NOR2_X1 MEM_stage_inst_dmem_U2592 ( .A1(MEM_stage_inst_dmem_n2424), .A2(MEM_stage_inst_dmem_n2423), .ZN(MEM_stage_inst_dmem_n2425) );
NAND2_X1 MEM_stage_inst_dmem_U2591 ( .A1(MEM_stage_inst_dmem_n2422), .A2(MEM_stage_inst_dmem_n2421), .ZN(MEM_stage_inst_dmem_n2423) );
NOR2_X1 MEM_stage_inst_dmem_U2590 ( .A1(MEM_stage_inst_dmem_n2420), .A2(MEM_stage_inst_dmem_n2419), .ZN(MEM_stage_inst_dmem_n2421) );
NAND2_X1 MEM_stage_inst_dmem_U2589 ( .A1(MEM_stage_inst_dmem_n2418), .A2(MEM_stage_inst_dmem_n2417), .ZN(MEM_stage_inst_dmem_n2419) );
NAND2_X1 MEM_stage_inst_dmem_U2588 ( .A1(MEM_stage_inst_dmem_ram_484), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n2417) );
NAND2_X1 MEM_stage_inst_dmem_U2587 ( .A1(MEM_stage_inst_dmem_ram_516), .A2(MEM_stage_inst_dmem_n71), .ZN(MEM_stage_inst_dmem_n2418) );
NAND2_X1 MEM_stage_inst_dmem_U2586 ( .A1(MEM_stage_inst_dmem_n2416), .A2(MEM_stage_inst_dmem_n2415), .ZN(MEM_stage_inst_dmem_n2420) );
NAND2_X1 MEM_stage_inst_dmem_U2585 ( .A1(MEM_stage_inst_dmem_ram_916), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n2415) );
NAND2_X1 MEM_stage_inst_dmem_U2584 ( .A1(MEM_stage_inst_dmem_ram_580), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n2416) );
NOR2_X1 MEM_stage_inst_dmem_U2583 ( .A1(MEM_stage_inst_dmem_n2414), .A2(MEM_stage_inst_dmem_n2413), .ZN(MEM_stage_inst_dmem_n2422) );
NAND2_X1 MEM_stage_inst_dmem_U2582 ( .A1(MEM_stage_inst_dmem_n2412), .A2(MEM_stage_inst_dmem_n2411), .ZN(MEM_stage_inst_dmem_n2413) );
NAND2_X1 MEM_stage_inst_dmem_U2581 ( .A1(MEM_stage_inst_dmem_ram_388), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n2411) );
NAND2_X1 MEM_stage_inst_dmem_U2580 ( .A1(MEM_stage_inst_dmem_ram_724), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n2412) );
NAND2_X1 MEM_stage_inst_dmem_U2579 ( .A1(MEM_stage_inst_dmem_n2410), .A2(MEM_stage_inst_dmem_n2409), .ZN(MEM_stage_inst_dmem_n2414) );
NAND2_X1 MEM_stage_inst_dmem_U2578 ( .A1(MEM_stage_inst_dmem_ram_836), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n2409) );
NAND2_X1 MEM_stage_inst_dmem_U2577 ( .A1(MEM_stage_inst_dmem_ram_372), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n2410) );
NAND2_X1 MEM_stage_inst_dmem_U2576 ( .A1(MEM_stage_inst_dmem_n2408), .A2(MEM_stage_inst_dmem_n2407), .ZN(MEM_stage_inst_dmem_n2424) );
NOR2_X1 MEM_stage_inst_dmem_U2575 ( .A1(MEM_stage_inst_dmem_n2406), .A2(MEM_stage_inst_dmem_n2405), .ZN(MEM_stage_inst_dmem_n2407) );
NAND2_X1 MEM_stage_inst_dmem_U2574 ( .A1(MEM_stage_inst_dmem_n2404), .A2(MEM_stage_inst_dmem_n2403), .ZN(MEM_stage_inst_dmem_n2405) );
NAND2_X1 MEM_stage_inst_dmem_U2573 ( .A1(MEM_stage_inst_dmem_ram_36), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n2403) );
NAND2_X1 MEM_stage_inst_dmem_U2572 ( .A1(MEM_stage_inst_dmem_ram_596), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n2404) );
NAND2_X1 MEM_stage_inst_dmem_U2571 ( .A1(MEM_stage_inst_dmem_n2402), .A2(MEM_stage_inst_dmem_n2401), .ZN(MEM_stage_inst_dmem_n2406) );
NAND2_X1 MEM_stage_inst_dmem_U2570 ( .A1(MEM_stage_inst_dmem_ram_772), .A2(MEM_stage_inst_dmem_n37), .ZN(MEM_stage_inst_dmem_n2401) );
NAND2_X1 MEM_stage_inst_dmem_U2569 ( .A1(MEM_stage_inst_dmem_ram_452), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n2402) );
NOR2_X1 MEM_stage_inst_dmem_U2568 ( .A1(MEM_stage_inst_dmem_n2400), .A2(MEM_stage_inst_dmem_n2399), .ZN(MEM_stage_inst_dmem_n2408) );
NAND2_X1 MEM_stage_inst_dmem_U2567 ( .A1(MEM_stage_inst_dmem_n2398), .A2(MEM_stage_inst_dmem_n2397), .ZN(MEM_stage_inst_dmem_n2399) );
NAND2_X1 MEM_stage_inst_dmem_U2566 ( .A1(MEM_stage_inst_dmem_ram_852), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n2397) );
NAND2_X1 MEM_stage_inst_dmem_U2565 ( .A1(MEM_stage_inst_dmem_ram_948), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n2398) );
NAND2_X1 MEM_stage_inst_dmem_U2564 ( .A1(MEM_stage_inst_dmem_n2396), .A2(MEM_stage_inst_dmem_n2395), .ZN(MEM_stage_inst_dmem_n2400) );
NAND2_X1 MEM_stage_inst_dmem_U2563 ( .A1(MEM_stage_inst_dmem_ram_148), .A2(MEM_stage_inst_dmem_n44), .ZN(MEM_stage_inst_dmem_n2395) );
NAND2_X1 MEM_stage_inst_dmem_U2562 ( .A1(MEM_stage_inst_dmem_ram_740), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n2396) );
NOR2_X1 MEM_stage_inst_dmem_U2561 ( .A1(MEM_stage_inst_dmem_n2394), .A2(MEM_stage_inst_dmem_n2393), .ZN(MEM_stage_inst_dmem_n2426) );
NAND2_X1 MEM_stage_inst_dmem_U2560 ( .A1(MEM_stage_inst_dmem_n2392), .A2(MEM_stage_inst_dmem_n2391), .ZN(MEM_stage_inst_dmem_n2393) );
NOR2_X1 MEM_stage_inst_dmem_U2559 ( .A1(MEM_stage_inst_dmem_n2390), .A2(MEM_stage_inst_dmem_n2389), .ZN(MEM_stage_inst_dmem_n2391) );
NAND2_X1 MEM_stage_inst_dmem_U2558 ( .A1(MEM_stage_inst_dmem_n2388), .A2(MEM_stage_inst_dmem_n2387), .ZN(MEM_stage_inst_dmem_n2389) );
NAND2_X1 MEM_stage_inst_dmem_U2557 ( .A1(MEM_stage_inst_dmem_ram_980), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n2387) );
NAND2_X1 MEM_stage_inst_dmem_U2556 ( .A1(MEM_stage_inst_dmem_ram_468), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n2388) );
NAND2_X1 MEM_stage_inst_dmem_U2555 ( .A1(MEM_stage_inst_dmem_n2386), .A2(MEM_stage_inst_dmem_n2385), .ZN(MEM_stage_inst_dmem_n2390) );
NAND2_X1 MEM_stage_inst_dmem_U2554 ( .A1(MEM_stage_inst_dmem_ram_884), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n2385) );
NAND2_X1 MEM_stage_inst_dmem_U2553 ( .A1(MEM_stage_inst_dmem_ram_420), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n2386) );
NOR2_X1 MEM_stage_inst_dmem_U2552 ( .A1(MEM_stage_inst_dmem_n2384), .A2(MEM_stage_inst_dmem_n2383), .ZN(MEM_stage_inst_dmem_n2392) );
NAND2_X1 MEM_stage_inst_dmem_U2551 ( .A1(MEM_stage_inst_dmem_n2382), .A2(MEM_stage_inst_dmem_n2381), .ZN(MEM_stage_inst_dmem_n2383) );
NAND2_X1 MEM_stage_inst_dmem_U2550 ( .A1(MEM_stage_inst_dmem_ram_996), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n2381) );
NAND2_X1 MEM_stage_inst_dmem_U2549 ( .A1(MEM_stage_inst_dmem_ram_212), .A2(MEM_stage_inst_dmem_n51), .ZN(MEM_stage_inst_dmem_n2382) );
NAND2_X1 MEM_stage_inst_dmem_U2548 ( .A1(MEM_stage_inst_dmem_n2380), .A2(MEM_stage_inst_dmem_n2379), .ZN(MEM_stage_inst_dmem_n2384) );
NAND2_X1 MEM_stage_inst_dmem_U2547 ( .A1(MEM_stage_inst_dmem_ram_324), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n2379) );
NAND2_X1 MEM_stage_inst_dmem_U2546 ( .A1(MEM_stage_inst_dmem_ram_292), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n2380) );
NAND2_X1 MEM_stage_inst_dmem_U2545 ( .A1(MEM_stage_inst_dmem_n2378), .A2(MEM_stage_inst_dmem_n2377), .ZN(MEM_stage_inst_dmem_n2394) );
NOR2_X1 MEM_stage_inst_dmem_U2544 ( .A1(MEM_stage_inst_dmem_n2376), .A2(MEM_stage_inst_dmem_n2375), .ZN(MEM_stage_inst_dmem_n2377) );
NAND2_X1 MEM_stage_inst_dmem_U2543 ( .A1(MEM_stage_inst_dmem_n2374), .A2(MEM_stage_inst_dmem_n2373), .ZN(MEM_stage_inst_dmem_n2375) );
NAND2_X1 MEM_stage_inst_dmem_U2542 ( .A1(MEM_stage_inst_dmem_ram_548), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n2373) );
NAND2_X1 MEM_stage_inst_dmem_U2541 ( .A1(MEM_stage_inst_dmem_ram_788), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n2374) );
NAND2_X1 MEM_stage_inst_dmem_U2540 ( .A1(MEM_stage_inst_dmem_n2372), .A2(MEM_stage_inst_dmem_n2371), .ZN(MEM_stage_inst_dmem_n2376) );
NAND2_X1 MEM_stage_inst_dmem_U2539 ( .A1(MEM_stage_inst_dmem_ram_68), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n2371) );
NAND2_X1 MEM_stage_inst_dmem_U2538 ( .A1(MEM_stage_inst_dmem_ram_756), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n2372) );
NOR2_X1 MEM_stage_inst_dmem_U2537 ( .A1(MEM_stage_inst_dmem_n2370), .A2(MEM_stage_inst_dmem_n2369), .ZN(MEM_stage_inst_dmem_n2378) );
NAND2_X1 MEM_stage_inst_dmem_U2536 ( .A1(MEM_stage_inst_dmem_n2368), .A2(MEM_stage_inst_dmem_n2367), .ZN(MEM_stage_inst_dmem_n2369) );
NAND2_X1 MEM_stage_inst_dmem_U2535 ( .A1(MEM_stage_inst_dmem_ram_868), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n2367) );
NAND2_X1 MEM_stage_inst_dmem_U2534 ( .A1(MEM_stage_inst_dmem_ram_804), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n2368) );
NAND2_X1 MEM_stage_inst_dmem_U2533 ( .A1(MEM_stage_inst_dmem_n2366), .A2(MEM_stage_inst_dmem_n2365), .ZN(MEM_stage_inst_dmem_n2370) );
NAND2_X1 MEM_stage_inst_dmem_U2532 ( .A1(MEM_stage_inst_dmem_ram_356), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n2365) );
NAND2_X1 MEM_stage_inst_dmem_U2531 ( .A1(MEM_stage_inst_dmem_ram_612), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n2366) );
NAND2_X1 MEM_stage_inst_dmem_U2530 ( .A1(MEM_stage_inst_dmem_n2364), .A2(MEM_stage_inst_dmem_n2363), .ZN(MEM_stage_inst_dmem_n2428) );
NOR2_X1 MEM_stage_inst_dmem_U2529 ( .A1(MEM_stage_inst_dmem_n2362), .A2(MEM_stage_inst_dmem_n2361), .ZN(MEM_stage_inst_dmem_n2363) );
NAND2_X1 MEM_stage_inst_dmem_U2528 ( .A1(MEM_stage_inst_dmem_n2360), .A2(MEM_stage_inst_dmem_n2359), .ZN(MEM_stage_inst_dmem_n2361) );
NOR2_X1 MEM_stage_inst_dmem_U2527 ( .A1(MEM_stage_inst_dmem_n2358), .A2(MEM_stage_inst_dmem_n2357), .ZN(MEM_stage_inst_dmem_n2359) );
NAND2_X1 MEM_stage_inst_dmem_U2526 ( .A1(MEM_stage_inst_dmem_n2356), .A2(MEM_stage_inst_dmem_n2355), .ZN(MEM_stage_inst_dmem_n2357) );
NAND2_X1 MEM_stage_inst_dmem_U2525 ( .A1(MEM_stage_inst_dmem_ram_692), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n2355) );
NAND2_X1 MEM_stage_inst_dmem_U2524 ( .A1(MEM_stage_inst_dmem_ram_660), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n2356) );
NAND2_X1 MEM_stage_inst_dmem_U2523 ( .A1(MEM_stage_inst_dmem_n2354), .A2(MEM_stage_inst_dmem_n2353), .ZN(MEM_stage_inst_dmem_n2358) );
NAND2_X1 MEM_stage_inst_dmem_U2522 ( .A1(MEM_stage_inst_dmem_ram_180), .A2(MEM_stage_inst_dmem_n55), .ZN(MEM_stage_inst_dmem_n2353) );
NAND2_X1 MEM_stage_inst_dmem_U2521 ( .A1(MEM_stage_inst_dmem_ram_532), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n2354) );
NOR2_X1 MEM_stage_inst_dmem_U2520 ( .A1(MEM_stage_inst_dmem_n2352), .A2(MEM_stage_inst_dmem_n2351), .ZN(MEM_stage_inst_dmem_n2360) );
NAND2_X1 MEM_stage_inst_dmem_U2519 ( .A1(MEM_stage_inst_dmem_n2350), .A2(MEM_stage_inst_dmem_n2349), .ZN(MEM_stage_inst_dmem_n2351) );
NAND2_X1 MEM_stage_inst_dmem_U2518 ( .A1(MEM_stage_inst_dmem_ram_644), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n2349) );
NAND2_X1 MEM_stage_inst_dmem_U2517 ( .A1(MEM_stage_inst_dmem_ram_244), .A2(MEM_stage_inst_dmem_n39), .ZN(MEM_stage_inst_dmem_n2350) );
NAND2_X1 MEM_stage_inst_dmem_U2516 ( .A1(MEM_stage_inst_dmem_n2348), .A2(MEM_stage_inst_dmem_n2347), .ZN(MEM_stage_inst_dmem_n2352) );
NAND2_X1 MEM_stage_inst_dmem_U2515 ( .A1(MEM_stage_inst_dmem_ram_964), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n2347) );
NAND2_X1 MEM_stage_inst_dmem_U2514 ( .A1(MEM_stage_inst_dmem_ram_100), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n2348) );
NAND2_X1 MEM_stage_inst_dmem_U2513 ( .A1(MEM_stage_inst_dmem_n2346), .A2(MEM_stage_inst_dmem_n2345), .ZN(MEM_stage_inst_dmem_n2362) );
NOR2_X1 MEM_stage_inst_dmem_U2512 ( .A1(MEM_stage_inst_dmem_n2344), .A2(MEM_stage_inst_dmem_n2343), .ZN(MEM_stage_inst_dmem_n2345) );
NAND2_X1 MEM_stage_inst_dmem_U2511 ( .A1(MEM_stage_inst_dmem_n2342), .A2(MEM_stage_inst_dmem_n2341), .ZN(MEM_stage_inst_dmem_n2343) );
NAND2_X1 MEM_stage_inst_dmem_U2510 ( .A1(MEM_stage_inst_dmem_ram_132), .A2(MEM_stage_inst_dmem_n61), .ZN(MEM_stage_inst_dmem_n2341) );
NAND2_X1 MEM_stage_inst_dmem_U2509 ( .A1(MEM_stage_inst_dmem_ram_676), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n2342) );
NAND2_X1 MEM_stage_inst_dmem_U2508 ( .A1(MEM_stage_inst_dmem_n2340), .A2(MEM_stage_inst_dmem_n2339), .ZN(MEM_stage_inst_dmem_n2344) );
NAND2_X1 MEM_stage_inst_dmem_U2507 ( .A1(MEM_stage_inst_dmem_ram_84), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n2339) );
NAND2_X1 MEM_stage_inst_dmem_U2506 ( .A1(MEM_stage_inst_dmem_ram_932), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n2340) );
NOR2_X1 MEM_stage_inst_dmem_U2505 ( .A1(MEM_stage_inst_dmem_n2338), .A2(MEM_stage_inst_dmem_n2337), .ZN(MEM_stage_inst_dmem_n2346) );
NAND2_X1 MEM_stage_inst_dmem_U2504 ( .A1(MEM_stage_inst_dmem_n2336), .A2(MEM_stage_inst_dmem_n2335), .ZN(MEM_stage_inst_dmem_n2337) );
NAND2_X1 MEM_stage_inst_dmem_U2503 ( .A1(MEM_stage_inst_dmem_ram_52), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n2335) );
NAND2_X1 MEM_stage_inst_dmem_U2502 ( .A1(MEM_stage_inst_dmem_ram_164), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n2336) );
NAND2_X1 MEM_stage_inst_dmem_U2501 ( .A1(MEM_stage_inst_dmem_n2334), .A2(MEM_stage_inst_dmem_n2333), .ZN(MEM_stage_inst_dmem_n2338) );
NAND2_X1 MEM_stage_inst_dmem_U2500 ( .A1(MEM_stage_inst_dmem_ram_820), .A2(MEM_stage_inst_dmem_n46), .ZN(MEM_stage_inst_dmem_n2333) );
NAND2_X1 MEM_stage_inst_dmem_U2499 ( .A1(MEM_stage_inst_dmem_ram_260), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n2334) );
NOR2_X1 MEM_stage_inst_dmem_U2498 ( .A1(MEM_stage_inst_dmem_n2332), .A2(MEM_stage_inst_dmem_n2331), .ZN(MEM_stage_inst_dmem_n2364) );
NAND2_X1 MEM_stage_inst_dmem_U2497 ( .A1(MEM_stage_inst_dmem_n2330), .A2(MEM_stage_inst_dmem_n2329), .ZN(MEM_stage_inst_dmem_n2331) );
NOR2_X1 MEM_stage_inst_dmem_U2496 ( .A1(MEM_stage_inst_dmem_n2328), .A2(MEM_stage_inst_dmem_n2327), .ZN(MEM_stage_inst_dmem_n2329) );
NAND2_X1 MEM_stage_inst_dmem_U2495 ( .A1(MEM_stage_inst_dmem_n2326), .A2(MEM_stage_inst_dmem_n2325), .ZN(MEM_stage_inst_dmem_n2327) );
NAND2_X1 MEM_stage_inst_dmem_U2494 ( .A1(MEM_stage_inst_dmem_ram_196), .A2(MEM_stage_inst_dmem_n36), .ZN(MEM_stage_inst_dmem_n2325) );
NAND2_X1 MEM_stage_inst_dmem_U2493 ( .A1(MEM_stage_inst_dmem_ram_228), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n2326) );
NAND2_X1 MEM_stage_inst_dmem_U2492 ( .A1(MEM_stage_inst_dmem_n2324), .A2(MEM_stage_inst_dmem_n2323), .ZN(MEM_stage_inst_dmem_n2328) );
NAND2_X1 MEM_stage_inst_dmem_U2491 ( .A1(MEM_stage_inst_dmem_ram_708), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n2323) );
NAND2_X1 MEM_stage_inst_dmem_U2490 ( .A1(MEM_stage_inst_dmem_ram_900), .A2(MEM_stage_inst_dmem_n72), .ZN(MEM_stage_inst_dmem_n2324) );
NOR2_X1 MEM_stage_inst_dmem_U2489 ( .A1(MEM_stage_inst_dmem_n2322), .A2(MEM_stage_inst_dmem_n2321), .ZN(MEM_stage_inst_dmem_n2330) );
NAND2_X1 MEM_stage_inst_dmem_U2488 ( .A1(MEM_stage_inst_dmem_n2320), .A2(MEM_stage_inst_dmem_n2319), .ZN(MEM_stage_inst_dmem_n2321) );
NAND2_X1 MEM_stage_inst_dmem_U2487 ( .A1(MEM_stage_inst_dmem_ram_308), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n2319) );
NAND2_X1 MEM_stage_inst_dmem_U2486 ( .A1(MEM_stage_inst_dmem_ram_628), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n2320) );
NAND2_X1 MEM_stage_inst_dmem_U2485 ( .A1(MEM_stage_inst_dmem_n2318), .A2(MEM_stage_inst_dmem_n2317), .ZN(MEM_stage_inst_dmem_n2322) );
NAND2_X1 MEM_stage_inst_dmem_U2484 ( .A1(MEM_stage_inst_dmem_ram_564), .A2(MEM_stage_inst_dmem_n41), .ZN(MEM_stage_inst_dmem_n2317) );
NAND2_X1 MEM_stage_inst_dmem_U2483 ( .A1(MEM_stage_inst_dmem_ram_1012), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n2318) );
NAND2_X1 MEM_stage_inst_dmem_U2482 ( .A1(MEM_stage_inst_dmem_n2316), .A2(MEM_stage_inst_dmem_n2315), .ZN(MEM_stage_inst_dmem_n2332) );
NOR2_X1 MEM_stage_inst_dmem_U2481 ( .A1(MEM_stage_inst_dmem_n2314), .A2(MEM_stage_inst_dmem_n2313), .ZN(MEM_stage_inst_dmem_n2315) );
NAND2_X1 MEM_stage_inst_dmem_U2480 ( .A1(MEM_stage_inst_dmem_n2312), .A2(MEM_stage_inst_dmem_n2311), .ZN(MEM_stage_inst_dmem_n2313) );
NAND2_X1 MEM_stage_inst_dmem_U2479 ( .A1(MEM_stage_inst_dmem_ram_500), .A2(MEM_stage_inst_dmem_n8535), .ZN(MEM_stage_inst_dmem_n2311) );
NAND2_X1 MEM_stage_inst_dmem_U2478 ( .A1(MEM_stage_inst_dmem_ram_116), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n2312) );
NAND2_X1 MEM_stage_inst_dmem_U2477 ( .A1(MEM_stage_inst_dmem_n2310), .A2(MEM_stage_inst_dmem_n2309), .ZN(MEM_stage_inst_dmem_n2314) );
NAND2_X1 MEM_stage_inst_dmem_U2476 ( .A1(MEM_stage_inst_dmem_ram_436), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n2309) );
NAND2_X1 MEM_stage_inst_dmem_U2475 ( .A1(MEM_stage_inst_dmem_ram_340), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n2310) );
NOR2_X1 MEM_stage_inst_dmem_U2474 ( .A1(MEM_stage_inst_dmem_n2308), .A2(MEM_stage_inst_dmem_n2307), .ZN(MEM_stage_inst_dmem_n2316) );
NAND2_X1 MEM_stage_inst_dmem_U2473 ( .A1(MEM_stage_inst_dmem_n2306), .A2(MEM_stage_inst_dmem_n2305), .ZN(MEM_stage_inst_dmem_n2307) );
NAND2_X1 MEM_stage_inst_dmem_U2472 ( .A1(MEM_stage_inst_dmem_ram_276), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n2305) );
NAND2_X1 MEM_stage_inst_dmem_U2471 ( .A1(MEM_stage_inst_dmem_ram_4), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n2306) );
NAND2_X1 MEM_stage_inst_dmem_U2470 ( .A1(MEM_stage_inst_dmem_n2304), .A2(MEM_stage_inst_dmem_n2303), .ZN(MEM_stage_inst_dmem_n2308) );
NAND2_X1 MEM_stage_inst_dmem_U2469 ( .A1(MEM_stage_inst_dmem_ram_404), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n2303) );
NAND2_X1 MEM_stage_inst_dmem_U2468 ( .A1(MEM_stage_inst_dmem_ram_20), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n2304) );
NAND2_X1 MEM_stage_inst_dmem_U2467 ( .A1(MEM_stage_inst_dmem_n2302), .A2(MEM_stage_inst_dmem_n2301), .ZN(MEM_stage_inst_mem_read_data_3) );
NOR2_X1 MEM_stage_inst_dmem_U2466 ( .A1(MEM_stage_inst_dmem_n2300), .A2(MEM_stage_inst_dmem_n2299), .ZN(MEM_stage_inst_dmem_n2301) );
NOR2_X1 MEM_stage_inst_dmem_U2465 ( .A1(MEM_stage_inst_dmem_n2298), .A2(MEM_stage_inst_dmem_n8286), .ZN(MEM_stage_inst_dmem_n2299) );
NOR2_X1 MEM_stage_inst_dmem_U2464 ( .A1(MEM_stage_inst_dmem_n2297), .A2(MEM_stage_inst_dmem_n2296), .ZN(MEM_stage_inst_dmem_n2298) );
NAND2_X1 MEM_stage_inst_dmem_U2463 ( .A1(MEM_stage_inst_dmem_n2295), .A2(MEM_stage_inst_dmem_n2294), .ZN(MEM_stage_inst_dmem_n2296) );
NOR2_X1 MEM_stage_inst_dmem_U2462 ( .A1(MEM_stage_inst_dmem_n2293), .A2(MEM_stage_inst_dmem_n2292), .ZN(MEM_stage_inst_dmem_n2294) );
NAND2_X1 MEM_stage_inst_dmem_U2461 ( .A1(MEM_stage_inst_dmem_n2291), .A2(MEM_stage_inst_dmem_n2290), .ZN(MEM_stage_inst_dmem_n2292) );
NOR2_X1 MEM_stage_inst_dmem_U2460 ( .A1(MEM_stage_inst_dmem_n2289), .A2(MEM_stage_inst_dmem_n2288), .ZN(MEM_stage_inst_dmem_n2290) );
NAND2_X1 MEM_stage_inst_dmem_U2459 ( .A1(MEM_stage_inst_dmem_n2287), .A2(MEM_stage_inst_dmem_n2286), .ZN(MEM_stage_inst_dmem_n2288) );
NAND2_X1 MEM_stage_inst_dmem_U2458 ( .A1(MEM_stage_inst_dmem_ram_2099), .A2(MEM_stage_inst_dmem_n3103), .ZN(MEM_stage_inst_dmem_n2286) );
NAND2_X1 MEM_stage_inst_dmem_U2457 ( .A1(MEM_stage_inst_dmem_ram_2467), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n2287) );
NAND2_X1 MEM_stage_inst_dmem_U2456 ( .A1(MEM_stage_inst_dmem_n2285), .A2(MEM_stage_inst_dmem_n2284), .ZN(MEM_stage_inst_dmem_n2289) );
NAND2_X1 MEM_stage_inst_dmem_U2455 ( .A1(MEM_stage_inst_dmem_ram_2483), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n2284) );
NAND2_X1 MEM_stage_inst_dmem_U2454 ( .A1(MEM_stage_inst_dmem_ram_2275), .A2(MEM_stage_inst_dmem_n3152), .ZN(MEM_stage_inst_dmem_n2285) );
NOR2_X1 MEM_stage_inst_dmem_U2453 ( .A1(MEM_stage_inst_dmem_n2283), .A2(MEM_stage_inst_dmem_n2282), .ZN(MEM_stage_inst_dmem_n2291) );
NAND2_X1 MEM_stage_inst_dmem_U2452 ( .A1(MEM_stage_inst_dmem_n2281), .A2(MEM_stage_inst_dmem_n2280), .ZN(MEM_stage_inst_dmem_n2282) );
NAND2_X1 MEM_stage_inst_dmem_U2451 ( .A1(MEM_stage_inst_dmem_ram_2563), .A2(MEM_stage_inst_dmem_n3182), .ZN(MEM_stage_inst_dmem_n2280) );
NAND2_X1 MEM_stage_inst_dmem_U2450 ( .A1(MEM_stage_inst_dmem_ram_2707), .A2(MEM_stage_inst_dmem_n3076), .ZN(MEM_stage_inst_dmem_n2281) );
NAND2_X1 MEM_stage_inst_dmem_U2449 ( .A1(MEM_stage_inst_dmem_n2279), .A2(MEM_stage_inst_dmem_n2278), .ZN(MEM_stage_inst_dmem_n2283) );
NAND2_X1 MEM_stage_inst_dmem_U2448 ( .A1(MEM_stage_inst_dmem_ram_2755), .A2(MEM_stage_inst_dmem_n3192), .ZN(MEM_stage_inst_dmem_n2278) );
NAND2_X1 MEM_stage_inst_dmem_U2447 ( .A1(MEM_stage_inst_dmem_ram_2963), .A2(MEM_stage_inst_dmem_n3073), .ZN(MEM_stage_inst_dmem_n2279) );
NAND2_X1 MEM_stage_inst_dmem_U2446 ( .A1(MEM_stage_inst_dmem_n2277), .A2(MEM_stage_inst_dmem_n2276), .ZN(MEM_stage_inst_dmem_n2293) );
NOR2_X1 MEM_stage_inst_dmem_U2445 ( .A1(MEM_stage_inst_dmem_n2275), .A2(MEM_stage_inst_dmem_n2274), .ZN(MEM_stage_inst_dmem_n2276) );
NAND2_X1 MEM_stage_inst_dmem_U2444 ( .A1(MEM_stage_inst_dmem_n2273), .A2(MEM_stage_inst_dmem_n2272), .ZN(MEM_stage_inst_dmem_n2274) );
NAND2_X1 MEM_stage_inst_dmem_U2443 ( .A1(MEM_stage_inst_dmem_ram_2403), .A2(MEM_stage_inst_dmem_n3217), .ZN(MEM_stage_inst_dmem_n2272) );
NAND2_X1 MEM_stage_inst_dmem_U2442 ( .A1(MEM_stage_inst_dmem_ram_2419), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n2273) );
NAND2_X1 MEM_stage_inst_dmem_U2441 ( .A1(MEM_stage_inst_dmem_n2271), .A2(MEM_stage_inst_dmem_n2270), .ZN(MEM_stage_inst_dmem_n2275) );
NAND2_X1 MEM_stage_inst_dmem_U2440 ( .A1(MEM_stage_inst_dmem_ram_2195), .A2(MEM_stage_inst_dmem_n44), .ZN(MEM_stage_inst_dmem_n2270) );
NAND2_X1 MEM_stage_inst_dmem_U2439 ( .A1(MEM_stage_inst_dmem_ram_2051), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n2271) );
NOR2_X1 MEM_stage_inst_dmem_U2438 ( .A1(MEM_stage_inst_dmem_n2269), .A2(MEM_stage_inst_dmem_n2268), .ZN(MEM_stage_inst_dmem_n2277) );
NAND2_X1 MEM_stage_inst_dmem_U2437 ( .A1(MEM_stage_inst_dmem_n2267), .A2(MEM_stage_inst_dmem_n2266), .ZN(MEM_stage_inst_dmem_n2268) );
NAND2_X1 MEM_stage_inst_dmem_U2436 ( .A1(MEM_stage_inst_dmem_ram_2995), .A2(MEM_stage_inst_dmem_n3163), .ZN(MEM_stage_inst_dmem_n2266) );
NAND2_X1 MEM_stage_inst_dmem_U2435 ( .A1(MEM_stage_inst_dmem_ram_2851), .A2(MEM_stage_inst_dmem_n3137), .ZN(MEM_stage_inst_dmem_n2267) );
NAND2_X1 MEM_stage_inst_dmem_U2434 ( .A1(MEM_stage_inst_dmem_n2265), .A2(MEM_stage_inst_dmem_n2264), .ZN(MEM_stage_inst_dmem_n2269) );
NAND2_X1 MEM_stage_inst_dmem_U2433 ( .A1(MEM_stage_inst_dmem_ram_2915), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n2264) );
NAND2_X1 MEM_stage_inst_dmem_U2432 ( .A1(MEM_stage_inst_dmem_ram_2339), .A2(MEM_stage_inst_dmem_n3209), .ZN(MEM_stage_inst_dmem_n2265) );
NOR2_X1 MEM_stage_inst_dmem_U2431 ( .A1(MEM_stage_inst_dmem_n2263), .A2(MEM_stage_inst_dmem_n2262), .ZN(MEM_stage_inst_dmem_n2295) );
NAND2_X1 MEM_stage_inst_dmem_U2430 ( .A1(MEM_stage_inst_dmem_n2261), .A2(MEM_stage_inst_dmem_n2260), .ZN(MEM_stage_inst_dmem_n2262) );
NOR2_X1 MEM_stage_inst_dmem_U2429 ( .A1(MEM_stage_inst_dmem_n2259), .A2(MEM_stage_inst_dmem_n2258), .ZN(MEM_stage_inst_dmem_n2260) );
NAND2_X1 MEM_stage_inst_dmem_U2428 ( .A1(MEM_stage_inst_dmem_n2257), .A2(MEM_stage_inst_dmem_n2256), .ZN(MEM_stage_inst_dmem_n2258) );
NAND2_X1 MEM_stage_inst_dmem_U2427 ( .A1(MEM_stage_inst_dmem_ram_2371), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n2256) );
NAND2_X1 MEM_stage_inst_dmem_U2426 ( .A1(MEM_stage_inst_dmem_ram_3059), .A2(MEM_stage_inst_dmem_n3199), .ZN(MEM_stage_inst_dmem_n2257) );
NAND2_X1 MEM_stage_inst_dmem_U2425 ( .A1(MEM_stage_inst_dmem_n2255), .A2(MEM_stage_inst_dmem_n2254), .ZN(MEM_stage_inst_dmem_n2259) );
NAND2_X1 MEM_stage_inst_dmem_U2424 ( .A1(MEM_stage_inst_dmem_ram_2307), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n2254) );
NAND2_X1 MEM_stage_inst_dmem_U2423 ( .A1(MEM_stage_inst_dmem_ram_2787), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n2255) );
NOR2_X1 MEM_stage_inst_dmem_U2422 ( .A1(MEM_stage_inst_dmem_n2253), .A2(MEM_stage_inst_dmem_n2252), .ZN(MEM_stage_inst_dmem_n2261) );
NAND2_X1 MEM_stage_inst_dmem_U2421 ( .A1(MEM_stage_inst_dmem_n2251), .A2(MEM_stage_inst_dmem_n2250), .ZN(MEM_stage_inst_dmem_n2252) );
NAND2_X1 MEM_stage_inst_dmem_U2420 ( .A1(MEM_stage_inst_dmem_ram_2243), .A2(MEM_stage_inst_dmem_n3082), .ZN(MEM_stage_inst_dmem_n2250) );
NAND2_X1 MEM_stage_inst_dmem_U2419 ( .A1(MEM_stage_inst_dmem_ram_2531), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n2251) );
NAND2_X1 MEM_stage_inst_dmem_U2418 ( .A1(MEM_stage_inst_dmem_n2249), .A2(MEM_stage_inst_dmem_n2248), .ZN(MEM_stage_inst_dmem_n2253) );
NAND2_X1 MEM_stage_inst_dmem_U2417 ( .A1(MEM_stage_inst_dmem_ram_2899), .A2(MEM_stage_inst_dmem_n3141), .ZN(MEM_stage_inst_dmem_n2248) );
NAND2_X1 MEM_stage_inst_dmem_U2416 ( .A1(MEM_stage_inst_dmem_ram_2147), .A2(MEM_stage_inst_dmem_n3179), .ZN(MEM_stage_inst_dmem_n2249) );
NAND2_X1 MEM_stage_inst_dmem_U2415 ( .A1(MEM_stage_inst_dmem_n2247), .A2(MEM_stage_inst_dmem_n2246), .ZN(MEM_stage_inst_dmem_n2263) );
NOR2_X1 MEM_stage_inst_dmem_U2414 ( .A1(MEM_stage_inst_dmem_n2245), .A2(MEM_stage_inst_dmem_n2244), .ZN(MEM_stage_inst_dmem_n2246) );
NAND2_X1 MEM_stage_inst_dmem_U2413 ( .A1(MEM_stage_inst_dmem_n2243), .A2(MEM_stage_inst_dmem_n2242), .ZN(MEM_stage_inst_dmem_n2244) );
NAND2_X1 MEM_stage_inst_dmem_U2412 ( .A1(MEM_stage_inst_dmem_ram_2163), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n2242) );
NAND2_X1 MEM_stage_inst_dmem_U2411 ( .A1(MEM_stage_inst_dmem_ram_2659), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n2243) );
NAND2_X1 MEM_stage_inst_dmem_U2410 ( .A1(MEM_stage_inst_dmem_n2241), .A2(MEM_stage_inst_dmem_n2240), .ZN(MEM_stage_inst_dmem_n2245) );
NAND2_X1 MEM_stage_inst_dmem_U2409 ( .A1(MEM_stage_inst_dmem_ram_2083), .A2(MEM_stage_inst_dmem_n3092), .ZN(MEM_stage_inst_dmem_n2240) );
NAND2_X1 MEM_stage_inst_dmem_U2408 ( .A1(MEM_stage_inst_dmem_ram_2387), .A2(MEM_stage_inst_dmem_n3216), .ZN(MEM_stage_inst_dmem_n2241) );
NOR2_X1 MEM_stage_inst_dmem_U2407 ( .A1(MEM_stage_inst_dmem_n2239), .A2(MEM_stage_inst_dmem_n2238), .ZN(MEM_stage_inst_dmem_n2247) );
NAND2_X1 MEM_stage_inst_dmem_U2406 ( .A1(MEM_stage_inst_dmem_n2237), .A2(MEM_stage_inst_dmem_n2236), .ZN(MEM_stage_inst_dmem_n2238) );
NAND2_X1 MEM_stage_inst_dmem_U2405 ( .A1(MEM_stage_inst_dmem_ram_2723), .A2(MEM_stage_inst_dmem_n3155), .ZN(MEM_stage_inst_dmem_n2236) );
NAND2_X1 MEM_stage_inst_dmem_U2404 ( .A1(MEM_stage_inst_dmem_ram_2131), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n2237) );
NAND2_X1 MEM_stage_inst_dmem_U2403 ( .A1(MEM_stage_inst_dmem_n2235), .A2(MEM_stage_inst_dmem_n2234), .ZN(MEM_stage_inst_dmem_n2239) );
NAND2_X1 MEM_stage_inst_dmem_U2402 ( .A1(MEM_stage_inst_dmem_ram_2931), .A2(MEM_stage_inst_dmem_n3099), .ZN(MEM_stage_inst_dmem_n2234) );
NAND2_X1 MEM_stage_inst_dmem_U2401 ( .A1(MEM_stage_inst_dmem_ram_2211), .A2(MEM_stage_inst_dmem_n3081), .ZN(MEM_stage_inst_dmem_n2235) );
NAND2_X1 MEM_stage_inst_dmem_U2400 ( .A1(MEM_stage_inst_dmem_n2233), .A2(MEM_stage_inst_dmem_n2232), .ZN(MEM_stage_inst_dmem_n2297) );
NOR2_X1 MEM_stage_inst_dmem_U2399 ( .A1(MEM_stage_inst_dmem_n2231), .A2(MEM_stage_inst_dmem_n2230), .ZN(MEM_stage_inst_dmem_n2232) );
NAND2_X1 MEM_stage_inst_dmem_U2398 ( .A1(MEM_stage_inst_dmem_n2229), .A2(MEM_stage_inst_dmem_n2228), .ZN(MEM_stage_inst_dmem_n2230) );
NOR2_X1 MEM_stage_inst_dmem_U2397 ( .A1(MEM_stage_inst_dmem_n2227), .A2(MEM_stage_inst_dmem_n2226), .ZN(MEM_stage_inst_dmem_n2228) );
NAND2_X1 MEM_stage_inst_dmem_U2396 ( .A1(MEM_stage_inst_dmem_n2225), .A2(MEM_stage_inst_dmem_n2224), .ZN(MEM_stage_inst_dmem_n2226) );
NAND2_X1 MEM_stage_inst_dmem_U2395 ( .A1(MEM_stage_inst_dmem_ram_3043), .A2(MEM_stage_inst_dmem_n3113), .ZN(MEM_stage_inst_dmem_n2224) );
NAND2_X1 MEM_stage_inst_dmem_U2394 ( .A1(MEM_stage_inst_dmem_ram_2179), .A2(MEM_stage_inst_dmem_n3130), .ZN(MEM_stage_inst_dmem_n2225) );
NAND2_X1 MEM_stage_inst_dmem_U2393 ( .A1(MEM_stage_inst_dmem_n2223), .A2(MEM_stage_inst_dmem_n2222), .ZN(MEM_stage_inst_dmem_n2227) );
NAND2_X1 MEM_stage_inst_dmem_U2392 ( .A1(MEM_stage_inst_dmem_ram_2819), .A2(MEM_stage_inst_dmem_n37), .ZN(MEM_stage_inst_dmem_n2222) );
NAND2_X1 MEM_stage_inst_dmem_U2391 ( .A1(MEM_stage_inst_dmem_ram_2675), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n2223) );
NOR2_X1 MEM_stage_inst_dmem_U2390 ( .A1(MEM_stage_inst_dmem_n2221), .A2(MEM_stage_inst_dmem_n2220), .ZN(MEM_stage_inst_dmem_n2229) );
NAND2_X1 MEM_stage_inst_dmem_U2389 ( .A1(MEM_stage_inst_dmem_n2219), .A2(MEM_stage_inst_dmem_n2218), .ZN(MEM_stage_inst_dmem_n2220) );
NAND2_X1 MEM_stage_inst_dmem_U2388 ( .A1(MEM_stage_inst_dmem_ram_2883), .A2(MEM_stage_inst_dmem_n3120), .ZN(MEM_stage_inst_dmem_n2218) );
NAND2_X1 MEM_stage_inst_dmem_U2387 ( .A1(MEM_stage_inst_dmem_ram_2451), .A2(MEM_stage_inst_dmem_n3160), .ZN(MEM_stage_inst_dmem_n2219) );
NAND2_X1 MEM_stage_inst_dmem_U2386 ( .A1(MEM_stage_inst_dmem_n2217), .A2(MEM_stage_inst_dmem_n2216), .ZN(MEM_stage_inst_dmem_n2221) );
NAND2_X1 MEM_stage_inst_dmem_U2385 ( .A1(MEM_stage_inst_dmem_ram_2355), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n2216) );
NAND2_X1 MEM_stage_inst_dmem_U2384 ( .A1(MEM_stage_inst_dmem_ram_3027), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n2217) );
NAND2_X1 MEM_stage_inst_dmem_U2383 ( .A1(MEM_stage_inst_dmem_n2215), .A2(MEM_stage_inst_dmem_n2214), .ZN(MEM_stage_inst_dmem_n2231) );
NOR2_X1 MEM_stage_inst_dmem_U2382 ( .A1(MEM_stage_inst_dmem_n2213), .A2(MEM_stage_inst_dmem_n2212), .ZN(MEM_stage_inst_dmem_n2214) );
NAND2_X1 MEM_stage_inst_dmem_U2381 ( .A1(MEM_stage_inst_dmem_n2211), .A2(MEM_stage_inst_dmem_n2210), .ZN(MEM_stage_inst_dmem_n2212) );
NAND2_X1 MEM_stage_inst_dmem_U2380 ( .A1(MEM_stage_inst_dmem_ram_2547), .A2(MEM_stage_inst_dmem_n3170), .ZN(MEM_stage_inst_dmem_n2210) );
NAND2_X1 MEM_stage_inst_dmem_U2379 ( .A1(MEM_stage_inst_dmem_ram_2227), .A2(MEM_stage_inst_dmem_n55), .ZN(MEM_stage_inst_dmem_n2211) );
NAND2_X1 MEM_stage_inst_dmem_U2378 ( .A1(MEM_stage_inst_dmem_n2209), .A2(MEM_stage_inst_dmem_n2208), .ZN(MEM_stage_inst_dmem_n2213) );
NAND2_X1 MEM_stage_inst_dmem_U2377 ( .A1(MEM_stage_inst_dmem_ram_3011), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n2208) );
NAND2_X1 MEM_stage_inst_dmem_U2376 ( .A1(MEM_stage_inst_dmem_ram_2579), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n2209) );
NOR2_X1 MEM_stage_inst_dmem_U2375 ( .A1(MEM_stage_inst_dmem_n2207), .A2(MEM_stage_inst_dmem_n2206), .ZN(MEM_stage_inst_dmem_n2215) );
NAND2_X1 MEM_stage_inst_dmem_U2374 ( .A1(MEM_stage_inst_dmem_n2205), .A2(MEM_stage_inst_dmem_n2204), .ZN(MEM_stage_inst_dmem_n2206) );
NAND2_X1 MEM_stage_inst_dmem_U2373 ( .A1(MEM_stage_inst_dmem_ram_2979), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n2204) );
NAND2_X1 MEM_stage_inst_dmem_U2372 ( .A1(MEM_stage_inst_dmem_ram_2643), .A2(MEM_stage_inst_dmem_n3140), .ZN(MEM_stage_inst_dmem_n2205) );
NAND2_X1 MEM_stage_inst_dmem_U2371 ( .A1(MEM_stage_inst_dmem_n2203), .A2(MEM_stage_inst_dmem_n2202), .ZN(MEM_stage_inst_dmem_n2207) );
NAND2_X1 MEM_stage_inst_dmem_U2370 ( .A1(MEM_stage_inst_dmem_ram_2611), .A2(MEM_stage_inst_dmem_n3085), .ZN(MEM_stage_inst_dmem_n2202) );
NAND2_X1 MEM_stage_inst_dmem_U2369 ( .A1(MEM_stage_inst_dmem_ram_2771), .A2(MEM_stage_inst_dmem_n3112), .ZN(MEM_stage_inst_dmem_n2203) );
NOR2_X1 MEM_stage_inst_dmem_U2368 ( .A1(MEM_stage_inst_dmem_n2201), .A2(MEM_stage_inst_dmem_n2200), .ZN(MEM_stage_inst_dmem_n2233) );
NAND2_X1 MEM_stage_inst_dmem_U2367 ( .A1(MEM_stage_inst_dmem_n2199), .A2(MEM_stage_inst_dmem_n2198), .ZN(MEM_stage_inst_dmem_n2200) );
NOR2_X1 MEM_stage_inst_dmem_U2366 ( .A1(MEM_stage_inst_dmem_n2197), .A2(MEM_stage_inst_dmem_n2196), .ZN(MEM_stage_inst_dmem_n2198) );
NAND2_X1 MEM_stage_inst_dmem_U2365 ( .A1(MEM_stage_inst_dmem_n2195), .A2(MEM_stage_inst_dmem_n2194), .ZN(MEM_stage_inst_dmem_n2196) );
NAND2_X1 MEM_stage_inst_dmem_U2364 ( .A1(MEM_stage_inst_dmem_ram_2947), .A2(MEM_stage_inst_dmem_n3123), .ZN(MEM_stage_inst_dmem_n2194) );
NAND2_X1 MEM_stage_inst_dmem_U2363 ( .A1(MEM_stage_inst_dmem_ram_2835), .A2(MEM_stage_inst_dmem_n3191), .ZN(MEM_stage_inst_dmem_n2195) );
NAND2_X1 MEM_stage_inst_dmem_U2362 ( .A1(MEM_stage_inst_dmem_n2193), .A2(MEM_stage_inst_dmem_n2192), .ZN(MEM_stage_inst_dmem_n2197) );
NAND2_X1 MEM_stage_inst_dmem_U2361 ( .A1(MEM_stage_inst_dmem_ram_2803), .A2(MEM_stage_inst_dmem_n3202), .ZN(MEM_stage_inst_dmem_n2192) );
NAND2_X1 MEM_stage_inst_dmem_U2360 ( .A1(MEM_stage_inst_dmem_ram_2739), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n2193) );
NOR2_X1 MEM_stage_inst_dmem_U2359 ( .A1(MEM_stage_inst_dmem_n2191), .A2(MEM_stage_inst_dmem_n2190), .ZN(MEM_stage_inst_dmem_n2199) );
NAND2_X1 MEM_stage_inst_dmem_U2358 ( .A1(MEM_stage_inst_dmem_n2189), .A2(MEM_stage_inst_dmem_n2188), .ZN(MEM_stage_inst_dmem_n2190) );
NAND2_X1 MEM_stage_inst_dmem_U2357 ( .A1(MEM_stage_inst_dmem_ram_2291), .A2(MEM_stage_inst_dmem_n39), .ZN(MEM_stage_inst_dmem_n2188) );
NAND2_X1 MEM_stage_inst_dmem_U2356 ( .A1(MEM_stage_inst_dmem_ram_2595), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n2189) );
NAND2_X1 MEM_stage_inst_dmem_U2355 ( .A1(MEM_stage_inst_dmem_n2187), .A2(MEM_stage_inst_dmem_n2186), .ZN(MEM_stage_inst_dmem_n2191) );
NAND2_X1 MEM_stage_inst_dmem_U2354 ( .A1(MEM_stage_inst_dmem_ram_2691), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n2186) );
NAND2_X1 MEM_stage_inst_dmem_U2353 ( .A1(MEM_stage_inst_dmem_ram_2435), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n2187) );
NAND2_X1 MEM_stage_inst_dmem_U2352 ( .A1(MEM_stage_inst_dmem_n2185), .A2(MEM_stage_inst_dmem_n2184), .ZN(MEM_stage_inst_dmem_n2201) );
NOR2_X1 MEM_stage_inst_dmem_U2351 ( .A1(MEM_stage_inst_dmem_n2183), .A2(MEM_stage_inst_dmem_n2182), .ZN(MEM_stage_inst_dmem_n2184) );
NAND2_X1 MEM_stage_inst_dmem_U2350 ( .A1(MEM_stage_inst_dmem_n2181), .A2(MEM_stage_inst_dmem_n2180), .ZN(MEM_stage_inst_dmem_n2182) );
NAND2_X1 MEM_stage_inst_dmem_U2349 ( .A1(MEM_stage_inst_dmem_ram_2867), .A2(MEM_stage_inst_dmem_n46), .ZN(MEM_stage_inst_dmem_n2180) );
NAND2_X1 MEM_stage_inst_dmem_U2348 ( .A1(MEM_stage_inst_dmem_ram_2259), .A2(MEM_stage_inst_dmem_n3220), .ZN(MEM_stage_inst_dmem_n2181) );
NAND2_X1 MEM_stage_inst_dmem_U2347 ( .A1(MEM_stage_inst_dmem_n2179), .A2(MEM_stage_inst_dmem_n2178), .ZN(MEM_stage_inst_dmem_n2183) );
NAND2_X1 MEM_stage_inst_dmem_U2346 ( .A1(MEM_stage_inst_dmem_ram_2515), .A2(MEM_stage_inst_dmem_n3174), .ZN(MEM_stage_inst_dmem_n2178) );
NAND2_X1 MEM_stage_inst_dmem_U2345 ( .A1(MEM_stage_inst_dmem_ram_2627), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n2179) );
NOR2_X1 MEM_stage_inst_dmem_U2344 ( .A1(MEM_stage_inst_dmem_n2177), .A2(MEM_stage_inst_dmem_n2176), .ZN(MEM_stage_inst_dmem_n2185) );
NAND2_X1 MEM_stage_inst_dmem_U2343 ( .A1(MEM_stage_inst_dmem_n2175), .A2(MEM_stage_inst_dmem_n2174), .ZN(MEM_stage_inst_dmem_n2176) );
NAND2_X1 MEM_stage_inst_dmem_U2342 ( .A1(MEM_stage_inst_dmem_ram_2115), .A2(MEM_stage_inst_dmem_n3102), .ZN(MEM_stage_inst_dmem_n2174) );
NAND2_X1 MEM_stage_inst_dmem_U2341 ( .A1(MEM_stage_inst_dmem_ram_2067), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n2175) );
NAND2_X1 MEM_stage_inst_dmem_U2340 ( .A1(MEM_stage_inst_dmem_n2173), .A2(MEM_stage_inst_dmem_n2172), .ZN(MEM_stage_inst_dmem_n2177) );
NAND2_X1 MEM_stage_inst_dmem_U2339 ( .A1(MEM_stage_inst_dmem_ram_2323), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n2172) );
NAND2_X1 MEM_stage_inst_dmem_U2338 ( .A1(MEM_stage_inst_dmem_ram_2499), .A2(MEM_stage_inst_dmem_n3173), .ZN(MEM_stage_inst_dmem_n2173) );
NOR2_X1 MEM_stage_inst_dmem_U2337 ( .A1(MEM_stage_inst_dmem_n2171), .A2(MEM_stage_inst_dmem_n8551), .ZN(MEM_stage_inst_dmem_n2300) );
NOR2_X1 MEM_stage_inst_dmem_U2336 ( .A1(MEM_stage_inst_dmem_n2170), .A2(MEM_stage_inst_dmem_n2169), .ZN(MEM_stage_inst_dmem_n2171) );
NAND2_X1 MEM_stage_inst_dmem_U2335 ( .A1(MEM_stage_inst_dmem_n2168), .A2(MEM_stage_inst_dmem_n2167), .ZN(MEM_stage_inst_dmem_n2169) );
NOR2_X1 MEM_stage_inst_dmem_U2334 ( .A1(MEM_stage_inst_dmem_n2166), .A2(MEM_stage_inst_dmem_n2165), .ZN(MEM_stage_inst_dmem_n2167) );
NAND2_X1 MEM_stage_inst_dmem_U2333 ( .A1(MEM_stage_inst_dmem_n2164), .A2(MEM_stage_inst_dmem_n2163), .ZN(MEM_stage_inst_dmem_n2165) );
NOR2_X1 MEM_stage_inst_dmem_U2332 ( .A1(MEM_stage_inst_dmem_n2162), .A2(MEM_stage_inst_dmem_n2161), .ZN(MEM_stage_inst_dmem_n2163) );
NAND2_X1 MEM_stage_inst_dmem_U2331 ( .A1(MEM_stage_inst_dmem_n2160), .A2(MEM_stage_inst_dmem_n2159), .ZN(MEM_stage_inst_dmem_n2161) );
NAND2_X1 MEM_stage_inst_dmem_U2330 ( .A1(MEM_stage_inst_dmem_ram_867), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n2159) );
NAND2_X1 MEM_stage_inst_dmem_U2329 ( .A1(MEM_stage_inst_dmem_ram_947), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n2160) );
NAND2_X1 MEM_stage_inst_dmem_U2328 ( .A1(MEM_stage_inst_dmem_n2158), .A2(MEM_stage_inst_dmem_n2157), .ZN(MEM_stage_inst_dmem_n2162) );
NAND2_X1 MEM_stage_inst_dmem_U2327 ( .A1(MEM_stage_inst_dmem_ram_979), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n2157) );
NAND2_X1 MEM_stage_inst_dmem_U2326 ( .A1(MEM_stage_inst_dmem_ram_371), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n2158) );
NOR2_X1 MEM_stage_inst_dmem_U2325 ( .A1(MEM_stage_inst_dmem_n2156), .A2(MEM_stage_inst_dmem_n2155), .ZN(MEM_stage_inst_dmem_n2164) );
NAND2_X1 MEM_stage_inst_dmem_U2324 ( .A1(MEM_stage_inst_dmem_n2154), .A2(MEM_stage_inst_dmem_n2153), .ZN(MEM_stage_inst_dmem_n2155) );
NAND2_X1 MEM_stage_inst_dmem_U2323 ( .A1(MEM_stage_inst_dmem_ram_291), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n2153) );
NAND2_X1 MEM_stage_inst_dmem_U2322 ( .A1(MEM_stage_inst_dmem_ram_531), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n2154) );
NAND2_X1 MEM_stage_inst_dmem_U2321 ( .A1(MEM_stage_inst_dmem_n2152), .A2(MEM_stage_inst_dmem_n2151), .ZN(MEM_stage_inst_dmem_n2156) );
NAND2_X1 MEM_stage_inst_dmem_U2320 ( .A1(MEM_stage_inst_dmem_ram_643), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n2151) );
NAND2_X1 MEM_stage_inst_dmem_U2319 ( .A1(MEM_stage_inst_dmem_ram_755), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n2152) );
NAND2_X1 MEM_stage_inst_dmem_U2318 ( .A1(MEM_stage_inst_dmem_n2150), .A2(MEM_stage_inst_dmem_n2149), .ZN(MEM_stage_inst_dmem_n2166) );
NOR2_X1 MEM_stage_inst_dmem_U2317 ( .A1(MEM_stage_inst_dmem_n2148), .A2(MEM_stage_inst_dmem_n2147), .ZN(MEM_stage_inst_dmem_n2149) );
NAND2_X1 MEM_stage_inst_dmem_U2316 ( .A1(MEM_stage_inst_dmem_n2146), .A2(MEM_stage_inst_dmem_n2145), .ZN(MEM_stage_inst_dmem_n2147) );
NAND2_X1 MEM_stage_inst_dmem_U2315 ( .A1(MEM_stage_inst_dmem_ram_131), .A2(MEM_stage_inst_dmem_n61), .ZN(MEM_stage_inst_dmem_n2145) );
NAND2_X1 MEM_stage_inst_dmem_U2314 ( .A1(MEM_stage_inst_dmem_ram_547), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n2146) );
NAND2_X1 MEM_stage_inst_dmem_U2313 ( .A1(MEM_stage_inst_dmem_n2144), .A2(MEM_stage_inst_dmem_n2143), .ZN(MEM_stage_inst_dmem_n2148) );
NAND2_X1 MEM_stage_inst_dmem_U2312 ( .A1(MEM_stage_inst_dmem_ram_883), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n2143) );
NAND2_X1 MEM_stage_inst_dmem_U2311 ( .A1(MEM_stage_inst_dmem_ram_899), .A2(MEM_stage_inst_dmem_n72), .ZN(MEM_stage_inst_dmem_n2144) );
NOR2_X1 MEM_stage_inst_dmem_U2310 ( .A1(MEM_stage_inst_dmem_n2142), .A2(MEM_stage_inst_dmem_n2141), .ZN(MEM_stage_inst_dmem_n2150) );
NAND2_X1 MEM_stage_inst_dmem_U2309 ( .A1(MEM_stage_inst_dmem_n2140), .A2(MEM_stage_inst_dmem_n2139), .ZN(MEM_stage_inst_dmem_n2141) );
NAND2_X1 MEM_stage_inst_dmem_U2308 ( .A1(MEM_stage_inst_dmem_ram_771), .A2(MEM_stage_inst_dmem_n37), .ZN(MEM_stage_inst_dmem_n2139) );
NAND2_X1 MEM_stage_inst_dmem_U2307 ( .A1(MEM_stage_inst_dmem_ram_275), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n2140) );
NAND2_X1 MEM_stage_inst_dmem_U2306 ( .A1(MEM_stage_inst_dmem_n2138), .A2(MEM_stage_inst_dmem_n2137), .ZN(MEM_stage_inst_dmem_n2142) );
NAND2_X1 MEM_stage_inst_dmem_U2305 ( .A1(MEM_stage_inst_dmem_ram_435), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n2137) );
NAND2_X1 MEM_stage_inst_dmem_U2304 ( .A1(MEM_stage_inst_dmem_ram_227), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n2138) );
NOR2_X1 MEM_stage_inst_dmem_U2303 ( .A1(MEM_stage_inst_dmem_n2136), .A2(MEM_stage_inst_dmem_n2135), .ZN(MEM_stage_inst_dmem_n2168) );
NAND2_X1 MEM_stage_inst_dmem_U2302 ( .A1(MEM_stage_inst_dmem_n2134), .A2(MEM_stage_inst_dmem_n2133), .ZN(MEM_stage_inst_dmem_n2135) );
NOR2_X1 MEM_stage_inst_dmem_U2301 ( .A1(MEM_stage_inst_dmem_n2132), .A2(MEM_stage_inst_dmem_n2131), .ZN(MEM_stage_inst_dmem_n2133) );
NAND2_X1 MEM_stage_inst_dmem_U2300 ( .A1(MEM_stage_inst_dmem_n2130), .A2(MEM_stage_inst_dmem_n2129), .ZN(MEM_stage_inst_dmem_n2131) );
NAND2_X1 MEM_stage_inst_dmem_U2299 ( .A1(MEM_stage_inst_dmem_ram_355), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n2129) );
NAND2_X1 MEM_stage_inst_dmem_U2298 ( .A1(MEM_stage_inst_dmem_ram_115), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n2130) );
NAND2_X1 MEM_stage_inst_dmem_U2297 ( .A1(MEM_stage_inst_dmem_n2128), .A2(MEM_stage_inst_dmem_n2127), .ZN(MEM_stage_inst_dmem_n2132) );
NAND2_X1 MEM_stage_inst_dmem_U2296 ( .A1(MEM_stage_inst_dmem_ram_963), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n2127) );
NAND2_X1 MEM_stage_inst_dmem_U2295 ( .A1(MEM_stage_inst_dmem_ram_595), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n2128) );
NOR2_X1 MEM_stage_inst_dmem_U2294 ( .A1(MEM_stage_inst_dmem_n2126), .A2(MEM_stage_inst_dmem_n2125), .ZN(MEM_stage_inst_dmem_n2134) );
NAND2_X1 MEM_stage_inst_dmem_U2293 ( .A1(MEM_stage_inst_dmem_n2124), .A2(MEM_stage_inst_dmem_n2123), .ZN(MEM_stage_inst_dmem_n2125) );
NAND2_X1 MEM_stage_inst_dmem_U2292 ( .A1(MEM_stage_inst_dmem_ram_195), .A2(MEM_stage_inst_dmem_n36), .ZN(MEM_stage_inst_dmem_n2123) );
NAND2_X1 MEM_stage_inst_dmem_U2291 ( .A1(MEM_stage_inst_dmem_ram_739), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n2124) );
NAND2_X1 MEM_stage_inst_dmem_U2290 ( .A1(MEM_stage_inst_dmem_n2122), .A2(MEM_stage_inst_dmem_n2121), .ZN(MEM_stage_inst_dmem_n2126) );
NAND2_X1 MEM_stage_inst_dmem_U2289 ( .A1(MEM_stage_inst_dmem_ram_835), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n2121) );
NAND2_X1 MEM_stage_inst_dmem_U2288 ( .A1(MEM_stage_inst_dmem_ram_995), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n2122) );
NAND2_X1 MEM_stage_inst_dmem_U2287 ( .A1(MEM_stage_inst_dmem_n2120), .A2(MEM_stage_inst_dmem_n2119), .ZN(MEM_stage_inst_dmem_n2136) );
NOR2_X1 MEM_stage_inst_dmem_U2286 ( .A1(MEM_stage_inst_dmem_n2118), .A2(MEM_stage_inst_dmem_n2117), .ZN(MEM_stage_inst_dmem_n2119) );
NAND2_X1 MEM_stage_inst_dmem_U2285 ( .A1(MEM_stage_inst_dmem_n2116), .A2(MEM_stage_inst_dmem_n2115), .ZN(MEM_stage_inst_dmem_n2117) );
NAND2_X1 MEM_stage_inst_dmem_U2284 ( .A1(MEM_stage_inst_dmem_ram_163), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n2115) );
NAND2_X1 MEM_stage_inst_dmem_U2283 ( .A1(MEM_stage_inst_dmem_ram_339), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n2116) );
NAND2_X1 MEM_stage_inst_dmem_U2282 ( .A1(MEM_stage_inst_dmem_n2114), .A2(MEM_stage_inst_dmem_n2113), .ZN(MEM_stage_inst_dmem_n2118) );
NAND2_X1 MEM_stage_inst_dmem_U2281 ( .A1(MEM_stage_inst_dmem_ram_403), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n2113) );
NAND2_X1 MEM_stage_inst_dmem_U2280 ( .A1(MEM_stage_inst_dmem_ram_675), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n2114) );
NOR2_X1 MEM_stage_inst_dmem_U2279 ( .A1(MEM_stage_inst_dmem_n2112), .A2(MEM_stage_inst_dmem_n2111), .ZN(MEM_stage_inst_dmem_n2120) );
NAND2_X1 MEM_stage_inst_dmem_U2278 ( .A1(MEM_stage_inst_dmem_n2110), .A2(MEM_stage_inst_dmem_n2109), .ZN(MEM_stage_inst_dmem_n2111) );
NAND2_X1 MEM_stage_inst_dmem_U2277 ( .A1(MEM_stage_inst_dmem_ram_307), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n2109) );
NAND2_X1 MEM_stage_inst_dmem_U2276 ( .A1(MEM_stage_inst_dmem_ram_51), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n2110) );
NAND2_X1 MEM_stage_inst_dmem_U2275 ( .A1(MEM_stage_inst_dmem_n2108), .A2(MEM_stage_inst_dmem_n2107), .ZN(MEM_stage_inst_dmem_n2112) );
NAND2_X1 MEM_stage_inst_dmem_U2274 ( .A1(MEM_stage_inst_dmem_ram_467), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n2107) );
NAND2_X1 MEM_stage_inst_dmem_U2273 ( .A1(MEM_stage_inst_dmem_ram_931), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n2108) );
NAND2_X1 MEM_stage_inst_dmem_U2272 ( .A1(MEM_stage_inst_dmem_n2106), .A2(MEM_stage_inst_dmem_n2105), .ZN(MEM_stage_inst_dmem_n2170) );
NOR2_X1 MEM_stage_inst_dmem_U2271 ( .A1(MEM_stage_inst_dmem_n2104), .A2(MEM_stage_inst_dmem_n2103), .ZN(MEM_stage_inst_dmem_n2105) );
NAND2_X1 MEM_stage_inst_dmem_U2270 ( .A1(MEM_stage_inst_dmem_n2102), .A2(MEM_stage_inst_dmem_n2101), .ZN(MEM_stage_inst_dmem_n2103) );
NOR2_X1 MEM_stage_inst_dmem_U2269 ( .A1(MEM_stage_inst_dmem_n2100), .A2(MEM_stage_inst_dmem_n2099), .ZN(MEM_stage_inst_dmem_n2101) );
NAND2_X1 MEM_stage_inst_dmem_U2268 ( .A1(MEM_stage_inst_dmem_n2098), .A2(MEM_stage_inst_dmem_n2097), .ZN(MEM_stage_inst_dmem_n2099) );
NAND2_X1 MEM_stage_inst_dmem_U2267 ( .A1(MEM_stage_inst_dmem_ram_691), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n2097) );
NAND2_X1 MEM_stage_inst_dmem_U2266 ( .A1(MEM_stage_inst_dmem_ram_451), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n2098) );
NAND2_X1 MEM_stage_inst_dmem_U2265 ( .A1(MEM_stage_inst_dmem_n2096), .A2(MEM_stage_inst_dmem_n2095), .ZN(MEM_stage_inst_dmem_n2100) );
NAND2_X1 MEM_stage_inst_dmem_U2264 ( .A1(MEM_stage_inst_dmem_ram_787), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n2095) );
NAND2_X1 MEM_stage_inst_dmem_U2263 ( .A1(MEM_stage_inst_dmem_ram_99), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n2096) );
NOR2_X1 MEM_stage_inst_dmem_U2262 ( .A1(MEM_stage_inst_dmem_n2094), .A2(MEM_stage_inst_dmem_n2093), .ZN(MEM_stage_inst_dmem_n2102) );
NAND2_X1 MEM_stage_inst_dmem_U2261 ( .A1(MEM_stage_inst_dmem_n2092), .A2(MEM_stage_inst_dmem_n2091), .ZN(MEM_stage_inst_dmem_n2093) );
NAND2_X1 MEM_stage_inst_dmem_U2260 ( .A1(MEM_stage_inst_dmem_ram_323), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n2091) );
NAND2_X1 MEM_stage_inst_dmem_U2259 ( .A1(MEM_stage_inst_dmem_ram_707), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n2092) );
NAND2_X1 MEM_stage_inst_dmem_U2258 ( .A1(MEM_stage_inst_dmem_n2090), .A2(MEM_stage_inst_dmem_n2089), .ZN(MEM_stage_inst_dmem_n2094) );
NAND2_X1 MEM_stage_inst_dmem_U2257 ( .A1(MEM_stage_inst_dmem_ram_819), .A2(MEM_stage_inst_dmem_n46), .ZN(MEM_stage_inst_dmem_n2089) );
NAND2_X1 MEM_stage_inst_dmem_U2256 ( .A1(MEM_stage_inst_dmem_ram_259), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n2090) );
NAND2_X1 MEM_stage_inst_dmem_U2255 ( .A1(MEM_stage_inst_dmem_n2088), .A2(MEM_stage_inst_dmem_n2087), .ZN(MEM_stage_inst_dmem_n2104) );
NOR2_X1 MEM_stage_inst_dmem_U2254 ( .A1(MEM_stage_inst_dmem_n2086), .A2(MEM_stage_inst_dmem_n2085), .ZN(MEM_stage_inst_dmem_n2087) );
NAND2_X1 MEM_stage_inst_dmem_U2253 ( .A1(MEM_stage_inst_dmem_n2084), .A2(MEM_stage_inst_dmem_n2083), .ZN(MEM_stage_inst_dmem_n2085) );
NAND2_X1 MEM_stage_inst_dmem_U2252 ( .A1(MEM_stage_inst_dmem_ram_243), .A2(MEM_stage_inst_dmem_n39), .ZN(MEM_stage_inst_dmem_n2083) );
NAND2_X1 MEM_stage_inst_dmem_U2251 ( .A1(MEM_stage_inst_dmem_ram_611), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n2084) );
NAND2_X1 MEM_stage_inst_dmem_U2250 ( .A1(MEM_stage_inst_dmem_n2082), .A2(MEM_stage_inst_dmem_n2081), .ZN(MEM_stage_inst_dmem_n2086) );
NAND2_X1 MEM_stage_inst_dmem_U2249 ( .A1(MEM_stage_inst_dmem_ram_563), .A2(MEM_stage_inst_dmem_n41), .ZN(MEM_stage_inst_dmem_n2081) );
NAND2_X1 MEM_stage_inst_dmem_U2248 ( .A1(MEM_stage_inst_dmem_ram_723), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n2082) );
NOR2_X1 MEM_stage_inst_dmem_U2247 ( .A1(MEM_stage_inst_dmem_n2080), .A2(MEM_stage_inst_dmem_n2079), .ZN(MEM_stage_inst_dmem_n2088) );
NAND2_X1 MEM_stage_inst_dmem_U2246 ( .A1(MEM_stage_inst_dmem_n2078), .A2(MEM_stage_inst_dmem_n2077), .ZN(MEM_stage_inst_dmem_n2079) );
NAND2_X1 MEM_stage_inst_dmem_U2245 ( .A1(MEM_stage_inst_dmem_ram_387), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n2077) );
NAND2_X1 MEM_stage_inst_dmem_U2244 ( .A1(MEM_stage_inst_dmem_ram_627), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n2078) );
NAND2_X1 MEM_stage_inst_dmem_U2243 ( .A1(MEM_stage_inst_dmem_n2076), .A2(MEM_stage_inst_dmem_n2075), .ZN(MEM_stage_inst_dmem_n2080) );
NAND2_X1 MEM_stage_inst_dmem_U2242 ( .A1(MEM_stage_inst_dmem_ram_35), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n2075) );
NAND2_X1 MEM_stage_inst_dmem_U2241 ( .A1(MEM_stage_inst_dmem_ram_147), .A2(MEM_stage_inst_dmem_n44), .ZN(MEM_stage_inst_dmem_n2076) );
NOR2_X1 MEM_stage_inst_dmem_U2240 ( .A1(MEM_stage_inst_dmem_n2074), .A2(MEM_stage_inst_dmem_n2073), .ZN(MEM_stage_inst_dmem_n2106) );
NAND2_X1 MEM_stage_inst_dmem_U2239 ( .A1(MEM_stage_inst_dmem_n2072), .A2(MEM_stage_inst_dmem_n2071), .ZN(MEM_stage_inst_dmem_n2073) );
NOR2_X1 MEM_stage_inst_dmem_U2238 ( .A1(MEM_stage_inst_dmem_n2070), .A2(MEM_stage_inst_dmem_n2069), .ZN(MEM_stage_inst_dmem_n2071) );
NAND2_X1 MEM_stage_inst_dmem_U2237 ( .A1(MEM_stage_inst_dmem_n2068), .A2(MEM_stage_inst_dmem_n2067), .ZN(MEM_stage_inst_dmem_n2069) );
NAND2_X1 MEM_stage_inst_dmem_U2236 ( .A1(MEM_stage_inst_dmem_ram_851), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n2067) );
NAND2_X1 MEM_stage_inst_dmem_U2235 ( .A1(MEM_stage_inst_dmem_ram_83), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n2068) );
NAND2_X1 MEM_stage_inst_dmem_U2234 ( .A1(MEM_stage_inst_dmem_n2066), .A2(MEM_stage_inst_dmem_n2065), .ZN(MEM_stage_inst_dmem_n2070) );
NAND2_X1 MEM_stage_inst_dmem_U2233 ( .A1(MEM_stage_inst_dmem_ram_67), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n2065) );
NAND2_X1 MEM_stage_inst_dmem_U2232 ( .A1(MEM_stage_inst_dmem_ram_1011), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n2066) );
NOR2_X1 MEM_stage_inst_dmem_U2231 ( .A1(MEM_stage_inst_dmem_n2064), .A2(MEM_stage_inst_dmem_n2063), .ZN(MEM_stage_inst_dmem_n2072) );
NAND2_X1 MEM_stage_inst_dmem_U2230 ( .A1(MEM_stage_inst_dmem_n2062), .A2(MEM_stage_inst_dmem_n2061), .ZN(MEM_stage_inst_dmem_n2063) );
NAND2_X1 MEM_stage_inst_dmem_U2229 ( .A1(MEM_stage_inst_dmem_ram_3), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n2061) );
NAND2_X1 MEM_stage_inst_dmem_U2228 ( .A1(MEM_stage_inst_dmem_ram_579), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n2062) );
NAND2_X1 MEM_stage_inst_dmem_U2227 ( .A1(MEM_stage_inst_dmem_n2060), .A2(MEM_stage_inst_dmem_n2059), .ZN(MEM_stage_inst_dmem_n2064) );
NAND2_X1 MEM_stage_inst_dmem_U2226 ( .A1(MEM_stage_inst_dmem_ram_803), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n2059) );
NAND2_X1 MEM_stage_inst_dmem_U2225 ( .A1(MEM_stage_inst_dmem_ram_515), .A2(MEM_stage_inst_dmem_n71), .ZN(MEM_stage_inst_dmem_n2060) );
NAND2_X1 MEM_stage_inst_dmem_U2224 ( .A1(MEM_stage_inst_dmem_n2058), .A2(MEM_stage_inst_dmem_n2057), .ZN(MEM_stage_inst_dmem_n2074) );
NOR2_X1 MEM_stage_inst_dmem_U2223 ( .A1(MEM_stage_inst_dmem_n2056), .A2(MEM_stage_inst_dmem_n2055), .ZN(MEM_stage_inst_dmem_n2057) );
NAND2_X1 MEM_stage_inst_dmem_U2222 ( .A1(MEM_stage_inst_dmem_n2054), .A2(MEM_stage_inst_dmem_n2053), .ZN(MEM_stage_inst_dmem_n2055) );
NAND2_X1 MEM_stage_inst_dmem_U2221 ( .A1(MEM_stage_inst_dmem_ram_915), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n2053) );
NAND2_X1 MEM_stage_inst_dmem_U2220 ( .A1(MEM_stage_inst_dmem_ram_179), .A2(MEM_stage_inst_dmem_n55), .ZN(MEM_stage_inst_dmem_n2054) );
NAND2_X1 MEM_stage_inst_dmem_U2219 ( .A1(MEM_stage_inst_dmem_n2052), .A2(MEM_stage_inst_dmem_n2051), .ZN(MEM_stage_inst_dmem_n2056) );
NAND2_X1 MEM_stage_inst_dmem_U2218 ( .A1(MEM_stage_inst_dmem_ram_19), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n2051) );
NAND2_X1 MEM_stage_inst_dmem_U2217 ( .A1(MEM_stage_inst_dmem_ram_659), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n2052) );
NOR2_X1 MEM_stage_inst_dmem_U2216 ( .A1(MEM_stage_inst_dmem_n2050), .A2(MEM_stage_inst_dmem_n2049), .ZN(MEM_stage_inst_dmem_n2058) );
NAND2_X1 MEM_stage_inst_dmem_U2215 ( .A1(MEM_stage_inst_dmem_n2048), .A2(MEM_stage_inst_dmem_n2047), .ZN(MEM_stage_inst_dmem_n2049) );
NAND2_X1 MEM_stage_inst_dmem_U2214 ( .A1(MEM_stage_inst_dmem_ram_499), .A2(MEM_stage_inst_dmem_n8535), .ZN(MEM_stage_inst_dmem_n2047) );
NAND2_X1 MEM_stage_inst_dmem_U2213 ( .A1(MEM_stage_inst_dmem_ram_419), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n2048) );
NAND2_X1 MEM_stage_inst_dmem_U2212 ( .A1(MEM_stage_inst_dmem_n2046), .A2(MEM_stage_inst_dmem_n2045), .ZN(MEM_stage_inst_dmem_n2050) );
NAND2_X1 MEM_stage_inst_dmem_U2211 ( .A1(MEM_stage_inst_dmem_ram_483), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n2045) );
NAND2_X1 MEM_stage_inst_dmem_U2210 ( .A1(MEM_stage_inst_dmem_ram_211), .A2(MEM_stage_inst_dmem_n51), .ZN(MEM_stage_inst_dmem_n2046) );
NOR2_X1 MEM_stage_inst_dmem_U2209 ( .A1(MEM_stage_inst_dmem_n2044), .A2(MEM_stage_inst_dmem_n2043), .ZN(MEM_stage_inst_dmem_n2302) );
NOR2_X1 MEM_stage_inst_dmem_U2208 ( .A1(MEM_stage_inst_dmem_n2042), .A2(MEM_stage_inst_dmem_n8417), .ZN(MEM_stage_inst_dmem_n2043) );
NOR2_X1 MEM_stage_inst_dmem_U2207 ( .A1(MEM_stage_inst_dmem_n2041), .A2(MEM_stage_inst_dmem_n2040), .ZN(MEM_stage_inst_dmem_n2042) );
NAND2_X1 MEM_stage_inst_dmem_U2206 ( .A1(MEM_stage_inst_dmem_n2039), .A2(MEM_stage_inst_dmem_n2038), .ZN(MEM_stage_inst_dmem_n2040) );
NOR2_X1 MEM_stage_inst_dmem_U2205 ( .A1(MEM_stage_inst_dmem_n2037), .A2(MEM_stage_inst_dmem_n2036), .ZN(MEM_stage_inst_dmem_n2038) );
NAND2_X1 MEM_stage_inst_dmem_U2204 ( .A1(MEM_stage_inst_dmem_n2035), .A2(MEM_stage_inst_dmem_n2034), .ZN(MEM_stage_inst_dmem_n2036) );
NOR2_X1 MEM_stage_inst_dmem_U2203 ( .A1(MEM_stage_inst_dmem_n2033), .A2(MEM_stage_inst_dmem_n2032), .ZN(MEM_stage_inst_dmem_n2034) );
NAND2_X1 MEM_stage_inst_dmem_U2202 ( .A1(MEM_stage_inst_dmem_n2031), .A2(MEM_stage_inst_dmem_n2030), .ZN(MEM_stage_inst_dmem_n2032) );
NAND2_X1 MEM_stage_inst_dmem_U2201 ( .A1(MEM_stage_inst_dmem_ram_3427), .A2(MEM_stage_inst_dmem_n3217), .ZN(MEM_stage_inst_dmem_n2030) );
NAND2_X1 MEM_stage_inst_dmem_U2200 ( .A1(MEM_stage_inst_dmem_ram_3107), .A2(MEM_stage_inst_dmem_n3092), .ZN(MEM_stage_inst_dmem_n2031) );
NAND2_X1 MEM_stage_inst_dmem_U2199 ( .A1(MEM_stage_inst_dmem_n2029), .A2(MEM_stage_inst_dmem_n2028), .ZN(MEM_stage_inst_dmem_n2033) );
NAND2_X1 MEM_stage_inst_dmem_U2198 ( .A1(MEM_stage_inst_dmem_ram_4019), .A2(MEM_stage_inst_dmem_n3163), .ZN(MEM_stage_inst_dmem_n2028) );
NAND2_X1 MEM_stage_inst_dmem_U2197 ( .A1(MEM_stage_inst_dmem_ram_3283), .A2(MEM_stage_inst_dmem_n3220), .ZN(MEM_stage_inst_dmem_n2029) );
NOR2_X1 MEM_stage_inst_dmem_U2196 ( .A1(MEM_stage_inst_dmem_n2027), .A2(MEM_stage_inst_dmem_n2026), .ZN(MEM_stage_inst_dmem_n2035) );
NAND2_X1 MEM_stage_inst_dmem_U2195 ( .A1(MEM_stage_inst_dmem_n2025), .A2(MEM_stage_inst_dmem_n2024), .ZN(MEM_stage_inst_dmem_n2026) );
NAND2_X1 MEM_stage_inst_dmem_U2194 ( .A1(MEM_stage_inst_dmem_ram_3939), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n2024) );
NAND2_X1 MEM_stage_inst_dmem_U2193 ( .A1(MEM_stage_inst_dmem_ram_3891), .A2(MEM_stage_inst_dmem_n8005), .ZN(MEM_stage_inst_dmem_n2025) );
NAND2_X1 MEM_stage_inst_dmem_U2192 ( .A1(MEM_stage_inst_dmem_n2023), .A2(MEM_stage_inst_dmem_n2022), .ZN(MEM_stage_inst_dmem_n2027) );
NAND2_X1 MEM_stage_inst_dmem_U2191 ( .A1(MEM_stage_inst_dmem_ram_3459), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n2022) );
NAND2_X1 MEM_stage_inst_dmem_U2190 ( .A1(MEM_stage_inst_dmem_ram_3251), .A2(MEM_stage_inst_dmem_n55), .ZN(MEM_stage_inst_dmem_n2023) );
NAND2_X1 MEM_stage_inst_dmem_U2189 ( .A1(MEM_stage_inst_dmem_n2021), .A2(MEM_stage_inst_dmem_n2020), .ZN(MEM_stage_inst_dmem_n2037) );
NOR2_X1 MEM_stage_inst_dmem_U2188 ( .A1(MEM_stage_inst_dmem_n2019), .A2(MEM_stage_inst_dmem_n2018), .ZN(MEM_stage_inst_dmem_n2020) );
NAND2_X1 MEM_stage_inst_dmem_U2187 ( .A1(MEM_stage_inst_dmem_n2017), .A2(MEM_stage_inst_dmem_n2016), .ZN(MEM_stage_inst_dmem_n2018) );
NAND2_X1 MEM_stage_inst_dmem_U2186 ( .A1(MEM_stage_inst_dmem_ram_3955), .A2(MEM_stage_inst_dmem_n3099), .ZN(MEM_stage_inst_dmem_n2016) );
NAND2_X1 MEM_stage_inst_dmem_U2185 ( .A1(MEM_stage_inst_dmem_ram_3523), .A2(MEM_stage_inst_dmem_n3173), .ZN(MEM_stage_inst_dmem_n2017) );
NAND2_X1 MEM_stage_inst_dmem_U2184 ( .A1(MEM_stage_inst_dmem_n2015), .A2(MEM_stage_inst_dmem_n2014), .ZN(MEM_stage_inst_dmem_n2019) );
NAND2_X1 MEM_stage_inst_dmem_U2183 ( .A1(MEM_stage_inst_dmem_ram_3235), .A2(MEM_stage_inst_dmem_n3081), .ZN(MEM_stage_inst_dmem_n2014) );
NAND2_X1 MEM_stage_inst_dmem_U2182 ( .A1(MEM_stage_inst_dmem_ram_3171), .A2(MEM_stage_inst_dmem_n3179), .ZN(MEM_stage_inst_dmem_n2015) );
NOR2_X1 MEM_stage_inst_dmem_U2181 ( .A1(MEM_stage_inst_dmem_n2013), .A2(MEM_stage_inst_dmem_n2012), .ZN(MEM_stage_inst_dmem_n2021) );
NAND2_X1 MEM_stage_inst_dmem_U2180 ( .A1(MEM_stage_inst_dmem_n2011), .A2(MEM_stage_inst_dmem_n2010), .ZN(MEM_stage_inst_dmem_n2012) );
NAND2_X1 MEM_stage_inst_dmem_U2179 ( .A1(MEM_stage_inst_dmem_ram_3379), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n2010) );
NAND2_X1 MEM_stage_inst_dmem_U2178 ( .A1(MEM_stage_inst_dmem_ram_3875), .A2(MEM_stage_inst_dmem_n3137), .ZN(MEM_stage_inst_dmem_n2011) );
NAND2_X1 MEM_stage_inst_dmem_U2177 ( .A1(MEM_stage_inst_dmem_n2009), .A2(MEM_stage_inst_dmem_n2008), .ZN(MEM_stage_inst_dmem_n2013) );
NAND2_X1 MEM_stage_inst_dmem_U2176 ( .A1(MEM_stage_inst_dmem_ram_3315), .A2(MEM_stage_inst_dmem_n7914), .ZN(MEM_stage_inst_dmem_n2008) );
NAND2_X1 MEM_stage_inst_dmem_U2175 ( .A1(MEM_stage_inst_dmem_ram_3347), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n2009) );
NOR2_X1 MEM_stage_inst_dmem_U2174 ( .A1(MEM_stage_inst_dmem_n2007), .A2(MEM_stage_inst_dmem_n2006), .ZN(MEM_stage_inst_dmem_n2039) );
NAND2_X1 MEM_stage_inst_dmem_U2173 ( .A1(MEM_stage_inst_dmem_n2005), .A2(MEM_stage_inst_dmem_n2004), .ZN(MEM_stage_inst_dmem_n2006) );
NOR2_X1 MEM_stage_inst_dmem_U2172 ( .A1(MEM_stage_inst_dmem_n2003), .A2(MEM_stage_inst_dmem_n2002), .ZN(MEM_stage_inst_dmem_n2004) );
NAND2_X1 MEM_stage_inst_dmem_U2171 ( .A1(MEM_stage_inst_dmem_n2001), .A2(MEM_stage_inst_dmem_n2000), .ZN(MEM_stage_inst_dmem_n2002) );
NAND2_X1 MEM_stage_inst_dmem_U2170 ( .A1(MEM_stage_inst_dmem_ram_3555), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n2000) );
NAND2_X1 MEM_stage_inst_dmem_U2169 ( .A1(MEM_stage_inst_dmem_ram_4051), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n2001) );
NAND2_X1 MEM_stage_inst_dmem_U2168 ( .A1(MEM_stage_inst_dmem_n1999), .A2(MEM_stage_inst_dmem_n1998), .ZN(MEM_stage_inst_dmem_n2003) );
NAND2_X1 MEM_stage_inst_dmem_U2167 ( .A1(MEM_stage_inst_dmem_ram_4067), .A2(MEM_stage_inst_dmem_n3113), .ZN(MEM_stage_inst_dmem_n1998) );
NAND2_X1 MEM_stage_inst_dmem_U2166 ( .A1(MEM_stage_inst_dmem_ram_3667), .A2(MEM_stage_inst_dmem_n3140), .ZN(MEM_stage_inst_dmem_n1999) );
NOR2_X1 MEM_stage_inst_dmem_U2165 ( .A1(MEM_stage_inst_dmem_n1997), .A2(MEM_stage_inst_dmem_n1996), .ZN(MEM_stage_inst_dmem_n2005) );
NAND2_X1 MEM_stage_inst_dmem_U2164 ( .A1(MEM_stage_inst_dmem_n1995), .A2(MEM_stage_inst_dmem_n1994), .ZN(MEM_stage_inst_dmem_n1996) );
NAND2_X1 MEM_stage_inst_dmem_U2163 ( .A1(MEM_stage_inst_dmem_ram_3971), .A2(MEM_stage_inst_dmem_n3123), .ZN(MEM_stage_inst_dmem_n1994) );
NAND2_X1 MEM_stage_inst_dmem_U2162 ( .A1(MEM_stage_inst_dmem_ram_3651), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n1995) );
NAND2_X1 MEM_stage_inst_dmem_U2161 ( .A1(MEM_stage_inst_dmem_n1993), .A2(MEM_stage_inst_dmem_n1992), .ZN(MEM_stage_inst_dmem_n1997) );
NAND2_X1 MEM_stage_inst_dmem_U2160 ( .A1(MEM_stage_inst_dmem_ram_3923), .A2(MEM_stage_inst_dmem_n3141), .ZN(MEM_stage_inst_dmem_n1992) );
NAND2_X1 MEM_stage_inst_dmem_U2159 ( .A1(MEM_stage_inst_dmem_ram_3491), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n1993) );
NAND2_X1 MEM_stage_inst_dmem_U2158 ( .A1(MEM_stage_inst_dmem_n1991), .A2(MEM_stage_inst_dmem_n1990), .ZN(MEM_stage_inst_dmem_n2007) );
NOR2_X1 MEM_stage_inst_dmem_U2157 ( .A1(MEM_stage_inst_dmem_n1989), .A2(MEM_stage_inst_dmem_n1988), .ZN(MEM_stage_inst_dmem_n1990) );
NAND2_X1 MEM_stage_inst_dmem_U2156 ( .A1(MEM_stage_inst_dmem_n1987), .A2(MEM_stage_inst_dmem_n1986), .ZN(MEM_stage_inst_dmem_n1988) );
NAND2_X1 MEM_stage_inst_dmem_U2155 ( .A1(MEM_stage_inst_dmem_ram_3747), .A2(MEM_stage_inst_dmem_n3155), .ZN(MEM_stage_inst_dmem_n1986) );
NAND2_X1 MEM_stage_inst_dmem_U2154 ( .A1(MEM_stage_inst_dmem_ram_3091), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n1987) );
NAND2_X1 MEM_stage_inst_dmem_U2153 ( .A1(MEM_stage_inst_dmem_n1985), .A2(MEM_stage_inst_dmem_n1984), .ZN(MEM_stage_inst_dmem_n1989) );
NAND2_X1 MEM_stage_inst_dmem_U2152 ( .A1(MEM_stage_inst_dmem_ram_3571), .A2(MEM_stage_inst_dmem_n3170), .ZN(MEM_stage_inst_dmem_n1984) );
NAND2_X1 MEM_stage_inst_dmem_U2151 ( .A1(MEM_stage_inst_dmem_ram_3859), .A2(MEM_stage_inst_dmem_n3191), .ZN(MEM_stage_inst_dmem_n1985) );
NOR2_X1 MEM_stage_inst_dmem_U2150 ( .A1(MEM_stage_inst_dmem_n1983), .A2(MEM_stage_inst_dmem_n1982), .ZN(MEM_stage_inst_dmem_n1991) );
NAND2_X1 MEM_stage_inst_dmem_U2149 ( .A1(MEM_stage_inst_dmem_n1981), .A2(MEM_stage_inst_dmem_n1980), .ZN(MEM_stage_inst_dmem_n1982) );
NAND2_X1 MEM_stage_inst_dmem_U2148 ( .A1(MEM_stage_inst_dmem_ram_3699), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n1980) );
NAND2_X1 MEM_stage_inst_dmem_U2147 ( .A1(MEM_stage_inst_dmem_ram_3603), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n1981) );
NAND2_X1 MEM_stage_inst_dmem_U2146 ( .A1(MEM_stage_inst_dmem_n1979), .A2(MEM_stage_inst_dmem_n1978), .ZN(MEM_stage_inst_dmem_n1983) );
NAND2_X1 MEM_stage_inst_dmem_U2145 ( .A1(MEM_stage_inst_dmem_ram_3187), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n1978) );
NAND2_X1 MEM_stage_inst_dmem_U2144 ( .A1(MEM_stage_inst_dmem_ram_4003), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n1979) );
NAND2_X1 MEM_stage_inst_dmem_U2143 ( .A1(MEM_stage_inst_dmem_n1977), .A2(MEM_stage_inst_dmem_n1976), .ZN(MEM_stage_inst_dmem_n2041) );
NOR2_X1 MEM_stage_inst_dmem_U2142 ( .A1(MEM_stage_inst_dmem_n1975), .A2(MEM_stage_inst_dmem_n1974), .ZN(MEM_stage_inst_dmem_n1976) );
NAND2_X1 MEM_stage_inst_dmem_U2141 ( .A1(MEM_stage_inst_dmem_n1973), .A2(MEM_stage_inst_dmem_n1972), .ZN(MEM_stage_inst_dmem_n1974) );
NOR2_X1 MEM_stage_inst_dmem_U2140 ( .A1(MEM_stage_inst_dmem_n1971), .A2(MEM_stage_inst_dmem_n1970), .ZN(MEM_stage_inst_dmem_n1972) );
NAND2_X1 MEM_stage_inst_dmem_U2139 ( .A1(MEM_stage_inst_dmem_n1969), .A2(MEM_stage_inst_dmem_n1968), .ZN(MEM_stage_inst_dmem_n1970) );
NAND2_X1 MEM_stage_inst_dmem_U2138 ( .A1(MEM_stage_inst_dmem_ram_3907), .A2(MEM_stage_inst_dmem_n3120), .ZN(MEM_stage_inst_dmem_n1968) );
NAND2_X1 MEM_stage_inst_dmem_U2137 ( .A1(MEM_stage_inst_dmem_ram_3795), .A2(MEM_stage_inst_dmem_n3112), .ZN(MEM_stage_inst_dmem_n1969) );
NAND2_X1 MEM_stage_inst_dmem_U2136 ( .A1(MEM_stage_inst_dmem_n1967), .A2(MEM_stage_inst_dmem_n1966), .ZN(MEM_stage_inst_dmem_n1971) );
NAND2_X1 MEM_stage_inst_dmem_U2135 ( .A1(MEM_stage_inst_dmem_ram_3395), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n1966) );
NAND2_X1 MEM_stage_inst_dmem_U2134 ( .A1(MEM_stage_inst_dmem_ram_3123), .A2(MEM_stage_inst_dmem_n3103), .ZN(MEM_stage_inst_dmem_n1967) );
NOR2_X1 MEM_stage_inst_dmem_U2133 ( .A1(MEM_stage_inst_dmem_n1965), .A2(MEM_stage_inst_dmem_n1964), .ZN(MEM_stage_inst_dmem_n1973) );
NAND2_X1 MEM_stage_inst_dmem_U2132 ( .A1(MEM_stage_inst_dmem_n1963), .A2(MEM_stage_inst_dmem_n1962), .ZN(MEM_stage_inst_dmem_n1964) );
NAND2_X1 MEM_stage_inst_dmem_U2131 ( .A1(MEM_stage_inst_dmem_ram_3411), .A2(MEM_stage_inst_dmem_n3216), .ZN(MEM_stage_inst_dmem_n1962) );
NAND2_X1 MEM_stage_inst_dmem_U2130 ( .A1(MEM_stage_inst_dmem_ram_3731), .A2(MEM_stage_inst_dmem_n3076), .ZN(MEM_stage_inst_dmem_n1963) );
NAND2_X1 MEM_stage_inst_dmem_U2129 ( .A1(MEM_stage_inst_dmem_n1961), .A2(MEM_stage_inst_dmem_n1960), .ZN(MEM_stage_inst_dmem_n1965) );
NAND2_X1 MEM_stage_inst_dmem_U2128 ( .A1(MEM_stage_inst_dmem_ram_3475), .A2(MEM_stage_inst_dmem_n3160), .ZN(MEM_stage_inst_dmem_n1960) );
NAND2_X1 MEM_stage_inst_dmem_U2127 ( .A1(MEM_stage_inst_dmem_ram_3155), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n1961) );
NAND2_X1 MEM_stage_inst_dmem_U2126 ( .A1(MEM_stage_inst_dmem_n1959), .A2(MEM_stage_inst_dmem_n1958), .ZN(MEM_stage_inst_dmem_n1975) );
NOR2_X1 MEM_stage_inst_dmem_U2125 ( .A1(MEM_stage_inst_dmem_n1957), .A2(MEM_stage_inst_dmem_n1956), .ZN(MEM_stage_inst_dmem_n1958) );
NAND2_X1 MEM_stage_inst_dmem_U2124 ( .A1(MEM_stage_inst_dmem_n1955), .A2(MEM_stage_inst_dmem_n1954), .ZN(MEM_stage_inst_dmem_n1956) );
NAND2_X1 MEM_stage_inst_dmem_U2123 ( .A1(MEM_stage_inst_dmem_ram_3779), .A2(MEM_stage_inst_dmem_n3192), .ZN(MEM_stage_inst_dmem_n1954) );
NAND2_X1 MEM_stage_inst_dmem_U2122 ( .A1(MEM_stage_inst_dmem_ram_3363), .A2(MEM_stage_inst_dmem_n3209), .ZN(MEM_stage_inst_dmem_n1955) );
NAND2_X1 MEM_stage_inst_dmem_U2121 ( .A1(MEM_stage_inst_dmem_n1953), .A2(MEM_stage_inst_dmem_n1952), .ZN(MEM_stage_inst_dmem_n1957) );
NAND2_X1 MEM_stage_inst_dmem_U2120 ( .A1(MEM_stage_inst_dmem_ram_4035), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n1952) );
NAND2_X1 MEM_stage_inst_dmem_U2119 ( .A1(MEM_stage_inst_dmem_ram_3587), .A2(MEM_stage_inst_dmem_n3182), .ZN(MEM_stage_inst_dmem_n1953) );
NOR2_X1 MEM_stage_inst_dmem_U2118 ( .A1(MEM_stage_inst_dmem_n1951), .A2(MEM_stage_inst_dmem_n1950), .ZN(MEM_stage_inst_dmem_n1959) );
NAND2_X1 MEM_stage_inst_dmem_U2117 ( .A1(MEM_stage_inst_dmem_n1949), .A2(MEM_stage_inst_dmem_n1948), .ZN(MEM_stage_inst_dmem_n1950) );
NAND2_X1 MEM_stage_inst_dmem_U2116 ( .A1(MEM_stage_inst_dmem_ram_3139), .A2(MEM_stage_inst_dmem_n3102), .ZN(MEM_stage_inst_dmem_n1948) );
NAND2_X1 MEM_stage_inst_dmem_U2115 ( .A1(MEM_stage_inst_dmem_ram_3219), .A2(MEM_stage_inst_dmem_n44), .ZN(MEM_stage_inst_dmem_n1949) );
NAND2_X1 MEM_stage_inst_dmem_U2114 ( .A1(MEM_stage_inst_dmem_n1947), .A2(MEM_stage_inst_dmem_n1946), .ZN(MEM_stage_inst_dmem_n1951) );
NAND2_X1 MEM_stage_inst_dmem_U2113 ( .A1(MEM_stage_inst_dmem_ram_3203), .A2(MEM_stage_inst_dmem_n3130), .ZN(MEM_stage_inst_dmem_n1946) );
NAND2_X1 MEM_stage_inst_dmem_U2112 ( .A1(MEM_stage_inst_dmem_ram_4083), .A2(MEM_stage_inst_dmem_n3199), .ZN(MEM_stage_inst_dmem_n1947) );
NOR2_X1 MEM_stage_inst_dmem_U2111 ( .A1(MEM_stage_inst_dmem_n1945), .A2(MEM_stage_inst_dmem_n1944), .ZN(MEM_stage_inst_dmem_n1977) );
NAND2_X1 MEM_stage_inst_dmem_U2110 ( .A1(MEM_stage_inst_dmem_n1943), .A2(MEM_stage_inst_dmem_n1942), .ZN(MEM_stage_inst_dmem_n1944) );
NOR2_X1 MEM_stage_inst_dmem_U2109 ( .A1(MEM_stage_inst_dmem_n1941), .A2(MEM_stage_inst_dmem_n1940), .ZN(MEM_stage_inst_dmem_n1942) );
NAND2_X1 MEM_stage_inst_dmem_U2108 ( .A1(MEM_stage_inst_dmem_n1939), .A2(MEM_stage_inst_dmem_n1938), .ZN(MEM_stage_inst_dmem_n1940) );
NAND2_X1 MEM_stage_inst_dmem_U2107 ( .A1(MEM_stage_inst_dmem_ram_3299), .A2(MEM_stage_inst_dmem_n3152), .ZN(MEM_stage_inst_dmem_n1938) );
NAND2_X1 MEM_stage_inst_dmem_U2106 ( .A1(MEM_stage_inst_dmem_ram_3443), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n1939) );
NAND2_X1 MEM_stage_inst_dmem_U2105 ( .A1(MEM_stage_inst_dmem_n1937), .A2(MEM_stage_inst_dmem_n1936), .ZN(MEM_stage_inst_dmem_n1941) );
NAND2_X1 MEM_stage_inst_dmem_U2104 ( .A1(MEM_stage_inst_dmem_ram_3715), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n1936) );
NAND2_X1 MEM_stage_inst_dmem_U2103 ( .A1(MEM_stage_inst_dmem_ram_3987), .A2(MEM_stage_inst_dmem_n3073), .ZN(MEM_stage_inst_dmem_n1937) );
NOR2_X1 MEM_stage_inst_dmem_U2102 ( .A1(MEM_stage_inst_dmem_n1935), .A2(MEM_stage_inst_dmem_n1934), .ZN(MEM_stage_inst_dmem_n1943) );
NAND2_X1 MEM_stage_inst_dmem_U2101 ( .A1(MEM_stage_inst_dmem_n1933), .A2(MEM_stage_inst_dmem_n1932), .ZN(MEM_stage_inst_dmem_n1934) );
NAND2_X1 MEM_stage_inst_dmem_U2100 ( .A1(MEM_stage_inst_dmem_ram_3267), .A2(MEM_stage_inst_dmem_n3082), .ZN(MEM_stage_inst_dmem_n1932) );
NAND2_X1 MEM_stage_inst_dmem_U2099 ( .A1(MEM_stage_inst_dmem_ram_3331), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n1933) );
NAND2_X1 MEM_stage_inst_dmem_U2098 ( .A1(MEM_stage_inst_dmem_n1931), .A2(MEM_stage_inst_dmem_n1930), .ZN(MEM_stage_inst_dmem_n1935) );
NAND2_X1 MEM_stage_inst_dmem_U2097 ( .A1(MEM_stage_inst_dmem_ram_3827), .A2(MEM_stage_inst_dmem_n3202), .ZN(MEM_stage_inst_dmem_n1930) );
NAND2_X1 MEM_stage_inst_dmem_U2096 ( .A1(MEM_stage_inst_dmem_ram_3619), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n1931) );
NAND2_X1 MEM_stage_inst_dmem_U2095 ( .A1(MEM_stage_inst_dmem_n1929), .A2(MEM_stage_inst_dmem_n1928), .ZN(MEM_stage_inst_dmem_n1945) );
NOR2_X1 MEM_stage_inst_dmem_U2094 ( .A1(MEM_stage_inst_dmem_n1927), .A2(MEM_stage_inst_dmem_n1926), .ZN(MEM_stage_inst_dmem_n1928) );
NAND2_X1 MEM_stage_inst_dmem_U2093 ( .A1(MEM_stage_inst_dmem_n1925), .A2(MEM_stage_inst_dmem_n1924), .ZN(MEM_stage_inst_dmem_n1926) );
NAND2_X1 MEM_stage_inst_dmem_U2092 ( .A1(MEM_stage_inst_dmem_ram_3843), .A2(MEM_stage_inst_dmem_n37), .ZN(MEM_stage_inst_dmem_n1924) );
NAND2_X1 MEM_stage_inst_dmem_U2091 ( .A1(MEM_stage_inst_dmem_ram_3075), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n1925) );
NAND2_X1 MEM_stage_inst_dmem_U2090 ( .A1(MEM_stage_inst_dmem_n1923), .A2(MEM_stage_inst_dmem_n1922), .ZN(MEM_stage_inst_dmem_n1927) );
NAND2_X1 MEM_stage_inst_dmem_U2089 ( .A1(MEM_stage_inst_dmem_ram_3763), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n1922) );
NAND2_X1 MEM_stage_inst_dmem_U2088 ( .A1(MEM_stage_inst_dmem_ram_3683), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n1923) );
NOR2_X1 MEM_stage_inst_dmem_U2087 ( .A1(MEM_stage_inst_dmem_n1921), .A2(MEM_stage_inst_dmem_n1920), .ZN(MEM_stage_inst_dmem_n1929) );
NAND2_X1 MEM_stage_inst_dmem_U2086 ( .A1(MEM_stage_inst_dmem_n1919), .A2(MEM_stage_inst_dmem_n1918), .ZN(MEM_stage_inst_dmem_n1920) );
NAND2_X1 MEM_stage_inst_dmem_U2085 ( .A1(MEM_stage_inst_dmem_ram_3507), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n1918) );
NAND2_X1 MEM_stage_inst_dmem_U2084 ( .A1(MEM_stage_inst_dmem_ram_3539), .A2(MEM_stage_inst_dmem_n3174), .ZN(MEM_stage_inst_dmem_n1919) );
NAND2_X1 MEM_stage_inst_dmem_U2083 ( .A1(MEM_stage_inst_dmem_n1917), .A2(MEM_stage_inst_dmem_n1916), .ZN(MEM_stage_inst_dmem_n1921) );
NAND2_X1 MEM_stage_inst_dmem_U2082 ( .A1(MEM_stage_inst_dmem_ram_3635), .A2(MEM_stage_inst_dmem_n3085), .ZN(MEM_stage_inst_dmem_n1916) );
NAND2_X1 MEM_stage_inst_dmem_U2081 ( .A1(MEM_stage_inst_dmem_ram_3811), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n1917) );
NOR2_X1 MEM_stage_inst_dmem_U2080 ( .A1(MEM_stage_inst_dmem_n1915), .A2(MEM_stage_inst_dmem_n8152), .ZN(MEM_stage_inst_dmem_n2044) );
NOR2_X1 MEM_stage_inst_dmem_U2079 ( .A1(MEM_stage_inst_dmem_n1914), .A2(MEM_stage_inst_dmem_n1913), .ZN(MEM_stage_inst_dmem_n1915) );
NAND2_X1 MEM_stage_inst_dmem_U2078 ( .A1(MEM_stage_inst_dmem_n1912), .A2(MEM_stage_inst_dmem_n1911), .ZN(MEM_stage_inst_dmem_n1913) );
NOR2_X1 MEM_stage_inst_dmem_U2077 ( .A1(MEM_stage_inst_dmem_n1910), .A2(MEM_stage_inst_dmem_n1909), .ZN(MEM_stage_inst_dmem_n1911) );
NAND2_X1 MEM_stage_inst_dmem_U2076 ( .A1(MEM_stage_inst_dmem_n1908), .A2(MEM_stage_inst_dmem_n1907), .ZN(MEM_stage_inst_dmem_n1909) );
NOR2_X1 MEM_stage_inst_dmem_U2075 ( .A1(MEM_stage_inst_dmem_n1906), .A2(MEM_stage_inst_dmem_n1905), .ZN(MEM_stage_inst_dmem_n1907) );
NAND2_X1 MEM_stage_inst_dmem_U2074 ( .A1(MEM_stage_inst_dmem_n1904), .A2(MEM_stage_inst_dmem_n1903), .ZN(MEM_stage_inst_dmem_n1905) );
NAND2_X1 MEM_stage_inst_dmem_U2073 ( .A1(MEM_stage_inst_dmem_ram_1251), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n1903) );
NAND2_X1 MEM_stage_inst_dmem_U2072 ( .A1(MEM_stage_inst_dmem_ram_1139), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n1904) );
NAND2_X1 MEM_stage_inst_dmem_U2071 ( .A1(MEM_stage_inst_dmem_n1902), .A2(MEM_stage_inst_dmem_n1901), .ZN(MEM_stage_inst_dmem_n1906) );
NAND2_X1 MEM_stage_inst_dmem_U2070 ( .A1(MEM_stage_inst_dmem_ram_1859), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n1901) );
NAND2_X1 MEM_stage_inst_dmem_U2069 ( .A1(MEM_stage_inst_dmem_ram_1411), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n1902) );
NOR2_X1 MEM_stage_inst_dmem_U2068 ( .A1(MEM_stage_inst_dmem_n1900), .A2(MEM_stage_inst_dmem_n1899), .ZN(MEM_stage_inst_dmem_n1908) );
NAND2_X1 MEM_stage_inst_dmem_U2067 ( .A1(MEM_stage_inst_dmem_n1898), .A2(MEM_stage_inst_dmem_n1897), .ZN(MEM_stage_inst_dmem_n1899) );
NAND2_X1 MEM_stage_inst_dmem_U2066 ( .A1(MEM_stage_inst_dmem_ram_1331), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n1897) );
NAND2_X1 MEM_stage_inst_dmem_U2065 ( .A1(MEM_stage_inst_dmem_ram_1107), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n1898) );
NAND2_X1 MEM_stage_inst_dmem_U2064 ( .A1(MEM_stage_inst_dmem_n1896), .A2(MEM_stage_inst_dmem_n1895), .ZN(MEM_stage_inst_dmem_n1900) );
NAND2_X1 MEM_stage_inst_dmem_U2063 ( .A1(MEM_stage_inst_dmem_ram_2035), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n1895) );
NAND2_X1 MEM_stage_inst_dmem_U2062 ( .A1(MEM_stage_inst_dmem_ram_1203), .A2(MEM_stage_inst_dmem_n55), .ZN(MEM_stage_inst_dmem_n1896) );
NAND2_X1 MEM_stage_inst_dmem_U2061 ( .A1(MEM_stage_inst_dmem_n1894), .A2(MEM_stage_inst_dmem_n1893), .ZN(MEM_stage_inst_dmem_n1910) );
NOR2_X1 MEM_stage_inst_dmem_U2060 ( .A1(MEM_stage_inst_dmem_n1892), .A2(MEM_stage_inst_dmem_n1891), .ZN(MEM_stage_inst_dmem_n1893) );
NAND2_X1 MEM_stage_inst_dmem_U2059 ( .A1(MEM_stage_inst_dmem_n1890), .A2(MEM_stage_inst_dmem_n1889), .ZN(MEM_stage_inst_dmem_n1891) );
NAND2_X1 MEM_stage_inst_dmem_U2058 ( .A1(MEM_stage_inst_dmem_ram_1123), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n1889) );
NAND2_X1 MEM_stage_inst_dmem_U2057 ( .A1(MEM_stage_inst_dmem_ram_1763), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n1890) );
NAND2_X1 MEM_stage_inst_dmem_U2056 ( .A1(MEM_stage_inst_dmem_n1888), .A2(MEM_stage_inst_dmem_n1887), .ZN(MEM_stage_inst_dmem_n1892) );
NAND2_X1 MEM_stage_inst_dmem_U2055 ( .A1(MEM_stage_inst_dmem_ram_1379), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n1887) );
NAND2_X1 MEM_stage_inst_dmem_U2054 ( .A1(MEM_stage_inst_dmem_ram_1187), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n1888) );
NOR2_X1 MEM_stage_inst_dmem_U2053 ( .A1(MEM_stage_inst_dmem_n1886), .A2(MEM_stage_inst_dmem_n1885), .ZN(MEM_stage_inst_dmem_n1894) );
NAND2_X1 MEM_stage_inst_dmem_U2052 ( .A1(MEM_stage_inst_dmem_n1884), .A2(MEM_stage_inst_dmem_n1883), .ZN(MEM_stage_inst_dmem_n1885) );
NAND2_X1 MEM_stage_inst_dmem_U2051 ( .A1(MEM_stage_inst_dmem_ram_1155), .A2(MEM_stage_inst_dmem_n61), .ZN(MEM_stage_inst_dmem_n1883) );
NAND2_X1 MEM_stage_inst_dmem_U2050 ( .A1(MEM_stage_inst_dmem_ram_1315), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n1884) );
NAND2_X1 MEM_stage_inst_dmem_U2049 ( .A1(MEM_stage_inst_dmem_n1882), .A2(MEM_stage_inst_dmem_n1881), .ZN(MEM_stage_inst_dmem_n1886) );
NAND2_X1 MEM_stage_inst_dmem_U2048 ( .A1(MEM_stage_inst_dmem_ram_1459), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n1881) );
NAND2_X1 MEM_stage_inst_dmem_U2047 ( .A1(MEM_stage_inst_dmem_ram_1587), .A2(MEM_stage_inst_dmem_n41), .ZN(MEM_stage_inst_dmem_n1882) );
NOR2_X1 MEM_stage_inst_dmem_U2046 ( .A1(MEM_stage_inst_dmem_n1880), .A2(MEM_stage_inst_dmem_n1879), .ZN(MEM_stage_inst_dmem_n1912) );
NAND2_X1 MEM_stage_inst_dmem_U2045 ( .A1(MEM_stage_inst_dmem_n1878), .A2(MEM_stage_inst_dmem_n1877), .ZN(MEM_stage_inst_dmem_n1879) );
NOR2_X1 MEM_stage_inst_dmem_U2044 ( .A1(MEM_stage_inst_dmem_n1876), .A2(MEM_stage_inst_dmem_n1875), .ZN(MEM_stage_inst_dmem_n1877) );
NAND2_X1 MEM_stage_inst_dmem_U2043 ( .A1(MEM_stage_inst_dmem_n1874), .A2(MEM_stage_inst_dmem_n1873), .ZN(MEM_stage_inst_dmem_n1875) );
NAND2_X1 MEM_stage_inst_dmem_U2042 ( .A1(MEM_stage_inst_dmem_ram_1955), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n1873) );
NAND2_X1 MEM_stage_inst_dmem_U2041 ( .A1(MEM_stage_inst_dmem_ram_1811), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n1874) );
NAND2_X1 MEM_stage_inst_dmem_U2040 ( .A1(MEM_stage_inst_dmem_n1872), .A2(MEM_stage_inst_dmem_n1871), .ZN(MEM_stage_inst_dmem_n1876) );
NAND2_X1 MEM_stage_inst_dmem_U2039 ( .A1(MEM_stage_inst_dmem_ram_1507), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n1871) );
NAND2_X1 MEM_stage_inst_dmem_U2038 ( .A1(MEM_stage_inst_dmem_ram_1603), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n1872) );
NOR2_X1 MEM_stage_inst_dmem_U2037 ( .A1(MEM_stage_inst_dmem_n1870), .A2(MEM_stage_inst_dmem_n1869), .ZN(MEM_stage_inst_dmem_n1878) );
NAND2_X1 MEM_stage_inst_dmem_U2036 ( .A1(MEM_stage_inst_dmem_n1868), .A2(MEM_stage_inst_dmem_n1867), .ZN(MEM_stage_inst_dmem_n1869) );
NAND2_X1 MEM_stage_inst_dmem_U2035 ( .A1(MEM_stage_inst_dmem_ram_1875), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n1867) );
NAND2_X1 MEM_stage_inst_dmem_U2034 ( .A1(MEM_stage_inst_dmem_ram_1843), .A2(MEM_stage_inst_dmem_n46), .ZN(MEM_stage_inst_dmem_n1868) );
NAND2_X1 MEM_stage_inst_dmem_U2033 ( .A1(MEM_stage_inst_dmem_n1866), .A2(MEM_stage_inst_dmem_n1865), .ZN(MEM_stage_inst_dmem_n1870) );
NAND2_X1 MEM_stage_inst_dmem_U2032 ( .A1(MEM_stage_inst_dmem_ram_1827), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n1865) );
NAND2_X1 MEM_stage_inst_dmem_U2031 ( .A1(MEM_stage_inst_dmem_ram_1363), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n1866) );
NAND2_X1 MEM_stage_inst_dmem_U2030 ( .A1(MEM_stage_inst_dmem_n1864), .A2(MEM_stage_inst_dmem_n1863), .ZN(MEM_stage_inst_dmem_n1880) );
NOR2_X1 MEM_stage_inst_dmem_U2029 ( .A1(MEM_stage_inst_dmem_n1862), .A2(MEM_stage_inst_dmem_n1861), .ZN(MEM_stage_inst_dmem_n1863) );
NAND2_X1 MEM_stage_inst_dmem_U2028 ( .A1(MEM_stage_inst_dmem_n1860), .A2(MEM_stage_inst_dmem_n1859), .ZN(MEM_stage_inst_dmem_n1861) );
NAND2_X1 MEM_stage_inst_dmem_U2027 ( .A1(MEM_stage_inst_dmem_ram_1443), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n1859) );
NAND2_X1 MEM_stage_inst_dmem_U2026 ( .A1(MEM_stage_inst_dmem_ram_1043), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n1860) );
NAND2_X1 MEM_stage_inst_dmem_U2025 ( .A1(MEM_stage_inst_dmem_n1858), .A2(MEM_stage_inst_dmem_n1857), .ZN(MEM_stage_inst_dmem_n1862) );
NAND2_X1 MEM_stage_inst_dmem_U2024 ( .A1(MEM_stage_inst_dmem_ram_1427), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n1857) );
NAND2_X1 MEM_stage_inst_dmem_U2023 ( .A1(MEM_stage_inst_dmem_ram_2019), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n1858) );
NOR2_X1 MEM_stage_inst_dmem_U2022 ( .A1(MEM_stage_inst_dmem_n1856), .A2(MEM_stage_inst_dmem_n1855), .ZN(MEM_stage_inst_dmem_n1864) );
NAND2_X1 MEM_stage_inst_dmem_U2021 ( .A1(MEM_stage_inst_dmem_n1854), .A2(MEM_stage_inst_dmem_n1853), .ZN(MEM_stage_inst_dmem_n1855) );
NAND2_X1 MEM_stage_inst_dmem_U2020 ( .A1(MEM_stage_inst_dmem_ram_1779), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n1853) );
NAND2_X1 MEM_stage_inst_dmem_U2019 ( .A1(MEM_stage_inst_dmem_ram_1283), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n1854) );
NAND2_X1 MEM_stage_inst_dmem_U2018 ( .A1(MEM_stage_inst_dmem_n1852), .A2(MEM_stage_inst_dmem_n1851), .ZN(MEM_stage_inst_dmem_n1856) );
NAND2_X1 MEM_stage_inst_dmem_U2017 ( .A1(MEM_stage_inst_dmem_ram_1891), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n1851) );
NAND2_X1 MEM_stage_inst_dmem_U2016 ( .A1(MEM_stage_inst_dmem_ram_1923), .A2(MEM_stage_inst_dmem_n72), .ZN(MEM_stage_inst_dmem_n1852) );
NAND2_X1 MEM_stage_inst_dmem_U2015 ( .A1(MEM_stage_inst_dmem_n1850), .A2(MEM_stage_inst_dmem_n1849), .ZN(MEM_stage_inst_dmem_n1914) );
NOR2_X1 MEM_stage_inst_dmem_U2014 ( .A1(MEM_stage_inst_dmem_n1848), .A2(MEM_stage_inst_dmem_n1847), .ZN(MEM_stage_inst_dmem_n1849) );
NAND2_X1 MEM_stage_inst_dmem_U2013 ( .A1(MEM_stage_inst_dmem_n1846), .A2(MEM_stage_inst_dmem_n1845), .ZN(MEM_stage_inst_dmem_n1847) );
NOR2_X1 MEM_stage_inst_dmem_U2012 ( .A1(MEM_stage_inst_dmem_n1844), .A2(MEM_stage_inst_dmem_n1843), .ZN(MEM_stage_inst_dmem_n1845) );
NAND2_X1 MEM_stage_inst_dmem_U2011 ( .A1(MEM_stage_inst_dmem_n1842), .A2(MEM_stage_inst_dmem_n1841), .ZN(MEM_stage_inst_dmem_n1843) );
NAND2_X1 MEM_stage_inst_dmem_U2010 ( .A1(MEM_stage_inst_dmem_ram_1667), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n1841) );
NAND2_X1 MEM_stage_inst_dmem_U2009 ( .A1(MEM_stage_inst_dmem_ram_1539), .A2(MEM_stage_inst_dmem_n71), .ZN(MEM_stage_inst_dmem_n1842) );
NAND2_X1 MEM_stage_inst_dmem_U2008 ( .A1(MEM_stage_inst_dmem_n1840), .A2(MEM_stage_inst_dmem_n1839), .ZN(MEM_stage_inst_dmem_n1844) );
NAND2_X1 MEM_stage_inst_dmem_U2007 ( .A1(MEM_stage_inst_dmem_ram_1731), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n1839) );
NAND2_X1 MEM_stage_inst_dmem_U2006 ( .A1(MEM_stage_inst_dmem_ram_1027), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n1840) );
NOR2_X1 MEM_stage_inst_dmem_U2005 ( .A1(MEM_stage_inst_dmem_n1838), .A2(MEM_stage_inst_dmem_n1837), .ZN(MEM_stage_inst_dmem_n1846) );
NAND2_X1 MEM_stage_inst_dmem_U2004 ( .A1(MEM_stage_inst_dmem_n1836), .A2(MEM_stage_inst_dmem_n1835), .ZN(MEM_stage_inst_dmem_n1837) );
NAND2_X1 MEM_stage_inst_dmem_U2003 ( .A1(MEM_stage_inst_dmem_ram_1987), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n1835) );
NAND2_X1 MEM_stage_inst_dmem_U2002 ( .A1(MEM_stage_inst_dmem_ram_1555), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n1836) );
NAND2_X1 MEM_stage_inst_dmem_U2001 ( .A1(MEM_stage_inst_dmem_n1834), .A2(MEM_stage_inst_dmem_n1833), .ZN(MEM_stage_inst_dmem_n1838) );
NAND2_X1 MEM_stage_inst_dmem_U2000 ( .A1(MEM_stage_inst_dmem_ram_1075), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n1833) );
NAND2_X1 MEM_stage_inst_dmem_U1999 ( .A1(MEM_stage_inst_dmem_ram_1491), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n1834) );
NAND2_X1 MEM_stage_inst_dmem_U1998 ( .A1(MEM_stage_inst_dmem_n1832), .A2(MEM_stage_inst_dmem_n1831), .ZN(MEM_stage_inst_dmem_n1848) );
NOR2_X1 MEM_stage_inst_dmem_U1997 ( .A1(MEM_stage_inst_dmem_n1830), .A2(MEM_stage_inst_dmem_n1829), .ZN(MEM_stage_inst_dmem_n1831) );
NAND2_X1 MEM_stage_inst_dmem_U1996 ( .A1(MEM_stage_inst_dmem_n1828), .A2(MEM_stage_inst_dmem_n1827), .ZN(MEM_stage_inst_dmem_n1829) );
NAND2_X1 MEM_stage_inst_dmem_U1995 ( .A1(MEM_stage_inst_dmem_ram_1219), .A2(MEM_stage_inst_dmem_n36), .ZN(MEM_stage_inst_dmem_n1827) );
NAND2_X1 MEM_stage_inst_dmem_U1994 ( .A1(MEM_stage_inst_dmem_ram_1347), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n1828) );
NAND2_X1 MEM_stage_inst_dmem_U1993 ( .A1(MEM_stage_inst_dmem_n1826), .A2(MEM_stage_inst_dmem_n1825), .ZN(MEM_stage_inst_dmem_n1830) );
NAND2_X1 MEM_stage_inst_dmem_U1992 ( .A1(MEM_stage_inst_dmem_ram_1059), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n1825) );
NAND2_X1 MEM_stage_inst_dmem_U1991 ( .A1(MEM_stage_inst_dmem_ram_1171), .A2(MEM_stage_inst_dmem_n44), .ZN(MEM_stage_inst_dmem_n1826) );
NOR2_X1 MEM_stage_inst_dmem_U1990 ( .A1(MEM_stage_inst_dmem_n1824), .A2(MEM_stage_inst_dmem_n1823), .ZN(MEM_stage_inst_dmem_n1832) );
NAND2_X1 MEM_stage_inst_dmem_U1989 ( .A1(MEM_stage_inst_dmem_n1822), .A2(MEM_stage_inst_dmem_n1821), .ZN(MEM_stage_inst_dmem_n1823) );
NAND2_X1 MEM_stage_inst_dmem_U1988 ( .A1(MEM_stage_inst_dmem_ram_1939), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n1821) );
NAND2_X1 MEM_stage_inst_dmem_U1987 ( .A1(MEM_stage_inst_dmem_ram_1651), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n1822) );
NAND2_X1 MEM_stage_inst_dmem_U1986 ( .A1(MEM_stage_inst_dmem_n1820), .A2(MEM_stage_inst_dmem_n1819), .ZN(MEM_stage_inst_dmem_n1824) );
NAND2_X1 MEM_stage_inst_dmem_U1985 ( .A1(MEM_stage_inst_dmem_ram_1267), .A2(MEM_stage_inst_dmem_n39), .ZN(MEM_stage_inst_dmem_n1819) );
NAND2_X1 MEM_stage_inst_dmem_U1984 ( .A1(MEM_stage_inst_dmem_ram_1747), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n1820) );
NOR2_X1 MEM_stage_inst_dmem_U1983 ( .A1(MEM_stage_inst_dmem_n1818), .A2(MEM_stage_inst_dmem_n1817), .ZN(MEM_stage_inst_dmem_n1850) );
NAND2_X1 MEM_stage_inst_dmem_U1982 ( .A1(MEM_stage_inst_dmem_n1816), .A2(MEM_stage_inst_dmem_n1815), .ZN(MEM_stage_inst_dmem_n1817) );
NOR2_X1 MEM_stage_inst_dmem_U1981 ( .A1(MEM_stage_inst_dmem_n1814), .A2(MEM_stage_inst_dmem_n1813), .ZN(MEM_stage_inst_dmem_n1815) );
NAND2_X1 MEM_stage_inst_dmem_U1980 ( .A1(MEM_stage_inst_dmem_n1812), .A2(MEM_stage_inst_dmem_n1811), .ZN(MEM_stage_inst_dmem_n1813) );
NAND2_X1 MEM_stage_inst_dmem_U1979 ( .A1(MEM_stage_inst_dmem_ram_1907), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n1811) );
NAND2_X1 MEM_stage_inst_dmem_U1978 ( .A1(MEM_stage_inst_dmem_ram_1971), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n1812) );
NAND2_X1 MEM_stage_inst_dmem_U1977 ( .A1(MEM_stage_inst_dmem_n1810), .A2(MEM_stage_inst_dmem_n1809), .ZN(MEM_stage_inst_dmem_n1814) );
NAND2_X1 MEM_stage_inst_dmem_U1976 ( .A1(MEM_stage_inst_dmem_ram_1091), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n1809) );
NAND2_X1 MEM_stage_inst_dmem_U1975 ( .A1(MEM_stage_inst_dmem_ram_1395), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n1810) );
NOR2_X1 MEM_stage_inst_dmem_U1974 ( .A1(MEM_stage_inst_dmem_n1808), .A2(MEM_stage_inst_dmem_n1807), .ZN(MEM_stage_inst_dmem_n1816) );
NAND2_X1 MEM_stage_inst_dmem_U1973 ( .A1(MEM_stage_inst_dmem_n1806), .A2(MEM_stage_inst_dmem_n1805), .ZN(MEM_stage_inst_dmem_n1807) );
NAND2_X1 MEM_stage_inst_dmem_U1972 ( .A1(MEM_stage_inst_dmem_ram_1699), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n1805) );
NAND2_X1 MEM_stage_inst_dmem_U1971 ( .A1(MEM_stage_inst_dmem_ram_1235), .A2(MEM_stage_inst_dmem_n51), .ZN(MEM_stage_inst_dmem_n1806) );
NAND2_X1 MEM_stage_inst_dmem_U1970 ( .A1(MEM_stage_inst_dmem_n1804), .A2(MEM_stage_inst_dmem_n1803), .ZN(MEM_stage_inst_dmem_n1808) );
NAND2_X1 MEM_stage_inst_dmem_U1969 ( .A1(MEM_stage_inst_dmem_ram_1571), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n1803) );
NAND2_X1 MEM_stage_inst_dmem_U1968 ( .A1(MEM_stage_inst_dmem_ram_1635), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n1804) );
NAND2_X1 MEM_stage_inst_dmem_U1967 ( .A1(MEM_stage_inst_dmem_n1802), .A2(MEM_stage_inst_dmem_n1801), .ZN(MEM_stage_inst_dmem_n1818) );
NOR2_X1 MEM_stage_inst_dmem_U1966 ( .A1(MEM_stage_inst_dmem_n1800), .A2(MEM_stage_inst_dmem_n1799), .ZN(MEM_stage_inst_dmem_n1801) );
NAND2_X1 MEM_stage_inst_dmem_U1965 ( .A1(MEM_stage_inst_dmem_n1798), .A2(MEM_stage_inst_dmem_n1797), .ZN(MEM_stage_inst_dmem_n1799) );
NAND2_X1 MEM_stage_inst_dmem_U1964 ( .A1(MEM_stage_inst_dmem_ram_1715), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n1797) );
NAND2_X1 MEM_stage_inst_dmem_U1963 ( .A1(MEM_stage_inst_dmem_ram_1683), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n1798) );
NAND2_X1 MEM_stage_inst_dmem_U1962 ( .A1(MEM_stage_inst_dmem_n1796), .A2(MEM_stage_inst_dmem_n1795), .ZN(MEM_stage_inst_dmem_n1800) );
NAND2_X1 MEM_stage_inst_dmem_U1961 ( .A1(MEM_stage_inst_dmem_ram_2003), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n1795) );
NAND2_X1 MEM_stage_inst_dmem_U1960 ( .A1(MEM_stage_inst_dmem_ram_1619), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n1796) );
NOR2_X1 MEM_stage_inst_dmem_U1959 ( .A1(MEM_stage_inst_dmem_n1794), .A2(MEM_stage_inst_dmem_n1793), .ZN(MEM_stage_inst_dmem_n1802) );
NAND2_X1 MEM_stage_inst_dmem_U1958 ( .A1(MEM_stage_inst_dmem_n1792), .A2(MEM_stage_inst_dmem_n1791), .ZN(MEM_stage_inst_dmem_n1793) );
NAND2_X1 MEM_stage_inst_dmem_U1957 ( .A1(MEM_stage_inst_dmem_ram_1795), .A2(MEM_stage_inst_dmem_n37), .ZN(MEM_stage_inst_dmem_n1791) );
NAND2_X1 MEM_stage_inst_dmem_U1956 ( .A1(MEM_stage_inst_dmem_ram_1523), .A2(MEM_stage_inst_dmem_n8535), .ZN(MEM_stage_inst_dmem_n1792) );
NAND2_X1 MEM_stage_inst_dmem_U1955 ( .A1(MEM_stage_inst_dmem_n1790), .A2(MEM_stage_inst_dmem_n1789), .ZN(MEM_stage_inst_dmem_n1794) );
NAND2_X1 MEM_stage_inst_dmem_U1954 ( .A1(MEM_stage_inst_dmem_ram_1299), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n1789) );
NAND2_X1 MEM_stage_inst_dmem_U1953 ( .A1(MEM_stage_inst_dmem_ram_1475), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n1790) );
NAND2_X1 MEM_stage_inst_dmem_U1952 ( .A1(MEM_stage_inst_dmem_n1788), .A2(MEM_stage_inst_dmem_n1787), .ZN(MEM_stage_inst_mem_read_data_2) );
NOR2_X1 MEM_stage_inst_dmem_U1951 ( .A1(MEM_stage_inst_dmem_n1786), .A2(MEM_stage_inst_dmem_n1785), .ZN(MEM_stage_inst_dmem_n1787) );
NOR2_X1 MEM_stage_inst_dmem_U1950 ( .A1(MEM_stage_inst_dmem_n1784), .A2(MEM_stage_inst_dmem_n8286), .ZN(MEM_stage_inst_dmem_n1785) );
NOR2_X1 MEM_stage_inst_dmem_U1949 ( .A1(MEM_stage_inst_dmem_n1783), .A2(MEM_stage_inst_dmem_n1782), .ZN(MEM_stage_inst_dmem_n1784) );
NAND2_X1 MEM_stage_inst_dmem_U1948 ( .A1(MEM_stage_inst_dmem_n1781), .A2(MEM_stage_inst_dmem_n1780), .ZN(MEM_stage_inst_dmem_n1782) );
NOR2_X1 MEM_stage_inst_dmem_U1947 ( .A1(MEM_stage_inst_dmem_n1779), .A2(MEM_stage_inst_dmem_n1778), .ZN(MEM_stage_inst_dmem_n1780) );
NAND2_X1 MEM_stage_inst_dmem_U1946 ( .A1(MEM_stage_inst_dmem_n1777), .A2(MEM_stage_inst_dmem_n1776), .ZN(MEM_stage_inst_dmem_n1778) );
NOR2_X1 MEM_stage_inst_dmem_U1945 ( .A1(MEM_stage_inst_dmem_n1775), .A2(MEM_stage_inst_dmem_n1774), .ZN(MEM_stage_inst_dmem_n1776) );
NAND2_X1 MEM_stage_inst_dmem_U1944 ( .A1(MEM_stage_inst_dmem_n1773), .A2(MEM_stage_inst_dmem_n1772), .ZN(MEM_stage_inst_dmem_n1774) );
NAND2_X1 MEM_stage_inst_dmem_U1943 ( .A1(MEM_stage_inst_dmem_ram_2354), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n1772) );
NAND2_X1 MEM_stage_inst_dmem_U1942 ( .A1(MEM_stage_inst_dmem_ram_2962), .A2(MEM_stage_inst_dmem_n3073), .ZN(MEM_stage_inst_dmem_n1773) );
NAND2_X1 MEM_stage_inst_dmem_U1941 ( .A1(MEM_stage_inst_dmem_n1771), .A2(MEM_stage_inst_dmem_n1770), .ZN(MEM_stage_inst_dmem_n1775) );
NAND2_X1 MEM_stage_inst_dmem_U1940 ( .A1(MEM_stage_inst_dmem_ram_2402), .A2(MEM_stage_inst_dmem_n3217), .ZN(MEM_stage_inst_dmem_n1770) );
NAND2_X1 MEM_stage_inst_dmem_U1939 ( .A1(MEM_stage_inst_dmem_ram_2674), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n1771) );
NOR2_X1 MEM_stage_inst_dmem_U1938 ( .A1(MEM_stage_inst_dmem_n1769), .A2(MEM_stage_inst_dmem_n1768), .ZN(MEM_stage_inst_dmem_n1777) );
NAND2_X1 MEM_stage_inst_dmem_U1937 ( .A1(MEM_stage_inst_dmem_n1767), .A2(MEM_stage_inst_dmem_n1766), .ZN(MEM_stage_inst_dmem_n1768) );
NAND2_X1 MEM_stage_inst_dmem_U1936 ( .A1(MEM_stage_inst_dmem_ram_2610), .A2(MEM_stage_inst_dmem_n3085), .ZN(MEM_stage_inst_dmem_n1766) );
NAND2_X1 MEM_stage_inst_dmem_U1935 ( .A1(MEM_stage_inst_dmem_ram_2066), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n1767) );
NAND2_X1 MEM_stage_inst_dmem_U1934 ( .A1(MEM_stage_inst_dmem_n1765), .A2(MEM_stage_inst_dmem_n1764), .ZN(MEM_stage_inst_dmem_n1769) );
NAND2_X1 MEM_stage_inst_dmem_U1933 ( .A1(MEM_stage_inst_dmem_ram_2098), .A2(MEM_stage_inst_dmem_n3103), .ZN(MEM_stage_inst_dmem_n1764) );
NAND2_X1 MEM_stage_inst_dmem_U1932 ( .A1(MEM_stage_inst_dmem_ram_2594), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n1765) );
NAND2_X1 MEM_stage_inst_dmem_U1931 ( .A1(MEM_stage_inst_dmem_n1763), .A2(MEM_stage_inst_dmem_n1762), .ZN(MEM_stage_inst_dmem_n1779) );
NOR2_X1 MEM_stage_inst_dmem_U1930 ( .A1(MEM_stage_inst_dmem_n1761), .A2(MEM_stage_inst_dmem_n1760), .ZN(MEM_stage_inst_dmem_n1762) );
NAND2_X1 MEM_stage_inst_dmem_U1929 ( .A1(MEM_stage_inst_dmem_n1759), .A2(MEM_stage_inst_dmem_n1758), .ZN(MEM_stage_inst_dmem_n1760) );
NAND2_X1 MEM_stage_inst_dmem_U1928 ( .A1(MEM_stage_inst_dmem_ram_2514), .A2(MEM_stage_inst_dmem_n3174), .ZN(MEM_stage_inst_dmem_n1758) );
NAND2_X1 MEM_stage_inst_dmem_U1927 ( .A1(MEM_stage_inst_dmem_ram_2770), .A2(MEM_stage_inst_dmem_n3112), .ZN(MEM_stage_inst_dmem_n1759) );
NAND2_X1 MEM_stage_inst_dmem_U1926 ( .A1(MEM_stage_inst_dmem_n1757), .A2(MEM_stage_inst_dmem_n1756), .ZN(MEM_stage_inst_dmem_n1761) );
NAND2_X1 MEM_stage_inst_dmem_U1925 ( .A1(MEM_stage_inst_dmem_ram_2482), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n1756) );
NAND2_X1 MEM_stage_inst_dmem_U1924 ( .A1(MEM_stage_inst_dmem_ram_3058), .A2(MEM_stage_inst_dmem_n3199), .ZN(MEM_stage_inst_dmem_n1757) );
NOR2_X1 MEM_stage_inst_dmem_U1923 ( .A1(MEM_stage_inst_dmem_n1755), .A2(MEM_stage_inst_dmem_n1754), .ZN(MEM_stage_inst_dmem_n1763) );
NAND2_X1 MEM_stage_inst_dmem_U1922 ( .A1(MEM_stage_inst_dmem_n1753), .A2(MEM_stage_inst_dmem_n1752), .ZN(MEM_stage_inst_dmem_n1754) );
NAND2_X1 MEM_stage_inst_dmem_U1921 ( .A1(MEM_stage_inst_dmem_ram_2898), .A2(MEM_stage_inst_dmem_n3141), .ZN(MEM_stage_inst_dmem_n1752) );
NAND2_X1 MEM_stage_inst_dmem_U1920 ( .A1(MEM_stage_inst_dmem_ram_2146), .A2(MEM_stage_inst_dmem_n3179), .ZN(MEM_stage_inst_dmem_n1753) );
NAND2_X1 MEM_stage_inst_dmem_U1919 ( .A1(MEM_stage_inst_dmem_n1751), .A2(MEM_stage_inst_dmem_n1750), .ZN(MEM_stage_inst_dmem_n1755) );
NAND2_X1 MEM_stage_inst_dmem_U1918 ( .A1(MEM_stage_inst_dmem_ram_2802), .A2(MEM_stage_inst_dmem_n3202), .ZN(MEM_stage_inst_dmem_n1750) );
NAND2_X1 MEM_stage_inst_dmem_U1917 ( .A1(MEM_stage_inst_dmem_ram_2338), .A2(MEM_stage_inst_dmem_n3209), .ZN(MEM_stage_inst_dmem_n1751) );
NOR2_X1 MEM_stage_inst_dmem_U1916 ( .A1(MEM_stage_inst_dmem_n1749), .A2(MEM_stage_inst_dmem_n1748), .ZN(MEM_stage_inst_dmem_n1781) );
NAND2_X1 MEM_stage_inst_dmem_U1915 ( .A1(MEM_stage_inst_dmem_n1747), .A2(MEM_stage_inst_dmem_n1746), .ZN(MEM_stage_inst_dmem_n1748) );
NOR2_X1 MEM_stage_inst_dmem_U1914 ( .A1(MEM_stage_inst_dmem_n1745), .A2(MEM_stage_inst_dmem_n1744), .ZN(MEM_stage_inst_dmem_n1746) );
NAND2_X1 MEM_stage_inst_dmem_U1913 ( .A1(MEM_stage_inst_dmem_n1743), .A2(MEM_stage_inst_dmem_n1742), .ZN(MEM_stage_inst_dmem_n1744) );
NAND2_X1 MEM_stage_inst_dmem_U1912 ( .A1(MEM_stage_inst_dmem_ram_2178), .A2(MEM_stage_inst_dmem_n3130), .ZN(MEM_stage_inst_dmem_n1742) );
NAND2_X1 MEM_stage_inst_dmem_U1911 ( .A1(MEM_stage_inst_dmem_ram_2210), .A2(MEM_stage_inst_dmem_n3081), .ZN(MEM_stage_inst_dmem_n1743) );
NAND2_X1 MEM_stage_inst_dmem_U1910 ( .A1(MEM_stage_inst_dmem_n1741), .A2(MEM_stage_inst_dmem_n1740), .ZN(MEM_stage_inst_dmem_n1745) );
NAND2_X1 MEM_stage_inst_dmem_U1909 ( .A1(MEM_stage_inst_dmem_ram_2930), .A2(MEM_stage_inst_dmem_n3099), .ZN(MEM_stage_inst_dmem_n1740) );
NAND2_X1 MEM_stage_inst_dmem_U1908 ( .A1(MEM_stage_inst_dmem_ram_2466), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n1741) );
NOR2_X1 MEM_stage_inst_dmem_U1907 ( .A1(MEM_stage_inst_dmem_n1739), .A2(MEM_stage_inst_dmem_n1738), .ZN(MEM_stage_inst_dmem_n1747) );
NAND2_X1 MEM_stage_inst_dmem_U1906 ( .A1(MEM_stage_inst_dmem_n1737), .A2(MEM_stage_inst_dmem_n1736), .ZN(MEM_stage_inst_dmem_n1738) );
NAND2_X1 MEM_stage_inst_dmem_U1905 ( .A1(MEM_stage_inst_dmem_ram_2754), .A2(MEM_stage_inst_dmem_n3192), .ZN(MEM_stage_inst_dmem_n1736) );
NAND2_X1 MEM_stage_inst_dmem_U1904 ( .A1(MEM_stage_inst_dmem_ram_2786), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n1737) );
NAND2_X1 MEM_stage_inst_dmem_U1903 ( .A1(MEM_stage_inst_dmem_n1735), .A2(MEM_stage_inst_dmem_n1734), .ZN(MEM_stage_inst_dmem_n1739) );
NAND2_X1 MEM_stage_inst_dmem_U1902 ( .A1(MEM_stage_inst_dmem_ram_2866), .A2(MEM_stage_inst_dmem_n8005), .ZN(MEM_stage_inst_dmem_n1734) );
NAND2_X1 MEM_stage_inst_dmem_U1901 ( .A1(MEM_stage_inst_dmem_ram_2658), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n1735) );
NAND2_X1 MEM_stage_inst_dmem_U1900 ( .A1(MEM_stage_inst_dmem_n1733), .A2(MEM_stage_inst_dmem_n1732), .ZN(MEM_stage_inst_dmem_n1749) );
NOR2_X1 MEM_stage_inst_dmem_U1899 ( .A1(MEM_stage_inst_dmem_n1731), .A2(MEM_stage_inst_dmem_n1730), .ZN(MEM_stage_inst_dmem_n1732) );
NAND2_X1 MEM_stage_inst_dmem_U1898 ( .A1(MEM_stage_inst_dmem_n1729), .A2(MEM_stage_inst_dmem_n1728), .ZN(MEM_stage_inst_dmem_n1730) );
NAND2_X1 MEM_stage_inst_dmem_U1897 ( .A1(MEM_stage_inst_dmem_ram_2434), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n1728) );
NAND2_X1 MEM_stage_inst_dmem_U1896 ( .A1(MEM_stage_inst_dmem_ram_2562), .A2(MEM_stage_inst_dmem_n3182), .ZN(MEM_stage_inst_dmem_n1729) );
NAND2_X1 MEM_stage_inst_dmem_U1895 ( .A1(MEM_stage_inst_dmem_n1727), .A2(MEM_stage_inst_dmem_n1726), .ZN(MEM_stage_inst_dmem_n1731) );
NAND2_X1 MEM_stage_inst_dmem_U1894 ( .A1(MEM_stage_inst_dmem_ram_2242), .A2(MEM_stage_inst_dmem_n3082), .ZN(MEM_stage_inst_dmem_n1726) );
NAND2_X1 MEM_stage_inst_dmem_U1893 ( .A1(MEM_stage_inst_dmem_ram_2946), .A2(MEM_stage_inst_dmem_n3123), .ZN(MEM_stage_inst_dmem_n1727) );
NOR2_X1 MEM_stage_inst_dmem_U1892 ( .A1(MEM_stage_inst_dmem_n1725), .A2(MEM_stage_inst_dmem_n1724), .ZN(MEM_stage_inst_dmem_n1733) );
NAND2_X1 MEM_stage_inst_dmem_U1891 ( .A1(MEM_stage_inst_dmem_n1723), .A2(MEM_stage_inst_dmem_n1722), .ZN(MEM_stage_inst_dmem_n1724) );
NAND2_X1 MEM_stage_inst_dmem_U1890 ( .A1(MEM_stage_inst_dmem_ram_3026), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n1722) );
NAND2_X1 MEM_stage_inst_dmem_U1889 ( .A1(MEM_stage_inst_dmem_ram_2386), .A2(MEM_stage_inst_dmem_n3216), .ZN(MEM_stage_inst_dmem_n1723) );
NAND2_X1 MEM_stage_inst_dmem_U1888 ( .A1(MEM_stage_inst_dmem_n1721), .A2(MEM_stage_inst_dmem_n1720), .ZN(MEM_stage_inst_dmem_n1725) );
NAND2_X1 MEM_stage_inst_dmem_U1887 ( .A1(MEM_stage_inst_dmem_ram_2322), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n1720) );
NAND2_X1 MEM_stage_inst_dmem_U1886 ( .A1(MEM_stage_inst_dmem_ram_2706), .A2(MEM_stage_inst_dmem_n3076), .ZN(MEM_stage_inst_dmem_n1721) );
NAND2_X1 MEM_stage_inst_dmem_U1885 ( .A1(MEM_stage_inst_dmem_n1719), .A2(MEM_stage_inst_dmem_n1718), .ZN(MEM_stage_inst_dmem_n1783) );
NOR2_X1 MEM_stage_inst_dmem_U1884 ( .A1(MEM_stage_inst_dmem_n1717), .A2(MEM_stage_inst_dmem_n1716), .ZN(MEM_stage_inst_dmem_n1718) );
NAND2_X1 MEM_stage_inst_dmem_U1883 ( .A1(MEM_stage_inst_dmem_n1715), .A2(MEM_stage_inst_dmem_n1714), .ZN(MEM_stage_inst_dmem_n1716) );
NOR2_X1 MEM_stage_inst_dmem_U1882 ( .A1(MEM_stage_inst_dmem_n1713), .A2(MEM_stage_inst_dmem_n1712), .ZN(MEM_stage_inst_dmem_n1714) );
NAND2_X1 MEM_stage_inst_dmem_U1881 ( .A1(MEM_stage_inst_dmem_n1711), .A2(MEM_stage_inst_dmem_n1710), .ZN(MEM_stage_inst_dmem_n1712) );
NAND2_X1 MEM_stage_inst_dmem_U1880 ( .A1(MEM_stage_inst_dmem_ram_2114), .A2(MEM_stage_inst_dmem_n3102), .ZN(MEM_stage_inst_dmem_n1710) );
NAND2_X1 MEM_stage_inst_dmem_U1879 ( .A1(MEM_stage_inst_dmem_ram_2626), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n1711) );
NAND2_X1 MEM_stage_inst_dmem_U1878 ( .A1(MEM_stage_inst_dmem_n1709), .A2(MEM_stage_inst_dmem_n1708), .ZN(MEM_stage_inst_dmem_n1713) );
NAND2_X1 MEM_stage_inst_dmem_U1877 ( .A1(MEM_stage_inst_dmem_ram_2546), .A2(MEM_stage_inst_dmem_n3170), .ZN(MEM_stage_inst_dmem_n1708) );
NAND2_X1 MEM_stage_inst_dmem_U1876 ( .A1(MEM_stage_inst_dmem_ram_2050), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n1709) );
NOR2_X1 MEM_stage_inst_dmem_U1875 ( .A1(MEM_stage_inst_dmem_n1707), .A2(MEM_stage_inst_dmem_n1706), .ZN(MEM_stage_inst_dmem_n1715) );
NAND2_X1 MEM_stage_inst_dmem_U1874 ( .A1(MEM_stage_inst_dmem_n1705), .A2(MEM_stage_inst_dmem_n1704), .ZN(MEM_stage_inst_dmem_n1706) );
NAND2_X1 MEM_stage_inst_dmem_U1873 ( .A1(MEM_stage_inst_dmem_ram_2530), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n1704) );
NAND2_X1 MEM_stage_inst_dmem_U1872 ( .A1(MEM_stage_inst_dmem_ram_2578), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n1705) );
NAND2_X1 MEM_stage_inst_dmem_U1871 ( .A1(MEM_stage_inst_dmem_n1703), .A2(MEM_stage_inst_dmem_n1702), .ZN(MEM_stage_inst_dmem_n1707) );
NAND2_X1 MEM_stage_inst_dmem_U1870 ( .A1(MEM_stage_inst_dmem_ram_2882), .A2(MEM_stage_inst_dmem_n3120), .ZN(MEM_stage_inst_dmem_n1702) );
NAND2_X1 MEM_stage_inst_dmem_U1869 ( .A1(MEM_stage_inst_dmem_ram_2498), .A2(MEM_stage_inst_dmem_n3173), .ZN(MEM_stage_inst_dmem_n1703) );
NAND2_X1 MEM_stage_inst_dmem_U1868 ( .A1(MEM_stage_inst_dmem_n1701), .A2(MEM_stage_inst_dmem_n1700), .ZN(MEM_stage_inst_dmem_n1717) );
NOR2_X1 MEM_stage_inst_dmem_U1867 ( .A1(MEM_stage_inst_dmem_n1699), .A2(MEM_stage_inst_dmem_n1698), .ZN(MEM_stage_inst_dmem_n1700) );
NAND2_X1 MEM_stage_inst_dmem_U1866 ( .A1(MEM_stage_inst_dmem_n1697), .A2(MEM_stage_inst_dmem_n1696), .ZN(MEM_stage_inst_dmem_n1698) );
NAND2_X1 MEM_stage_inst_dmem_U1865 ( .A1(MEM_stage_inst_dmem_ram_2274), .A2(MEM_stage_inst_dmem_n3152), .ZN(MEM_stage_inst_dmem_n1696) );
NAND2_X1 MEM_stage_inst_dmem_U1864 ( .A1(MEM_stage_inst_dmem_ram_2738), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n1697) );
NAND2_X1 MEM_stage_inst_dmem_U1863 ( .A1(MEM_stage_inst_dmem_n1695), .A2(MEM_stage_inst_dmem_n1694), .ZN(MEM_stage_inst_dmem_n1699) );
NAND2_X1 MEM_stage_inst_dmem_U1862 ( .A1(MEM_stage_inst_dmem_ram_2850), .A2(MEM_stage_inst_dmem_n3137), .ZN(MEM_stage_inst_dmem_n1694) );
NAND2_X1 MEM_stage_inst_dmem_U1861 ( .A1(MEM_stage_inst_dmem_ram_2418), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n1695) );
NOR2_X1 MEM_stage_inst_dmem_U1860 ( .A1(MEM_stage_inst_dmem_n1693), .A2(MEM_stage_inst_dmem_n1692), .ZN(MEM_stage_inst_dmem_n1701) );
NAND2_X1 MEM_stage_inst_dmem_U1859 ( .A1(MEM_stage_inst_dmem_n1691), .A2(MEM_stage_inst_dmem_n1690), .ZN(MEM_stage_inst_dmem_n1692) );
NAND2_X1 MEM_stage_inst_dmem_U1858 ( .A1(MEM_stage_inst_dmem_ram_2370), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n1690) );
NAND2_X1 MEM_stage_inst_dmem_U1857 ( .A1(MEM_stage_inst_dmem_ram_2994), .A2(MEM_stage_inst_dmem_n3163), .ZN(MEM_stage_inst_dmem_n1691) );
NAND2_X1 MEM_stage_inst_dmem_U1856 ( .A1(MEM_stage_inst_dmem_n1689), .A2(MEM_stage_inst_dmem_n1688), .ZN(MEM_stage_inst_dmem_n1693) );
NAND2_X1 MEM_stage_inst_dmem_U1855 ( .A1(MEM_stage_inst_dmem_ram_2818), .A2(MEM_stage_inst_dmem_n37), .ZN(MEM_stage_inst_dmem_n1688) );
NAND2_X1 MEM_stage_inst_dmem_U1854 ( .A1(MEM_stage_inst_dmem_ram_2450), .A2(MEM_stage_inst_dmem_n3160), .ZN(MEM_stage_inst_dmem_n1689) );
NOR2_X1 MEM_stage_inst_dmem_U1853 ( .A1(MEM_stage_inst_dmem_n1687), .A2(MEM_stage_inst_dmem_n1686), .ZN(MEM_stage_inst_dmem_n1719) );
NAND2_X1 MEM_stage_inst_dmem_U1852 ( .A1(MEM_stage_inst_dmem_n1685), .A2(MEM_stage_inst_dmem_n1684), .ZN(MEM_stage_inst_dmem_n1686) );
NOR2_X1 MEM_stage_inst_dmem_U1851 ( .A1(MEM_stage_inst_dmem_n1683), .A2(MEM_stage_inst_dmem_n1682), .ZN(MEM_stage_inst_dmem_n1684) );
NAND2_X1 MEM_stage_inst_dmem_U1850 ( .A1(MEM_stage_inst_dmem_n1681), .A2(MEM_stage_inst_dmem_n1680), .ZN(MEM_stage_inst_dmem_n1682) );
NAND2_X1 MEM_stage_inst_dmem_U1849 ( .A1(MEM_stage_inst_dmem_ram_2258), .A2(MEM_stage_inst_dmem_n3220), .ZN(MEM_stage_inst_dmem_n1680) );
NAND2_X1 MEM_stage_inst_dmem_U1848 ( .A1(MEM_stage_inst_dmem_ram_2834), .A2(MEM_stage_inst_dmem_n3191), .ZN(MEM_stage_inst_dmem_n1681) );
NAND2_X1 MEM_stage_inst_dmem_U1847 ( .A1(MEM_stage_inst_dmem_n1679), .A2(MEM_stage_inst_dmem_n1678), .ZN(MEM_stage_inst_dmem_n1683) );
NAND2_X1 MEM_stage_inst_dmem_U1846 ( .A1(MEM_stage_inst_dmem_ram_2690), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n1678) );
NAND2_X1 MEM_stage_inst_dmem_U1845 ( .A1(MEM_stage_inst_dmem_ram_2306), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n1679) );
NOR2_X1 MEM_stage_inst_dmem_U1844 ( .A1(MEM_stage_inst_dmem_n1677), .A2(MEM_stage_inst_dmem_n1676), .ZN(MEM_stage_inst_dmem_n1685) );
NAND2_X1 MEM_stage_inst_dmem_U1843 ( .A1(MEM_stage_inst_dmem_n1675), .A2(MEM_stage_inst_dmem_n1674), .ZN(MEM_stage_inst_dmem_n1676) );
NAND2_X1 MEM_stage_inst_dmem_U1842 ( .A1(MEM_stage_inst_dmem_ram_2290), .A2(MEM_stage_inst_dmem_n7914), .ZN(MEM_stage_inst_dmem_n1674) );
NAND2_X1 MEM_stage_inst_dmem_U1841 ( .A1(MEM_stage_inst_dmem_ram_2978), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n1675) );
NAND2_X1 MEM_stage_inst_dmem_U1840 ( .A1(MEM_stage_inst_dmem_n1673), .A2(MEM_stage_inst_dmem_n1672), .ZN(MEM_stage_inst_dmem_n1677) );
NAND2_X1 MEM_stage_inst_dmem_U1839 ( .A1(MEM_stage_inst_dmem_ram_2082), .A2(MEM_stage_inst_dmem_n3092), .ZN(MEM_stage_inst_dmem_n1672) );
NAND2_X1 MEM_stage_inst_dmem_U1838 ( .A1(MEM_stage_inst_dmem_ram_2226), .A2(MEM_stage_inst_dmem_n55), .ZN(MEM_stage_inst_dmem_n1673) );
NAND2_X1 MEM_stage_inst_dmem_U1837 ( .A1(MEM_stage_inst_dmem_n1671), .A2(MEM_stage_inst_dmem_n1670), .ZN(MEM_stage_inst_dmem_n1687) );
NOR2_X1 MEM_stage_inst_dmem_U1836 ( .A1(MEM_stage_inst_dmem_n1669), .A2(MEM_stage_inst_dmem_n1668), .ZN(MEM_stage_inst_dmem_n1670) );
NAND2_X1 MEM_stage_inst_dmem_U1835 ( .A1(MEM_stage_inst_dmem_n1667), .A2(MEM_stage_inst_dmem_n1666), .ZN(MEM_stage_inst_dmem_n1668) );
NAND2_X1 MEM_stage_inst_dmem_U1834 ( .A1(MEM_stage_inst_dmem_ram_3042), .A2(MEM_stage_inst_dmem_n3113), .ZN(MEM_stage_inst_dmem_n1666) );
NAND2_X1 MEM_stage_inst_dmem_U1833 ( .A1(MEM_stage_inst_dmem_ram_3010), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n1667) );
NAND2_X1 MEM_stage_inst_dmem_U1832 ( .A1(MEM_stage_inst_dmem_n1665), .A2(MEM_stage_inst_dmem_n1664), .ZN(MEM_stage_inst_dmem_n1669) );
NAND2_X1 MEM_stage_inst_dmem_U1831 ( .A1(MEM_stage_inst_dmem_ram_2914), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n1664) );
NAND2_X1 MEM_stage_inst_dmem_U1830 ( .A1(MEM_stage_inst_dmem_ram_2722), .A2(MEM_stage_inst_dmem_n3155), .ZN(MEM_stage_inst_dmem_n1665) );
NOR2_X1 MEM_stage_inst_dmem_U1829 ( .A1(MEM_stage_inst_dmem_n1663), .A2(MEM_stage_inst_dmem_n1662), .ZN(MEM_stage_inst_dmem_n1671) );
NAND2_X1 MEM_stage_inst_dmem_U1828 ( .A1(MEM_stage_inst_dmem_n1661), .A2(MEM_stage_inst_dmem_n1660), .ZN(MEM_stage_inst_dmem_n1662) );
NAND2_X1 MEM_stage_inst_dmem_U1827 ( .A1(MEM_stage_inst_dmem_ram_2130), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n1660) );
NAND2_X1 MEM_stage_inst_dmem_U1826 ( .A1(MEM_stage_inst_dmem_ram_2194), .A2(MEM_stage_inst_dmem_n5807), .ZN(MEM_stage_inst_dmem_n1661) );
NAND2_X1 MEM_stage_inst_dmem_U1825 ( .A1(MEM_stage_inst_dmem_n1659), .A2(MEM_stage_inst_dmem_n1658), .ZN(MEM_stage_inst_dmem_n1663) );
NAND2_X1 MEM_stage_inst_dmem_U1824 ( .A1(MEM_stage_inst_dmem_ram_2162), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n1658) );
NAND2_X1 MEM_stage_inst_dmem_U1823 ( .A1(MEM_stage_inst_dmem_ram_2642), .A2(MEM_stage_inst_dmem_n3140), .ZN(MEM_stage_inst_dmem_n1659) );
NOR2_X1 MEM_stage_inst_dmem_U1822 ( .A1(MEM_stage_inst_dmem_n1657), .A2(MEM_stage_inst_dmem_n8152), .ZN(MEM_stage_inst_dmem_n1786) );
NOR2_X1 MEM_stage_inst_dmem_U1821 ( .A1(MEM_stage_inst_dmem_n1656), .A2(MEM_stage_inst_dmem_n1655), .ZN(MEM_stage_inst_dmem_n1657) );
NAND2_X1 MEM_stage_inst_dmem_U1820 ( .A1(MEM_stage_inst_dmem_n1654), .A2(MEM_stage_inst_dmem_n1653), .ZN(MEM_stage_inst_dmem_n1655) );
NOR2_X1 MEM_stage_inst_dmem_U1819 ( .A1(MEM_stage_inst_dmem_n1652), .A2(MEM_stage_inst_dmem_n1651), .ZN(MEM_stage_inst_dmem_n1653) );
NAND2_X1 MEM_stage_inst_dmem_U1818 ( .A1(MEM_stage_inst_dmem_n1650), .A2(MEM_stage_inst_dmem_n1649), .ZN(MEM_stage_inst_dmem_n1651) );
NOR2_X1 MEM_stage_inst_dmem_U1817 ( .A1(MEM_stage_inst_dmem_n1648), .A2(MEM_stage_inst_dmem_n1647), .ZN(MEM_stage_inst_dmem_n1649) );
NAND2_X1 MEM_stage_inst_dmem_U1816 ( .A1(MEM_stage_inst_dmem_n1646), .A2(MEM_stage_inst_dmem_n1645), .ZN(MEM_stage_inst_dmem_n1647) );
NAND2_X1 MEM_stage_inst_dmem_U1815 ( .A1(MEM_stage_inst_dmem_ram_1858), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n1645) );
NAND2_X1 MEM_stage_inst_dmem_U1814 ( .A1(MEM_stage_inst_dmem_ram_1090), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n1646) );
NAND2_X1 MEM_stage_inst_dmem_U1813 ( .A1(MEM_stage_inst_dmem_n1644), .A2(MEM_stage_inst_dmem_n1643), .ZN(MEM_stage_inst_dmem_n1648) );
NAND2_X1 MEM_stage_inst_dmem_U1812 ( .A1(MEM_stage_inst_dmem_ram_1410), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n1643) );
NAND2_X1 MEM_stage_inst_dmem_U1811 ( .A1(MEM_stage_inst_dmem_ram_1602), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n1644) );
NOR2_X1 MEM_stage_inst_dmem_U1810 ( .A1(MEM_stage_inst_dmem_n1642), .A2(MEM_stage_inst_dmem_n1641), .ZN(MEM_stage_inst_dmem_n1650) );
NAND2_X1 MEM_stage_inst_dmem_U1809 ( .A1(MEM_stage_inst_dmem_n1640), .A2(MEM_stage_inst_dmem_n1639), .ZN(MEM_stage_inst_dmem_n1641) );
NAND2_X1 MEM_stage_inst_dmem_U1808 ( .A1(MEM_stage_inst_dmem_ram_1426), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n1639) );
NAND2_X1 MEM_stage_inst_dmem_U1807 ( .A1(MEM_stage_inst_dmem_ram_1394), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n1640) );
NAND2_X1 MEM_stage_inst_dmem_U1806 ( .A1(MEM_stage_inst_dmem_n1638), .A2(MEM_stage_inst_dmem_n1637), .ZN(MEM_stage_inst_dmem_n1642) );
NAND2_X1 MEM_stage_inst_dmem_U1805 ( .A1(MEM_stage_inst_dmem_ram_1490), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n1637) );
NAND2_X1 MEM_stage_inst_dmem_U1804 ( .A1(MEM_stage_inst_dmem_ram_1234), .A2(MEM_stage_inst_dmem_n51), .ZN(MEM_stage_inst_dmem_n1638) );
NAND2_X1 MEM_stage_inst_dmem_U1803 ( .A1(MEM_stage_inst_dmem_n1636), .A2(MEM_stage_inst_dmem_n1635), .ZN(MEM_stage_inst_dmem_n1652) );
NOR2_X1 MEM_stage_inst_dmem_U1802 ( .A1(MEM_stage_inst_dmem_n1634), .A2(MEM_stage_inst_dmem_n1633), .ZN(MEM_stage_inst_dmem_n1635) );
NAND2_X1 MEM_stage_inst_dmem_U1801 ( .A1(MEM_stage_inst_dmem_n1632), .A2(MEM_stage_inst_dmem_n1631), .ZN(MEM_stage_inst_dmem_n1633) );
NAND2_X1 MEM_stage_inst_dmem_U1800 ( .A1(MEM_stage_inst_dmem_ram_2034), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n1631) );
NAND2_X1 MEM_stage_inst_dmem_U1799 ( .A1(MEM_stage_inst_dmem_ram_1810), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n1632) );
NAND2_X1 MEM_stage_inst_dmem_U1798 ( .A1(MEM_stage_inst_dmem_n1630), .A2(MEM_stage_inst_dmem_n1629), .ZN(MEM_stage_inst_dmem_n1634) );
NAND2_X1 MEM_stage_inst_dmem_U1797 ( .A1(MEM_stage_inst_dmem_ram_1170), .A2(MEM_stage_inst_dmem_n44), .ZN(MEM_stage_inst_dmem_n1629) );
NAND2_X1 MEM_stage_inst_dmem_U1796 ( .A1(MEM_stage_inst_dmem_ram_1762), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n1630) );
NOR2_X1 MEM_stage_inst_dmem_U1795 ( .A1(MEM_stage_inst_dmem_n1628), .A2(MEM_stage_inst_dmem_n1627), .ZN(MEM_stage_inst_dmem_n1636) );
NAND2_X1 MEM_stage_inst_dmem_U1794 ( .A1(MEM_stage_inst_dmem_n1626), .A2(MEM_stage_inst_dmem_n1625), .ZN(MEM_stage_inst_dmem_n1627) );
NAND2_X1 MEM_stage_inst_dmem_U1793 ( .A1(MEM_stage_inst_dmem_ram_2018), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n1625) );
NAND2_X1 MEM_stage_inst_dmem_U1792 ( .A1(MEM_stage_inst_dmem_ram_1138), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n1626) );
NAND2_X1 MEM_stage_inst_dmem_U1791 ( .A1(MEM_stage_inst_dmem_n1624), .A2(MEM_stage_inst_dmem_n1623), .ZN(MEM_stage_inst_dmem_n1628) );
NAND2_X1 MEM_stage_inst_dmem_U1790 ( .A1(MEM_stage_inst_dmem_ram_1218), .A2(MEM_stage_inst_dmem_n36), .ZN(MEM_stage_inst_dmem_n1623) );
NAND2_X1 MEM_stage_inst_dmem_U1789 ( .A1(MEM_stage_inst_dmem_ram_1986), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n1624) );
NOR2_X1 MEM_stage_inst_dmem_U1788 ( .A1(MEM_stage_inst_dmem_n1622), .A2(MEM_stage_inst_dmem_n1621), .ZN(MEM_stage_inst_dmem_n1654) );
NAND2_X1 MEM_stage_inst_dmem_U1787 ( .A1(MEM_stage_inst_dmem_n1620), .A2(MEM_stage_inst_dmem_n1619), .ZN(MEM_stage_inst_dmem_n1621) );
NOR2_X1 MEM_stage_inst_dmem_U1786 ( .A1(MEM_stage_inst_dmem_n1618), .A2(MEM_stage_inst_dmem_n1617), .ZN(MEM_stage_inst_dmem_n1619) );
NAND2_X1 MEM_stage_inst_dmem_U1785 ( .A1(MEM_stage_inst_dmem_n1616), .A2(MEM_stage_inst_dmem_n1615), .ZN(MEM_stage_inst_dmem_n1617) );
NAND2_X1 MEM_stage_inst_dmem_U1784 ( .A1(MEM_stage_inst_dmem_ram_1666), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n1615) );
NAND2_X1 MEM_stage_inst_dmem_U1783 ( .A1(MEM_stage_inst_dmem_ram_1714), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n1616) );
NAND2_X1 MEM_stage_inst_dmem_U1782 ( .A1(MEM_stage_inst_dmem_n1614), .A2(MEM_stage_inst_dmem_n1613), .ZN(MEM_stage_inst_dmem_n1618) );
NAND2_X1 MEM_stage_inst_dmem_U1781 ( .A1(MEM_stage_inst_dmem_ram_1314), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n1613) );
NAND2_X1 MEM_stage_inst_dmem_U1780 ( .A1(MEM_stage_inst_dmem_ram_1282), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n1614) );
NOR2_X1 MEM_stage_inst_dmem_U1779 ( .A1(MEM_stage_inst_dmem_n1612), .A2(MEM_stage_inst_dmem_n1611), .ZN(MEM_stage_inst_dmem_n1620) );
NAND2_X1 MEM_stage_inst_dmem_U1778 ( .A1(MEM_stage_inst_dmem_n1610), .A2(MEM_stage_inst_dmem_n1609), .ZN(MEM_stage_inst_dmem_n1611) );
NAND2_X1 MEM_stage_inst_dmem_U1777 ( .A1(MEM_stage_inst_dmem_ram_1938), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n1609) );
NAND2_X1 MEM_stage_inst_dmem_U1776 ( .A1(MEM_stage_inst_dmem_ram_1746), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n1610) );
NAND2_X1 MEM_stage_inst_dmem_U1775 ( .A1(MEM_stage_inst_dmem_n1608), .A2(MEM_stage_inst_dmem_n1607), .ZN(MEM_stage_inst_dmem_n1612) );
NAND2_X1 MEM_stage_inst_dmem_U1774 ( .A1(MEM_stage_inst_dmem_ram_1506), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n1607) );
NAND2_X1 MEM_stage_inst_dmem_U1773 ( .A1(MEM_stage_inst_dmem_ram_1970), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n1608) );
NAND2_X1 MEM_stage_inst_dmem_U1772 ( .A1(MEM_stage_inst_dmem_n1606), .A2(MEM_stage_inst_dmem_n1605), .ZN(MEM_stage_inst_dmem_n1622) );
NOR2_X1 MEM_stage_inst_dmem_U1771 ( .A1(MEM_stage_inst_dmem_n1604), .A2(MEM_stage_inst_dmem_n1603), .ZN(MEM_stage_inst_dmem_n1605) );
NAND2_X1 MEM_stage_inst_dmem_U1770 ( .A1(MEM_stage_inst_dmem_n1602), .A2(MEM_stage_inst_dmem_n1601), .ZN(MEM_stage_inst_dmem_n1603) );
NAND2_X1 MEM_stage_inst_dmem_U1769 ( .A1(MEM_stage_inst_dmem_ram_1874), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n1601) );
NAND2_X1 MEM_stage_inst_dmem_U1768 ( .A1(MEM_stage_inst_dmem_ram_1250), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n1602) );
NAND2_X1 MEM_stage_inst_dmem_U1767 ( .A1(MEM_stage_inst_dmem_n1600), .A2(MEM_stage_inst_dmem_n1599), .ZN(MEM_stage_inst_dmem_n1604) );
NAND2_X1 MEM_stage_inst_dmem_U1766 ( .A1(MEM_stage_inst_dmem_ram_1890), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n1599) );
NAND2_X1 MEM_stage_inst_dmem_U1765 ( .A1(MEM_stage_inst_dmem_ram_1794), .A2(MEM_stage_inst_dmem_n8472), .ZN(MEM_stage_inst_dmem_n1600) );
NOR2_X1 MEM_stage_inst_dmem_U1764 ( .A1(MEM_stage_inst_dmem_n1598), .A2(MEM_stage_inst_dmem_n1597), .ZN(MEM_stage_inst_dmem_n1606) );
NAND2_X1 MEM_stage_inst_dmem_U1763 ( .A1(MEM_stage_inst_dmem_n1596), .A2(MEM_stage_inst_dmem_n1595), .ZN(MEM_stage_inst_dmem_n1597) );
NAND2_X1 MEM_stage_inst_dmem_U1762 ( .A1(MEM_stage_inst_dmem_ram_1922), .A2(MEM_stage_inst_dmem_n72), .ZN(MEM_stage_inst_dmem_n1595) );
NAND2_X1 MEM_stage_inst_dmem_U1761 ( .A1(MEM_stage_inst_dmem_ram_1634), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n1596) );
NAND2_X1 MEM_stage_inst_dmem_U1760 ( .A1(MEM_stage_inst_dmem_n1594), .A2(MEM_stage_inst_dmem_n1593), .ZN(MEM_stage_inst_dmem_n1598) );
NAND2_X1 MEM_stage_inst_dmem_U1759 ( .A1(MEM_stage_inst_dmem_ram_1906), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n1593) );
NAND2_X1 MEM_stage_inst_dmem_U1758 ( .A1(MEM_stage_inst_dmem_ram_1650), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n1594) );
NAND2_X1 MEM_stage_inst_dmem_U1757 ( .A1(MEM_stage_inst_dmem_n1592), .A2(MEM_stage_inst_dmem_n1591), .ZN(MEM_stage_inst_dmem_n1656) );
NOR2_X1 MEM_stage_inst_dmem_U1756 ( .A1(MEM_stage_inst_dmem_n1590), .A2(MEM_stage_inst_dmem_n1589), .ZN(MEM_stage_inst_dmem_n1591) );
NAND2_X1 MEM_stage_inst_dmem_U1755 ( .A1(MEM_stage_inst_dmem_n1588), .A2(MEM_stage_inst_dmem_n1587), .ZN(MEM_stage_inst_dmem_n1589) );
NOR2_X1 MEM_stage_inst_dmem_U1754 ( .A1(MEM_stage_inst_dmem_n1586), .A2(MEM_stage_inst_dmem_n1585), .ZN(MEM_stage_inst_dmem_n1587) );
NAND2_X1 MEM_stage_inst_dmem_U1753 ( .A1(MEM_stage_inst_dmem_n1584), .A2(MEM_stage_inst_dmem_n1583), .ZN(MEM_stage_inst_dmem_n1585) );
NAND2_X1 MEM_stage_inst_dmem_U1752 ( .A1(MEM_stage_inst_dmem_ram_1954), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n1583) );
NAND2_X1 MEM_stage_inst_dmem_U1751 ( .A1(MEM_stage_inst_dmem_ram_1554), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n1584) );
NAND2_X1 MEM_stage_inst_dmem_U1750 ( .A1(MEM_stage_inst_dmem_n1582), .A2(MEM_stage_inst_dmem_n1581), .ZN(MEM_stage_inst_dmem_n1586) );
NAND2_X1 MEM_stage_inst_dmem_U1749 ( .A1(MEM_stage_inst_dmem_ram_1362), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n1581) );
NAND2_X1 MEM_stage_inst_dmem_U1748 ( .A1(MEM_stage_inst_dmem_ram_1122), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n1582) );
NOR2_X1 MEM_stage_inst_dmem_U1747 ( .A1(MEM_stage_inst_dmem_n1580), .A2(MEM_stage_inst_dmem_n1579), .ZN(MEM_stage_inst_dmem_n1588) );
NAND2_X1 MEM_stage_inst_dmem_U1746 ( .A1(MEM_stage_inst_dmem_n1578), .A2(MEM_stage_inst_dmem_n1577), .ZN(MEM_stage_inst_dmem_n1579) );
NAND2_X1 MEM_stage_inst_dmem_U1745 ( .A1(MEM_stage_inst_dmem_ram_1298), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n1577) );
NAND2_X1 MEM_stage_inst_dmem_U1744 ( .A1(MEM_stage_inst_dmem_ram_1026), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n1578) );
NAND2_X1 MEM_stage_inst_dmem_U1743 ( .A1(MEM_stage_inst_dmem_n1576), .A2(MEM_stage_inst_dmem_n1575), .ZN(MEM_stage_inst_dmem_n1580) );
NAND2_X1 MEM_stage_inst_dmem_U1742 ( .A1(MEM_stage_inst_dmem_ram_1778), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n1575) );
NAND2_X1 MEM_stage_inst_dmem_U1741 ( .A1(MEM_stage_inst_dmem_ram_1698), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n1576) );
NAND2_X1 MEM_stage_inst_dmem_U1740 ( .A1(MEM_stage_inst_dmem_n1574), .A2(MEM_stage_inst_dmem_n1573), .ZN(MEM_stage_inst_dmem_n1590) );
NOR2_X1 MEM_stage_inst_dmem_U1739 ( .A1(MEM_stage_inst_dmem_n1572), .A2(MEM_stage_inst_dmem_n1571), .ZN(MEM_stage_inst_dmem_n1573) );
NAND2_X1 MEM_stage_inst_dmem_U1738 ( .A1(MEM_stage_inst_dmem_n1570), .A2(MEM_stage_inst_dmem_n1569), .ZN(MEM_stage_inst_dmem_n1571) );
NAND2_X1 MEM_stage_inst_dmem_U1737 ( .A1(MEM_stage_inst_dmem_ram_1042), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n1569) );
NAND2_X1 MEM_stage_inst_dmem_U1736 ( .A1(MEM_stage_inst_dmem_ram_1202), .A2(MEM_stage_inst_dmem_n8434), .ZN(MEM_stage_inst_dmem_n1570) );
NAND2_X1 MEM_stage_inst_dmem_U1735 ( .A1(MEM_stage_inst_dmem_n1568), .A2(MEM_stage_inst_dmem_n1567), .ZN(MEM_stage_inst_dmem_n1572) );
NAND2_X1 MEM_stage_inst_dmem_U1734 ( .A1(MEM_stage_inst_dmem_ram_1522), .A2(MEM_stage_inst_dmem_n8535), .ZN(MEM_stage_inst_dmem_n1567) );
NAND2_X1 MEM_stage_inst_dmem_U1733 ( .A1(MEM_stage_inst_dmem_ram_1570), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n1568) );
NOR2_X1 MEM_stage_inst_dmem_U1732 ( .A1(MEM_stage_inst_dmem_n1566), .A2(MEM_stage_inst_dmem_n1565), .ZN(MEM_stage_inst_dmem_n1574) );
NAND2_X1 MEM_stage_inst_dmem_U1731 ( .A1(MEM_stage_inst_dmem_n1564), .A2(MEM_stage_inst_dmem_n1563), .ZN(MEM_stage_inst_dmem_n1565) );
NAND2_X1 MEM_stage_inst_dmem_U1730 ( .A1(MEM_stage_inst_dmem_ram_1442), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n1563) );
NAND2_X1 MEM_stage_inst_dmem_U1729 ( .A1(MEM_stage_inst_dmem_ram_1842), .A2(MEM_stage_inst_dmem_n46), .ZN(MEM_stage_inst_dmem_n1564) );
NAND2_X1 MEM_stage_inst_dmem_U1728 ( .A1(MEM_stage_inst_dmem_n1562), .A2(MEM_stage_inst_dmem_n1561), .ZN(MEM_stage_inst_dmem_n1566) );
NAND2_X1 MEM_stage_inst_dmem_U1727 ( .A1(MEM_stage_inst_dmem_ram_1058), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n1561) );
NAND2_X1 MEM_stage_inst_dmem_U1726 ( .A1(MEM_stage_inst_dmem_ram_1682), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n1562) );
NOR2_X1 MEM_stage_inst_dmem_U1725 ( .A1(MEM_stage_inst_dmem_n1560), .A2(MEM_stage_inst_dmem_n1559), .ZN(MEM_stage_inst_dmem_n1592) );
NAND2_X1 MEM_stage_inst_dmem_U1724 ( .A1(MEM_stage_inst_dmem_n1558), .A2(MEM_stage_inst_dmem_n1557), .ZN(MEM_stage_inst_dmem_n1559) );
NOR2_X1 MEM_stage_inst_dmem_U1723 ( .A1(MEM_stage_inst_dmem_n1556), .A2(MEM_stage_inst_dmem_n1555), .ZN(MEM_stage_inst_dmem_n1557) );
NAND2_X1 MEM_stage_inst_dmem_U1722 ( .A1(MEM_stage_inst_dmem_n1554), .A2(MEM_stage_inst_dmem_n1553), .ZN(MEM_stage_inst_dmem_n1555) );
NAND2_X1 MEM_stage_inst_dmem_U1721 ( .A1(MEM_stage_inst_dmem_ram_1378), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n1553) );
NAND2_X1 MEM_stage_inst_dmem_U1720 ( .A1(MEM_stage_inst_dmem_ram_1538), .A2(MEM_stage_inst_dmem_n71), .ZN(MEM_stage_inst_dmem_n1554) );
NAND2_X1 MEM_stage_inst_dmem_U1719 ( .A1(MEM_stage_inst_dmem_n1552), .A2(MEM_stage_inst_dmem_n1551), .ZN(MEM_stage_inst_dmem_n1556) );
NAND2_X1 MEM_stage_inst_dmem_U1718 ( .A1(MEM_stage_inst_dmem_ram_1586), .A2(MEM_stage_inst_dmem_n41), .ZN(MEM_stage_inst_dmem_n1551) );
NAND2_X1 MEM_stage_inst_dmem_U1717 ( .A1(MEM_stage_inst_dmem_ram_1618), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n1552) );
NOR2_X1 MEM_stage_inst_dmem_U1716 ( .A1(MEM_stage_inst_dmem_n1550), .A2(MEM_stage_inst_dmem_n1549), .ZN(MEM_stage_inst_dmem_n1558) );
NAND2_X1 MEM_stage_inst_dmem_U1715 ( .A1(MEM_stage_inst_dmem_n1548), .A2(MEM_stage_inst_dmem_n1547), .ZN(MEM_stage_inst_dmem_n1549) );
NAND2_X1 MEM_stage_inst_dmem_U1714 ( .A1(MEM_stage_inst_dmem_ram_1730), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n1547) );
NAND2_X1 MEM_stage_inst_dmem_U1713 ( .A1(MEM_stage_inst_dmem_ram_2002), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n1548) );
NAND2_X1 MEM_stage_inst_dmem_U1712 ( .A1(MEM_stage_inst_dmem_n1546), .A2(MEM_stage_inst_dmem_n1545), .ZN(MEM_stage_inst_dmem_n1550) );
NAND2_X1 MEM_stage_inst_dmem_U1711 ( .A1(MEM_stage_inst_dmem_ram_1346), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n1545) );
NAND2_X1 MEM_stage_inst_dmem_U1710 ( .A1(MEM_stage_inst_dmem_ram_1826), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n1546) );
NAND2_X1 MEM_stage_inst_dmem_U1709 ( .A1(MEM_stage_inst_dmem_n1544), .A2(MEM_stage_inst_dmem_n1543), .ZN(MEM_stage_inst_dmem_n1560) );
NOR2_X1 MEM_stage_inst_dmem_U1708 ( .A1(MEM_stage_inst_dmem_n1542), .A2(MEM_stage_inst_dmem_n1541), .ZN(MEM_stage_inst_dmem_n1543) );
NAND2_X1 MEM_stage_inst_dmem_U1707 ( .A1(MEM_stage_inst_dmem_n1540), .A2(MEM_stage_inst_dmem_n1539), .ZN(MEM_stage_inst_dmem_n1541) );
NAND2_X1 MEM_stage_inst_dmem_U1706 ( .A1(MEM_stage_inst_dmem_ram_1458), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n1539) );
NAND2_X1 MEM_stage_inst_dmem_U1705 ( .A1(MEM_stage_inst_dmem_ram_1106), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n1540) );
NAND2_X1 MEM_stage_inst_dmem_U1704 ( .A1(MEM_stage_inst_dmem_n1538), .A2(MEM_stage_inst_dmem_n1537), .ZN(MEM_stage_inst_dmem_n1542) );
NAND2_X1 MEM_stage_inst_dmem_U1703 ( .A1(MEM_stage_inst_dmem_ram_1074), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n1537) );
NAND2_X1 MEM_stage_inst_dmem_U1702 ( .A1(MEM_stage_inst_dmem_ram_1154), .A2(MEM_stage_inst_dmem_n61), .ZN(MEM_stage_inst_dmem_n1538) );
NOR2_X1 MEM_stage_inst_dmem_U1701 ( .A1(MEM_stage_inst_dmem_n1536), .A2(MEM_stage_inst_dmem_n1535), .ZN(MEM_stage_inst_dmem_n1544) );
NAND2_X1 MEM_stage_inst_dmem_U1700 ( .A1(MEM_stage_inst_dmem_n1534), .A2(MEM_stage_inst_dmem_n1533), .ZN(MEM_stage_inst_dmem_n1535) );
NAND2_X1 MEM_stage_inst_dmem_U1699 ( .A1(MEM_stage_inst_dmem_ram_1330), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n1533) );
NAND2_X1 MEM_stage_inst_dmem_U1698 ( .A1(MEM_stage_inst_dmem_ram_1474), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n1534) );
NAND2_X1 MEM_stage_inst_dmem_U1697 ( .A1(MEM_stage_inst_dmem_n1532), .A2(MEM_stage_inst_dmem_n1531), .ZN(MEM_stage_inst_dmem_n1536) );
NAND2_X1 MEM_stage_inst_dmem_U1696 ( .A1(MEM_stage_inst_dmem_ram_1266), .A2(MEM_stage_inst_dmem_n39), .ZN(MEM_stage_inst_dmem_n1531) );
NAND2_X1 MEM_stage_inst_dmem_U1695 ( .A1(MEM_stage_inst_dmem_ram_1186), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n1532) );
NOR2_X1 MEM_stage_inst_dmem_U1694 ( .A1(MEM_stage_inst_dmem_n1530), .A2(MEM_stage_inst_dmem_n1529), .ZN(MEM_stage_inst_dmem_n1788) );
NOR2_X1 MEM_stage_inst_dmem_U1693 ( .A1(MEM_stage_inst_dmem_n1528), .A2(MEM_stage_inst_dmem_n8417), .ZN(MEM_stage_inst_dmem_n1529) );
NOR2_X1 MEM_stage_inst_dmem_U1692 ( .A1(MEM_stage_inst_dmem_n1527), .A2(MEM_stage_inst_dmem_n1526), .ZN(MEM_stage_inst_dmem_n1528) );
NAND2_X1 MEM_stage_inst_dmem_U1691 ( .A1(MEM_stage_inst_dmem_n1525), .A2(MEM_stage_inst_dmem_n1524), .ZN(MEM_stage_inst_dmem_n1526) );
NOR2_X1 MEM_stage_inst_dmem_U1690 ( .A1(MEM_stage_inst_dmem_n1523), .A2(MEM_stage_inst_dmem_n1522), .ZN(MEM_stage_inst_dmem_n1524) );
NAND2_X1 MEM_stage_inst_dmem_U1689 ( .A1(MEM_stage_inst_dmem_n1521), .A2(MEM_stage_inst_dmem_n1520), .ZN(MEM_stage_inst_dmem_n1522) );
NOR2_X1 MEM_stage_inst_dmem_U1688 ( .A1(MEM_stage_inst_dmem_n1519), .A2(MEM_stage_inst_dmem_n1518), .ZN(MEM_stage_inst_dmem_n1520) );
NAND2_X1 MEM_stage_inst_dmem_U1687 ( .A1(MEM_stage_inst_dmem_n1517), .A2(MEM_stage_inst_dmem_n1516), .ZN(MEM_stage_inst_dmem_n1518) );
NAND2_X1 MEM_stage_inst_dmem_U1686 ( .A1(MEM_stage_inst_dmem_ram_3938), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n1516) );
NAND2_X1 MEM_stage_inst_dmem_U1685 ( .A1(MEM_stage_inst_dmem_ram_3234), .A2(MEM_stage_inst_dmem_n3081), .ZN(MEM_stage_inst_dmem_n1517) );
NAND2_X1 MEM_stage_inst_dmem_U1684 ( .A1(MEM_stage_inst_dmem_n1515), .A2(MEM_stage_inst_dmem_n1514), .ZN(MEM_stage_inst_dmem_n1519) );
NAND2_X1 MEM_stage_inst_dmem_U1683 ( .A1(MEM_stage_inst_dmem_ram_3970), .A2(MEM_stage_inst_dmem_n3123), .ZN(MEM_stage_inst_dmem_n1514) );
NAND2_X1 MEM_stage_inst_dmem_U1682 ( .A1(MEM_stage_inst_dmem_ram_3250), .A2(MEM_stage_inst_dmem_n55), .ZN(MEM_stage_inst_dmem_n1515) );
NOR2_X1 MEM_stage_inst_dmem_U1681 ( .A1(MEM_stage_inst_dmem_n1513), .A2(MEM_stage_inst_dmem_n1512), .ZN(MEM_stage_inst_dmem_n1521) );
NAND2_X1 MEM_stage_inst_dmem_U1680 ( .A1(MEM_stage_inst_dmem_n1511), .A2(MEM_stage_inst_dmem_n1510), .ZN(MEM_stage_inst_dmem_n1512) );
NAND2_X1 MEM_stage_inst_dmem_U1679 ( .A1(MEM_stage_inst_dmem_ram_3122), .A2(MEM_stage_inst_dmem_n3103), .ZN(MEM_stage_inst_dmem_n1510) );
NAND2_X1 MEM_stage_inst_dmem_U1678 ( .A1(MEM_stage_inst_dmem_ram_3074), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n1511) );
NAND2_X1 MEM_stage_inst_dmem_U1677 ( .A1(MEM_stage_inst_dmem_n1509), .A2(MEM_stage_inst_dmem_n1508), .ZN(MEM_stage_inst_dmem_n1513) );
NAND2_X1 MEM_stage_inst_dmem_U1676 ( .A1(MEM_stage_inst_dmem_ram_4082), .A2(MEM_stage_inst_dmem_n3199), .ZN(MEM_stage_inst_dmem_n1508) );
NAND2_X1 MEM_stage_inst_dmem_U1675 ( .A1(MEM_stage_inst_dmem_ram_3650), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n1509) );
NAND2_X1 MEM_stage_inst_dmem_U1674 ( .A1(MEM_stage_inst_dmem_n1507), .A2(MEM_stage_inst_dmem_n1506), .ZN(MEM_stage_inst_dmem_n1523) );
NOR2_X1 MEM_stage_inst_dmem_U1673 ( .A1(MEM_stage_inst_dmem_n1505), .A2(MEM_stage_inst_dmem_n1504), .ZN(MEM_stage_inst_dmem_n1506) );
NAND2_X1 MEM_stage_inst_dmem_U1672 ( .A1(MEM_stage_inst_dmem_n1503), .A2(MEM_stage_inst_dmem_n1502), .ZN(MEM_stage_inst_dmem_n1504) );
NAND2_X1 MEM_stage_inst_dmem_U1671 ( .A1(MEM_stage_inst_dmem_ram_3858), .A2(MEM_stage_inst_dmem_n3191), .ZN(MEM_stage_inst_dmem_n1502) );
NAND2_X1 MEM_stage_inst_dmem_U1670 ( .A1(MEM_stage_inst_dmem_ram_3810), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n1503) );
NAND2_X1 MEM_stage_inst_dmem_U1669 ( .A1(MEM_stage_inst_dmem_n1501), .A2(MEM_stage_inst_dmem_n1500), .ZN(MEM_stage_inst_dmem_n1505) );
NAND2_X1 MEM_stage_inst_dmem_U1668 ( .A1(MEM_stage_inst_dmem_ram_4018), .A2(MEM_stage_inst_dmem_n3163), .ZN(MEM_stage_inst_dmem_n1500) );
NAND2_X1 MEM_stage_inst_dmem_U1667 ( .A1(MEM_stage_inst_dmem_ram_3698), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n1501) );
NOR2_X1 MEM_stage_inst_dmem_U1666 ( .A1(MEM_stage_inst_dmem_n1499), .A2(MEM_stage_inst_dmem_n1498), .ZN(MEM_stage_inst_dmem_n1507) );
NAND2_X1 MEM_stage_inst_dmem_U1665 ( .A1(MEM_stage_inst_dmem_n1497), .A2(MEM_stage_inst_dmem_n1496), .ZN(MEM_stage_inst_dmem_n1498) );
NAND2_X1 MEM_stage_inst_dmem_U1664 ( .A1(MEM_stage_inst_dmem_ram_3394), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n1496) );
NAND2_X1 MEM_stage_inst_dmem_U1663 ( .A1(MEM_stage_inst_dmem_ram_4034), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n1497) );
NAND2_X1 MEM_stage_inst_dmem_U1662 ( .A1(MEM_stage_inst_dmem_n1495), .A2(MEM_stage_inst_dmem_n1494), .ZN(MEM_stage_inst_dmem_n1499) );
NAND2_X1 MEM_stage_inst_dmem_U1661 ( .A1(MEM_stage_inst_dmem_ram_3986), .A2(MEM_stage_inst_dmem_n3073), .ZN(MEM_stage_inst_dmem_n1494) );
NAND2_X1 MEM_stage_inst_dmem_U1660 ( .A1(MEM_stage_inst_dmem_ram_3666), .A2(MEM_stage_inst_dmem_n3140), .ZN(MEM_stage_inst_dmem_n1495) );
NOR2_X1 MEM_stage_inst_dmem_U1659 ( .A1(MEM_stage_inst_dmem_n1493), .A2(MEM_stage_inst_dmem_n1492), .ZN(MEM_stage_inst_dmem_n1525) );
NAND2_X1 MEM_stage_inst_dmem_U1658 ( .A1(MEM_stage_inst_dmem_n1491), .A2(MEM_stage_inst_dmem_n1490), .ZN(MEM_stage_inst_dmem_n1492) );
NOR2_X1 MEM_stage_inst_dmem_U1657 ( .A1(MEM_stage_inst_dmem_n1489), .A2(MEM_stage_inst_dmem_n1488), .ZN(MEM_stage_inst_dmem_n1490) );
NAND2_X1 MEM_stage_inst_dmem_U1656 ( .A1(MEM_stage_inst_dmem_n1487), .A2(MEM_stage_inst_dmem_n1486), .ZN(MEM_stage_inst_dmem_n1488) );
NAND2_X1 MEM_stage_inst_dmem_U1655 ( .A1(MEM_stage_inst_dmem_ram_3106), .A2(MEM_stage_inst_dmem_n3092), .ZN(MEM_stage_inst_dmem_n1486) );
NAND2_X1 MEM_stage_inst_dmem_U1654 ( .A1(MEM_stage_inst_dmem_ram_3218), .A2(MEM_stage_inst_dmem_n44), .ZN(MEM_stage_inst_dmem_n1487) );
NAND2_X1 MEM_stage_inst_dmem_U1653 ( .A1(MEM_stage_inst_dmem_n1485), .A2(MEM_stage_inst_dmem_n1484), .ZN(MEM_stage_inst_dmem_n1489) );
NAND2_X1 MEM_stage_inst_dmem_U1652 ( .A1(MEM_stage_inst_dmem_ram_3314), .A2(MEM_stage_inst_dmem_n39), .ZN(MEM_stage_inst_dmem_n1484) );
NAND2_X1 MEM_stage_inst_dmem_U1651 ( .A1(MEM_stage_inst_dmem_ram_3282), .A2(MEM_stage_inst_dmem_n3220), .ZN(MEM_stage_inst_dmem_n1485) );
NOR2_X1 MEM_stage_inst_dmem_U1650 ( .A1(MEM_stage_inst_dmem_n1483), .A2(MEM_stage_inst_dmem_n1482), .ZN(MEM_stage_inst_dmem_n1491) );
NAND2_X1 MEM_stage_inst_dmem_U1649 ( .A1(MEM_stage_inst_dmem_n1481), .A2(MEM_stage_inst_dmem_n1480), .ZN(MEM_stage_inst_dmem_n1482) );
NAND2_X1 MEM_stage_inst_dmem_U1648 ( .A1(MEM_stage_inst_dmem_ram_3906), .A2(MEM_stage_inst_dmem_n3120), .ZN(MEM_stage_inst_dmem_n1480) );
NAND2_X1 MEM_stage_inst_dmem_U1647 ( .A1(MEM_stage_inst_dmem_ram_3362), .A2(MEM_stage_inst_dmem_n3209), .ZN(MEM_stage_inst_dmem_n1481) );
NAND2_X1 MEM_stage_inst_dmem_U1646 ( .A1(MEM_stage_inst_dmem_n1479), .A2(MEM_stage_inst_dmem_n1478), .ZN(MEM_stage_inst_dmem_n1483) );
NAND2_X1 MEM_stage_inst_dmem_U1645 ( .A1(MEM_stage_inst_dmem_ram_3266), .A2(MEM_stage_inst_dmem_n3082), .ZN(MEM_stage_inst_dmem_n1478) );
NAND2_X1 MEM_stage_inst_dmem_U1644 ( .A1(MEM_stage_inst_dmem_ram_3570), .A2(MEM_stage_inst_dmem_n3170), .ZN(MEM_stage_inst_dmem_n1479) );
NAND2_X1 MEM_stage_inst_dmem_U1643 ( .A1(MEM_stage_inst_dmem_n1477), .A2(MEM_stage_inst_dmem_n1476), .ZN(MEM_stage_inst_dmem_n1493) );
NOR2_X1 MEM_stage_inst_dmem_U1642 ( .A1(MEM_stage_inst_dmem_n1475), .A2(MEM_stage_inst_dmem_n1474), .ZN(MEM_stage_inst_dmem_n1476) );
NAND2_X1 MEM_stage_inst_dmem_U1641 ( .A1(MEM_stage_inst_dmem_n1473), .A2(MEM_stage_inst_dmem_n1472), .ZN(MEM_stage_inst_dmem_n1474) );
NAND2_X1 MEM_stage_inst_dmem_U1640 ( .A1(MEM_stage_inst_dmem_ram_3634), .A2(MEM_stage_inst_dmem_n3085), .ZN(MEM_stage_inst_dmem_n1472) );
NAND2_X1 MEM_stage_inst_dmem_U1639 ( .A1(MEM_stage_inst_dmem_ram_3330), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n1473) );
NAND2_X1 MEM_stage_inst_dmem_U1638 ( .A1(MEM_stage_inst_dmem_n1471), .A2(MEM_stage_inst_dmem_n1470), .ZN(MEM_stage_inst_dmem_n1475) );
NAND2_X1 MEM_stage_inst_dmem_U1637 ( .A1(MEM_stage_inst_dmem_ram_3138), .A2(MEM_stage_inst_dmem_n3102), .ZN(MEM_stage_inst_dmem_n1470) );
NAND2_X1 MEM_stage_inst_dmem_U1636 ( .A1(MEM_stage_inst_dmem_ram_3618), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n1471) );
NOR2_X1 MEM_stage_inst_dmem_U1635 ( .A1(MEM_stage_inst_dmem_n1469), .A2(MEM_stage_inst_dmem_n1468), .ZN(MEM_stage_inst_dmem_n1477) );
NAND2_X1 MEM_stage_inst_dmem_U1634 ( .A1(MEM_stage_inst_dmem_n1467), .A2(MEM_stage_inst_dmem_n1466), .ZN(MEM_stage_inst_dmem_n1468) );
NAND2_X1 MEM_stage_inst_dmem_U1633 ( .A1(MEM_stage_inst_dmem_ram_3954), .A2(MEM_stage_inst_dmem_n3099), .ZN(MEM_stage_inst_dmem_n1466) );
NAND2_X1 MEM_stage_inst_dmem_U1632 ( .A1(MEM_stage_inst_dmem_ram_3922), .A2(MEM_stage_inst_dmem_n3141), .ZN(MEM_stage_inst_dmem_n1467) );
NAND2_X1 MEM_stage_inst_dmem_U1631 ( .A1(MEM_stage_inst_dmem_n1465), .A2(MEM_stage_inst_dmem_n1464), .ZN(MEM_stage_inst_dmem_n1469) );
NAND2_X1 MEM_stage_inst_dmem_U1630 ( .A1(MEM_stage_inst_dmem_ram_3346), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n1464) );
NAND2_X1 MEM_stage_inst_dmem_U1629 ( .A1(MEM_stage_inst_dmem_ram_3090), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n1465) );
NAND2_X1 MEM_stage_inst_dmem_U1628 ( .A1(MEM_stage_inst_dmem_n1463), .A2(MEM_stage_inst_dmem_n1462), .ZN(MEM_stage_inst_dmem_n1527) );
NOR2_X1 MEM_stage_inst_dmem_U1627 ( .A1(MEM_stage_inst_dmem_n1461), .A2(MEM_stage_inst_dmem_n1460), .ZN(MEM_stage_inst_dmem_n1462) );
NAND2_X1 MEM_stage_inst_dmem_U1626 ( .A1(MEM_stage_inst_dmem_n1459), .A2(MEM_stage_inst_dmem_n1458), .ZN(MEM_stage_inst_dmem_n1460) );
NOR2_X1 MEM_stage_inst_dmem_U1625 ( .A1(MEM_stage_inst_dmem_n1457), .A2(MEM_stage_inst_dmem_n1456), .ZN(MEM_stage_inst_dmem_n1458) );
NAND2_X1 MEM_stage_inst_dmem_U1624 ( .A1(MEM_stage_inst_dmem_n1455), .A2(MEM_stage_inst_dmem_n1454), .ZN(MEM_stage_inst_dmem_n1456) );
NAND2_X1 MEM_stage_inst_dmem_U1623 ( .A1(MEM_stage_inst_dmem_ram_3506), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n1454) );
NAND2_X1 MEM_stage_inst_dmem_U1622 ( .A1(MEM_stage_inst_dmem_ram_3490), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n1455) );
NAND2_X1 MEM_stage_inst_dmem_U1621 ( .A1(MEM_stage_inst_dmem_n1453), .A2(MEM_stage_inst_dmem_n1452), .ZN(MEM_stage_inst_dmem_n1457) );
NAND2_X1 MEM_stage_inst_dmem_U1620 ( .A1(MEM_stage_inst_dmem_ram_3826), .A2(MEM_stage_inst_dmem_n3202), .ZN(MEM_stage_inst_dmem_n1452) );
NAND2_X1 MEM_stage_inst_dmem_U1619 ( .A1(MEM_stage_inst_dmem_ram_3170), .A2(MEM_stage_inst_dmem_n3179), .ZN(MEM_stage_inst_dmem_n1453) );
NOR2_X1 MEM_stage_inst_dmem_U1618 ( .A1(MEM_stage_inst_dmem_n1451), .A2(MEM_stage_inst_dmem_n1450), .ZN(MEM_stage_inst_dmem_n1459) );
NAND2_X1 MEM_stage_inst_dmem_U1617 ( .A1(MEM_stage_inst_dmem_n1449), .A2(MEM_stage_inst_dmem_n1448), .ZN(MEM_stage_inst_dmem_n1450) );
NAND2_X1 MEM_stage_inst_dmem_U1616 ( .A1(MEM_stage_inst_dmem_ram_3522), .A2(MEM_stage_inst_dmem_n3173), .ZN(MEM_stage_inst_dmem_n1448) );
NAND2_X1 MEM_stage_inst_dmem_U1615 ( .A1(MEM_stage_inst_dmem_ram_3730), .A2(MEM_stage_inst_dmem_n3076), .ZN(MEM_stage_inst_dmem_n1449) );
NAND2_X1 MEM_stage_inst_dmem_U1614 ( .A1(MEM_stage_inst_dmem_n1447), .A2(MEM_stage_inst_dmem_n1446), .ZN(MEM_stage_inst_dmem_n1451) );
NAND2_X1 MEM_stage_inst_dmem_U1613 ( .A1(MEM_stage_inst_dmem_ram_3842), .A2(MEM_stage_inst_dmem_n37), .ZN(MEM_stage_inst_dmem_n1446) );
NAND2_X1 MEM_stage_inst_dmem_U1612 ( .A1(MEM_stage_inst_dmem_ram_3890), .A2(MEM_stage_inst_dmem_n46), .ZN(MEM_stage_inst_dmem_n1447) );
NAND2_X1 MEM_stage_inst_dmem_U1611 ( .A1(MEM_stage_inst_dmem_n1445), .A2(MEM_stage_inst_dmem_n1444), .ZN(MEM_stage_inst_dmem_n1461) );
NOR2_X1 MEM_stage_inst_dmem_U1610 ( .A1(MEM_stage_inst_dmem_n1443), .A2(MEM_stage_inst_dmem_n1442), .ZN(MEM_stage_inst_dmem_n1444) );
NAND2_X1 MEM_stage_inst_dmem_U1609 ( .A1(MEM_stage_inst_dmem_n1441), .A2(MEM_stage_inst_dmem_n1440), .ZN(MEM_stage_inst_dmem_n1442) );
NAND2_X1 MEM_stage_inst_dmem_U1608 ( .A1(MEM_stage_inst_dmem_ram_3426), .A2(MEM_stage_inst_dmem_n3217), .ZN(MEM_stage_inst_dmem_n1440) );
NAND2_X1 MEM_stage_inst_dmem_U1607 ( .A1(MEM_stage_inst_dmem_ram_3298), .A2(MEM_stage_inst_dmem_n3152), .ZN(MEM_stage_inst_dmem_n1441) );
NAND2_X1 MEM_stage_inst_dmem_U1606 ( .A1(MEM_stage_inst_dmem_n1439), .A2(MEM_stage_inst_dmem_n1438), .ZN(MEM_stage_inst_dmem_n1443) );
NAND2_X1 MEM_stage_inst_dmem_U1605 ( .A1(MEM_stage_inst_dmem_ram_3154), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n1438) );
NAND2_X1 MEM_stage_inst_dmem_U1604 ( .A1(MEM_stage_inst_dmem_ram_3538), .A2(MEM_stage_inst_dmem_n3174), .ZN(MEM_stage_inst_dmem_n1439) );
NOR2_X1 MEM_stage_inst_dmem_U1603 ( .A1(MEM_stage_inst_dmem_n1437), .A2(MEM_stage_inst_dmem_n1436), .ZN(MEM_stage_inst_dmem_n1445) );
NAND2_X1 MEM_stage_inst_dmem_U1602 ( .A1(MEM_stage_inst_dmem_n1435), .A2(MEM_stage_inst_dmem_n1434), .ZN(MEM_stage_inst_dmem_n1436) );
NAND2_X1 MEM_stage_inst_dmem_U1601 ( .A1(MEM_stage_inst_dmem_ram_3458), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n1434) );
NAND2_X1 MEM_stage_inst_dmem_U1600 ( .A1(MEM_stage_inst_dmem_ram_3602), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n1435) );
NAND2_X1 MEM_stage_inst_dmem_U1599 ( .A1(MEM_stage_inst_dmem_n1433), .A2(MEM_stage_inst_dmem_n1432), .ZN(MEM_stage_inst_dmem_n1437) );
NAND2_X1 MEM_stage_inst_dmem_U1598 ( .A1(MEM_stage_inst_dmem_ram_4066), .A2(MEM_stage_inst_dmem_n3113), .ZN(MEM_stage_inst_dmem_n1432) );
NAND2_X1 MEM_stage_inst_dmem_U1597 ( .A1(MEM_stage_inst_dmem_ram_4002), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n1433) );
NOR2_X1 MEM_stage_inst_dmem_U1596 ( .A1(MEM_stage_inst_dmem_n1431), .A2(MEM_stage_inst_dmem_n1430), .ZN(MEM_stage_inst_dmem_n1463) );
NAND2_X1 MEM_stage_inst_dmem_U1595 ( .A1(MEM_stage_inst_dmem_n1429), .A2(MEM_stage_inst_dmem_n1428), .ZN(MEM_stage_inst_dmem_n1430) );
NOR2_X1 MEM_stage_inst_dmem_U1594 ( .A1(MEM_stage_inst_dmem_n1427), .A2(MEM_stage_inst_dmem_n1426), .ZN(MEM_stage_inst_dmem_n1428) );
NAND2_X1 MEM_stage_inst_dmem_U1593 ( .A1(MEM_stage_inst_dmem_n1425), .A2(MEM_stage_inst_dmem_n1424), .ZN(MEM_stage_inst_dmem_n1426) );
NAND2_X1 MEM_stage_inst_dmem_U1592 ( .A1(MEM_stage_inst_dmem_ram_3474), .A2(MEM_stage_inst_dmem_n3160), .ZN(MEM_stage_inst_dmem_n1424) );
NAND2_X1 MEM_stage_inst_dmem_U1591 ( .A1(MEM_stage_inst_dmem_ram_3762), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n1425) );
NAND2_X1 MEM_stage_inst_dmem_U1590 ( .A1(MEM_stage_inst_dmem_n1423), .A2(MEM_stage_inst_dmem_n1422), .ZN(MEM_stage_inst_dmem_n1427) );
NAND2_X1 MEM_stage_inst_dmem_U1589 ( .A1(MEM_stage_inst_dmem_ram_3554), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n1422) );
NAND2_X1 MEM_stage_inst_dmem_U1588 ( .A1(MEM_stage_inst_dmem_ram_3410), .A2(MEM_stage_inst_dmem_n3216), .ZN(MEM_stage_inst_dmem_n1423) );
NOR2_X1 MEM_stage_inst_dmem_U1587 ( .A1(MEM_stage_inst_dmem_n1421), .A2(MEM_stage_inst_dmem_n1420), .ZN(MEM_stage_inst_dmem_n1429) );
NAND2_X1 MEM_stage_inst_dmem_U1586 ( .A1(MEM_stage_inst_dmem_n1419), .A2(MEM_stage_inst_dmem_n1418), .ZN(MEM_stage_inst_dmem_n1420) );
NAND2_X1 MEM_stage_inst_dmem_U1585 ( .A1(MEM_stage_inst_dmem_ram_3778), .A2(MEM_stage_inst_dmem_n3192), .ZN(MEM_stage_inst_dmem_n1418) );
NAND2_X1 MEM_stage_inst_dmem_U1584 ( .A1(MEM_stage_inst_dmem_ram_3794), .A2(MEM_stage_inst_dmem_n3112), .ZN(MEM_stage_inst_dmem_n1419) );
NAND2_X1 MEM_stage_inst_dmem_U1583 ( .A1(MEM_stage_inst_dmem_n1417), .A2(MEM_stage_inst_dmem_n1416), .ZN(MEM_stage_inst_dmem_n1421) );
NAND2_X1 MEM_stage_inst_dmem_U1582 ( .A1(MEM_stage_inst_dmem_ram_3746), .A2(MEM_stage_inst_dmem_n3155), .ZN(MEM_stage_inst_dmem_n1416) );
NAND2_X1 MEM_stage_inst_dmem_U1581 ( .A1(MEM_stage_inst_dmem_ram_3186), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n1417) );
NAND2_X1 MEM_stage_inst_dmem_U1580 ( .A1(MEM_stage_inst_dmem_n1415), .A2(MEM_stage_inst_dmem_n1414), .ZN(MEM_stage_inst_dmem_n1431) );
NOR2_X1 MEM_stage_inst_dmem_U1579 ( .A1(MEM_stage_inst_dmem_n1413), .A2(MEM_stage_inst_dmem_n1412), .ZN(MEM_stage_inst_dmem_n1414) );
NAND2_X1 MEM_stage_inst_dmem_U1578 ( .A1(MEM_stage_inst_dmem_n1411), .A2(MEM_stage_inst_dmem_n1410), .ZN(MEM_stage_inst_dmem_n1412) );
NAND2_X1 MEM_stage_inst_dmem_U1577 ( .A1(MEM_stage_inst_dmem_ram_3378), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n1410) );
NAND2_X1 MEM_stage_inst_dmem_U1576 ( .A1(MEM_stage_inst_dmem_ram_3682), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n1411) );
NAND2_X1 MEM_stage_inst_dmem_U1575 ( .A1(MEM_stage_inst_dmem_n1409), .A2(MEM_stage_inst_dmem_n1408), .ZN(MEM_stage_inst_dmem_n1413) );
NAND2_X1 MEM_stage_inst_dmem_U1574 ( .A1(MEM_stage_inst_dmem_ram_3202), .A2(MEM_stage_inst_dmem_n3130), .ZN(MEM_stage_inst_dmem_n1408) );
NAND2_X1 MEM_stage_inst_dmem_U1573 ( .A1(MEM_stage_inst_dmem_ram_3442), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n1409) );
NOR2_X1 MEM_stage_inst_dmem_U1572 ( .A1(MEM_stage_inst_dmem_n1407), .A2(MEM_stage_inst_dmem_n1406), .ZN(MEM_stage_inst_dmem_n1415) );
NAND2_X1 MEM_stage_inst_dmem_U1571 ( .A1(MEM_stage_inst_dmem_n1405), .A2(MEM_stage_inst_dmem_n1404), .ZN(MEM_stage_inst_dmem_n1406) );
NAND2_X1 MEM_stage_inst_dmem_U1570 ( .A1(MEM_stage_inst_dmem_ram_3714), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n1404) );
NAND2_X1 MEM_stage_inst_dmem_U1569 ( .A1(MEM_stage_inst_dmem_ram_4050), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n1405) );
NAND2_X1 MEM_stage_inst_dmem_U1568 ( .A1(MEM_stage_inst_dmem_n1403), .A2(MEM_stage_inst_dmem_n1402), .ZN(MEM_stage_inst_dmem_n1407) );
NAND2_X1 MEM_stage_inst_dmem_U1567 ( .A1(MEM_stage_inst_dmem_ram_3874), .A2(MEM_stage_inst_dmem_n3137), .ZN(MEM_stage_inst_dmem_n1402) );
NAND2_X1 MEM_stage_inst_dmem_U1566 ( .A1(MEM_stage_inst_dmem_ram_3586), .A2(MEM_stage_inst_dmem_n3182), .ZN(MEM_stage_inst_dmem_n1403) );
NOR2_X1 MEM_stage_inst_dmem_U1565 ( .A1(MEM_stage_inst_dmem_n1401), .A2(MEM_stage_inst_dmem_n8551), .ZN(MEM_stage_inst_dmem_n1530) );
NOR2_X1 MEM_stage_inst_dmem_U1564 ( .A1(MEM_stage_inst_dmem_n1400), .A2(MEM_stage_inst_dmem_n1399), .ZN(MEM_stage_inst_dmem_n1401) );
NAND2_X1 MEM_stage_inst_dmem_U1563 ( .A1(MEM_stage_inst_dmem_n1398), .A2(MEM_stage_inst_dmem_n1397), .ZN(MEM_stage_inst_dmem_n1399) );
NOR2_X1 MEM_stage_inst_dmem_U1562 ( .A1(MEM_stage_inst_dmem_n1396), .A2(MEM_stage_inst_dmem_n1395), .ZN(MEM_stage_inst_dmem_n1397) );
NAND2_X1 MEM_stage_inst_dmem_U1561 ( .A1(MEM_stage_inst_dmem_n1394), .A2(MEM_stage_inst_dmem_n1393), .ZN(MEM_stage_inst_dmem_n1395) );
NOR2_X1 MEM_stage_inst_dmem_U1560 ( .A1(MEM_stage_inst_dmem_n1392), .A2(MEM_stage_inst_dmem_n1391), .ZN(MEM_stage_inst_dmem_n1393) );
NAND2_X1 MEM_stage_inst_dmem_U1559 ( .A1(MEM_stage_inst_dmem_n1390), .A2(MEM_stage_inst_dmem_n1389), .ZN(MEM_stage_inst_dmem_n1391) );
NAND2_X1 MEM_stage_inst_dmem_U1558 ( .A1(MEM_stage_inst_dmem_ram_962), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n1389) );
NAND2_X1 MEM_stage_inst_dmem_U1557 ( .A1(MEM_stage_inst_dmem_ram_370), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n1390) );
NAND2_X1 MEM_stage_inst_dmem_U1556 ( .A1(MEM_stage_inst_dmem_n1388), .A2(MEM_stage_inst_dmem_n1387), .ZN(MEM_stage_inst_dmem_n1392) );
NAND2_X1 MEM_stage_inst_dmem_U1555 ( .A1(MEM_stage_inst_dmem_ram_162), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n1387) );
NAND2_X1 MEM_stage_inst_dmem_U1554 ( .A1(MEM_stage_inst_dmem_ram_2), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n1388) );
NOR2_X1 MEM_stage_inst_dmem_U1553 ( .A1(MEM_stage_inst_dmem_n1386), .A2(MEM_stage_inst_dmem_n1385), .ZN(MEM_stage_inst_dmem_n1394) );
NAND2_X1 MEM_stage_inst_dmem_U1552 ( .A1(MEM_stage_inst_dmem_n1384), .A2(MEM_stage_inst_dmem_n1383), .ZN(MEM_stage_inst_dmem_n1385) );
NAND2_X1 MEM_stage_inst_dmem_U1551 ( .A1(MEM_stage_inst_dmem_ram_482), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n1383) );
NAND2_X1 MEM_stage_inst_dmem_U1550 ( .A1(MEM_stage_inst_dmem_ram_34), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n1384) );
NAND2_X1 MEM_stage_inst_dmem_U1549 ( .A1(MEM_stage_inst_dmem_n1382), .A2(MEM_stage_inst_dmem_n1381), .ZN(MEM_stage_inst_dmem_n1386) );
NAND2_X1 MEM_stage_inst_dmem_U1548 ( .A1(MEM_stage_inst_dmem_ram_818), .A2(MEM_stage_inst_dmem_n8005), .ZN(MEM_stage_inst_dmem_n1381) );
NAND2_X1 MEM_stage_inst_dmem_U1547 ( .A1(MEM_stage_inst_dmem_ram_178), .A2(MEM_stage_inst_dmem_n55), .ZN(MEM_stage_inst_dmem_n1382) );
NAND2_X1 MEM_stage_inst_dmem_U1546 ( .A1(MEM_stage_inst_dmem_n1380), .A2(MEM_stage_inst_dmem_n1379), .ZN(MEM_stage_inst_dmem_n1396) );
NOR2_X1 MEM_stage_inst_dmem_U1545 ( .A1(MEM_stage_inst_dmem_n1378), .A2(MEM_stage_inst_dmem_n1377), .ZN(MEM_stage_inst_dmem_n1379) );
NAND2_X1 MEM_stage_inst_dmem_U1544 ( .A1(MEM_stage_inst_dmem_n1376), .A2(MEM_stage_inst_dmem_n1375), .ZN(MEM_stage_inst_dmem_n1377) );
NAND2_X1 MEM_stage_inst_dmem_U1543 ( .A1(MEM_stage_inst_dmem_ram_114), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n1375) );
NAND2_X1 MEM_stage_inst_dmem_U1542 ( .A1(MEM_stage_inst_dmem_ram_258), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n1376) );
NAND2_X1 MEM_stage_inst_dmem_U1541 ( .A1(MEM_stage_inst_dmem_n1374), .A2(MEM_stage_inst_dmem_n1373), .ZN(MEM_stage_inst_dmem_n1378) );
NAND2_X1 MEM_stage_inst_dmem_U1540 ( .A1(MEM_stage_inst_dmem_ram_850), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n1373) );
NAND2_X1 MEM_stage_inst_dmem_U1539 ( .A1(MEM_stage_inst_dmem_ram_98), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n1374) );
NOR2_X1 MEM_stage_inst_dmem_U1538 ( .A1(MEM_stage_inst_dmem_n1372), .A2(MEM_stage_inst_dmem_n1371), .ZN(MEM_stage_inst_dmem_n1380) );
NAND2_X1 MEM_stage_inst_dmem_U1537 ( .A1(MEM_stage_inst_dmem_n1370), .A2(MEM_stage_inst_dmem_n1369), .ZN(MEM_stage_inst_dmem_n1371) );
NAND2_X1 MEM_stage_inst_dmem_U1536 ( .A1(MEM_stage_inst_dmem_ram_866), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n1369) );
NAND2_X1 MEM_stage_inst_dmem_U1535 ( .A1(MEM_stage_inst_dmem_ram_450), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n1370) );
NAND2_X1 MEM_stage_inst_dmem_U1534 ( .A1(MEM_stage_inst_dmem_n1368), .A2(MEM_stage_inst_dmem_n1367), .ZN(MEM_stage_inst_dmem_n1372) );
NAND2_X1 MEM_stage_inst_dmem_U1533 ( .A1(MEM_stage_inst_dmem_ram_754), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n1367) );
NAND2_X1 MEM_stage_inst_dmem_U1532 ( .A1(MEM_stage_inst_dmem_ram_386), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n1368) );
NOR2_X1 MEM_stage_inst_dmem_U1531 ( .A1(MEM_stage_inst_dmem_n1366), .A2(MEM_stage_inst_dmem_n1365), .ZN(MEM_stage_inst_dmem_n1398) );
NAND2_X1 MEM_stage_inst_dmem_U1530 ( .A1(MEM_stage_inst_dmem_n1364), .A2(MEM_stage_inst_dmem_n1363), .ZN(MEM_stage_inst_dmem_n1365) );
NOR2_X1 MEM_stage_inst_dmem_U1529 ( .A1(MEM_stage_inst_dmem_n1362), .A2(MEM_stage_inst_dmem_n1361), .ZN(MEM_stage_inst_dmem_n1363) );
NAND2_X1 MEM_stage_inst_dmem_U1528 ( .A1(MEM_stage_inst_dmem_n1360), .A2(MEM_stage_inst_dmem_n1359), .ZN(MEM_stage_inst_dmem_n1361) );
NAND2_X1 MEM_stage_inst_dmem_U1527 ( .A1(MEM_stage_inst_dmem_ram_130), .A2(MEM_stage_inst_dmem_n61), .ZN(MEM_stage_inst_dmem_n1359) );
NAND2_X1 MEM_stage_inst_dmem_U1526 ( .A1(MEM_stage_inst_dmem_ram_514), .A2(MEM_stage_inst_dmem_n71), .ZN(MEM_stage_inst_dmem_n1360) );
NAND2_X1 MEM_stage_inst_dmem_U1525 ( .A1(MEM_stage_inst_dmem_n1358), .A2(MEM_stage_inst_dmem_n1357), .ZN(MEM_stage_inst_dmem_n1362) );
NAND2_X1 MEM_stage_inst_dmem_U1524 ( .A1(MEM_stage_inst_dmem_ram_642), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n1357) );
NAND2_X1 MEM_stage_inst_dmem_U1523 ( .A1(MEM_stage_inst_dmem_ram_146), .A2(MEM_stage_inst_dmem_n5807), .ZN(MEM_stage_inst_dmem_n1358) );
NOR2_X1 MEM_stage_inst_dmem_U1522 ( .A1(MEM_stage_inst_dmem_n1356), .A2(MEM_stage_inst_dmem_n1355), .ZN(MEM_stage_inst_dmem_n1364) );
NAND2_X1 MEM_stage_inst_dmem_U1521 ( .A1(MEM_stage_inst_dmem_n1354), .A2(MEM_stage_inst_dmem_n1353), .ZN(MEM_stage_inst_dmem_n1355) );
NAND2_X1 MEM_stage_inst_dmem_U1520 ( .A1(MEM_stage_inst_dmem_ram_402), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n1353) );
NAND2_X1 MEM_stage_inst_dmem_U1519 ( .A1(MEM_stage_inst_dmem_ram_994), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n1354) );
NAND2_X1 MEM_stage_inst_dmem_U1518 ( .A1(MEM_stage_inst_dmem_n1352), .A2(MEM_stage_inst_dmem_n1351), .ZN(MEM_stage_inst_dmem_n1356) );
NAND2_X1 MEM_stage_inst_dmem_U1517 ( .A1(MEM_stage_inst_dmem_ram_306), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n1351) );
NAND2_X1 MEM_stage_inst_dmem_U1516 ( .A1(MEM_stage_inst_dmem_ram_418), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n1352) );
NAND2_X1 MEM_stage_inst_dmem_U1515 ( .A1(MEM_stage_inst_dmem_n1350), .A2(MEM_stage_inst_dmem_n1349), .ZN(MEM_stage_inst_dmem_n1366) );
NOR2_X1 MEM_stage_inst_dmem_U1514 ( .A1(MEM_stage_inst_dmem_n1348), .A2(MEM_stage_inst_dmem_n1347), .ZN(MEM_stage_inst_dmem_n1349) );
NAND2_X1 MEM_stage_inst_dmem_U1513 ( .A1(MEM_stage_inst_dmem_n1346), .A2(MEM_stage_inst_dmem_n1345), .ZN(MEM_stage_inst_dmem_n1347) );
NAND2_X1 MEM_stage_inst_dmem_U1512 ( .A1(MEM_stage_inst_dmem_ram_194), .A2(MEM_stage_inst_dmem_n36), .ZN(MEM_stage_inst_dmem_n1345) );
NAND2_X1 MEM_stage_inst_dmem_U1511 ( .A1(MEM_stage_inst_dmem_ram_978), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n1346) );
NAND2_X1 MEM_stage_inst_dmem_U1510 ( .A1(MEM_stage_inst_dmem_n1344), .A2(MEM_stage_inst_dmem_n1343), .ZN(MEM_stage_inst_dmem_n1348) );
NAND2_X1 MEM_stage_inst_dmem_U1509 ( .A1(MEM_stage_inst_dmem_ram_1010), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n1343) );
NAND2_X1 MEM_stage_inst_dmem_U1508 ( .A1(MEM_stage_inst_dmem_ram_658), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n1344) );
NOR2_X1 MEM_stage_inst_dmem_U1507 ( .A1(MEM_stage_inst_dmem_n1342), .A2(MEM_stage_inst_dmem_n1341), .ZN(MEM_stage_inst_dmem_n1350) );
NAND2_X1 MEM_stage_inst_dmem_U1506 ( .A1(MEM_stage_inst_dmem_n1340), .A2(MEM_stage_inst_dmem_n1339), .ZN(MEM_stage_inst_dmem_n1341) );
NAND2_X1 MEM_stage_inst_dmem_U1505 ( .A1(MEM_stage_inst_dmem_ram_274), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n1339) );
NAND2_X1 MEM_stage_inst_dmem_U1504 ( .A1(MEM_stage_inst_dmem_ram_674), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n1340) );
NAND2_X1 MEM_stage_inst_dmem_U1503 ( .A1(MEM_stage_inst_dmem_n1338), .A2(MEM_stage_inst_dmem_n1337), .ZN(MEM_stage_inst_dmem_n1342) );
NAND2_X1 MEM_stage_inst_dmem_U1502 ( .A1(MEM_stage_inst_dmem_ram_898), .A2(MEM_stage_inst_dmem_n72), .ZN(MEM_stage_inst_dmem_n1337) );
NAND2_X1 MEM_stage_inst_dmem_U1501 ( .A1(MEM_stage_inst_dmem_ram_82), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n1338) );
NAND2_X1 MEM_stage_inst_dmem_U1500 ( .A1(MEM_stage_inst_dmem_n1336), .A2(MEM_stage_inst_dmem_n1335), .ZN(MEM_stage_inst_dmem_n1400) );
NOR2_X1 MEM_stage_inst_dmem_U1499 ( .A1(MEM_stage_inst_dmem_n1334), .A2(MEM_stage_inst_dmem_n1333), .ZN(MEM_stage_inst_dmem_n1335) );
NAND2_X1 MEM_stage_inst_dmem_U1498 ( .A1(MEM_stage_inst_dmem_n1332), .A2(MEM_stage_inst_dmem_n1331), .ZN(MEM_stage_inst_dmem_n1333) );
NOR2_X1 MEM_stage_inst_dmem_U1497 ( .A1(MEM_stage_inst_dmem_n1330), .A2(MEM_stage_inst_dmem_n1329), .ZN(MEM_stage_inst_dmem_n1331) );
NAND2_X1 MEM_stage_inst_dmem_U1496 ( .A1(MEM_stage_inst_dmem_n1328), .A2(MEM_stage_inst_dmem_n1327), .ZN(MEM_stage_inst_dmem_n1329) );
NAND2_X1 MEM_stage_inst_dmem_U1495 ( .A1(MEM_stage_inst_dmem_ram_802), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n1327) );
NAND2_X1 MEM_stage_inst_dmem_U1494 ( .A1(MEM_stage_inst_dmem_ram_338), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n1328) );
NAND2_X1 MEM_stage_inst_dmem_U1493 ( .A1(MEM_stage_inst_dmem_n1326), .A2(MEM_stage_inst_dmem_n1325), .ZN(MEM_stage_inst_dmem_n1330) );
NAND2_X1 MEM_stage_inst_dmem_U1492 ( .A1(MEM_stage_inst_dmem_ram_770), .A2(MEM_stage_inst_dmem_n37), .ZN(MEM_stage_inst_dmem_n1325) );
NAND2_X1 MEM_stage_inst_dmem_U1491 ( .A1(MEM_stage_inst_dmem_ram_546), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n1326) );
NOR2_X1 MEM_stage_inst_dmem_U1490 ( .A1(MEM_stage_inst_dmem_n1324), .A2(MEM_stage_inst_dmem_n1323), .ZN(MEM_stage_inst_dmem_n1332) );
NAND2_X1 MEM_stage_inst_dmem_U1489 ( .A1(MEM_stage_inst_dmem_n1322), .A2(MEM_stage_inst_dmem_n1321), .ZN(MEM_stage_inst_dmem_n1323) );
NAND2_X1 MEM_stage_inst_dmem_U1488 ( .A1(MEM_stage_inst_dmem_ram_354), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n1321) );
NAND2_X1 MEM_stage_inst_dmem_U1487 ( .A1(MEM_stage_inst_dmem_ram_210), .A2(MEM_stage_inst_dmem_n51), .ZN(MEM_stage_inst_dmem_n1322) );
NAND2_X1 MEM_stage_inst_dmem_U1486 ( .A1(MEM_stage_inst_dmem_n1320), .A2(MEM_stage_inst_dmem_n1319), .ZN(MEM_stage_inst_dmem_n1324) );
NAND2_X1 MEM_stage_inst_dmem_U1485 ( .A1(MEM_stage_inst_dmem_ram_562), .A2(MEM_stage_inst_dmem_n41), .ZN(MEM_stage_inst_dmem_n1319) );
NAND2_X1 MEM_stage_inst_dmem_U1484 ( .A1(MEM_stage_inst_dmem_ram_50), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n1320) );
NAND2_X1 MEM_stage_inst_dmem_U1483 ( .A1(MEM_stage_inst_dmem_n1318), .A2(MEM_stage_inst_dmem_n1317), .ZN(MEM_stage_inst_dmem_n1334) );
NOR2_X1 MEM_stage_inst_dmem_U1482 ( .A1(MEM_stage_inst_dmem_n1316), .A2(MEM_stage_inst_dmem_n1315), .ZN(MEM_stage_inst_dmem_n1317) );
NAND2_X1 MEM_stage_inst_dmem_U1481 ( .A1(MEM_stage_inst_dmem_n1314), .A2(MEM_stage_inst_dmem_n1313), .ZN(MEM_stage_inst_dmem_n1315) );
NAND2_X1 MEM_stage_inst_dmem_U1480 ( .A1(MEM_stage_inst_dmem_ram_242), .A2(MEM_stage_inst_dmem_n7914), .ZN(MEM_stage_inst_dmem_n1313) );
NAND2_X1 MEM_stage_inst_dmem_U1479 ( .A1(MEM_stage_inst_dmem_ram_290), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n1314) );
NAND2_X1 MEM_stage_inst_dmem_U1478 ( .A1(MEM_stage_inst_dmem_n1312), .A2(MEM_stage_inst_dmem_n1311), .ZN(MEM_stage_inst_dmem_n1316) );
NAND2_X1 MEM_stage_inst_dmem_U1477 ( .A1(MEM_stage_inst_dmem_ram_594), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n1311) );
NAND2_X1 MEM_stage_inst_dmem_U1476 ( .A1(MEM_stage_inst_dmem_ram_722), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n1312) );
NOR2_X1 MEM_stage_inst_dmem_U1475 ( .A1(MEM_stage_inst_dmem_n1310), .A2(MEM_stage_inst_dmem_n1309), .ZN(MEM_stage_inst_dmem_n1318) );
NAND2_X1 MEM_stage_inst_dmem_U1474 ( .A1(MEM_stage_inst_dmem_n1308), .A2(MEM_stage_inst_dmem_n1307), .ZN(MEM_stage_inst_dmem_n1309) );
NAND2_X1 MEM_stage_inst_dmem_U1473 ( .A1(MEM_stage_inst_dmem_ram_226), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n1307) );
NAND2_X1 MEM_stage_inst_dmem_U1472 ( .A1(MEM_stage_inst_dmem_ram_930), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n1308) );
NAND2_X1 MEM_stage_inst_dmem_U1471 ( .A1(MEM_stage_inst_dmem_n1306), .A2(MEM_stage_inst_dmem_n1305), .ZN(MEM_stage_inst_dmem_n1310) );
NAND2_X1 MEM_stage_inst_dmem_U1470 ( .A1(MEM_stage_inst_dmem_ram_914), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n1305) );
NAND2_X1 MEM_stage_inst_dmem_U1469 ( .A1(MEM_stage_inst_dmem_ram_610), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n1306) );
NOR2_X1 MEM_stage_inst_dmem_U1468 ( .A1(MEM_stage_inst_dmem_n1304), .A2(MEM_stage_inst_dmem_n1303), .ZN(MEM_stage_inst_dmem_n1336) );
NAND2_X1 MEM_stage_inst_dmem_U1467 ( .A1(MEM_stage_inst_dmem_n1302), .A2(MEM_stage_inst_dmem_n1301), .ZN(MEM_stage_inst_dmem_n1303) );
NOR2_X1 MEM_stage_inst_dmem_U1466 ( .A1(MEM_stage_inst_dmem_n1300), .A2(MEM_stage_inst_dmem_n1299), .ZN(MEM_stage_inst_dmem_n1301) );
NAND2_X1 MEM_stage_inst_dmem_U1465 ( .A1(MEM_stage_inst_dmem_n1298), .A2(MEM_stage_inst_dmem_n1297), .ZN(MEM_stage_inst_dmem_n1299) );
NAND2_X1 MEM_stage_inst_dmem_U1464 ( .A1(MEM_stage_inst_dmem_ram_498), .A2(MEM_stage_inst_dmem_n8535), .ZN(MEM_stage_inst_dmem_n1297) );
NAND2_X1 MEM_stage_inst_dmem_U1463 ( .A1(MEM_stage_inst_dmem_ram_66), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n1298) );
NAND2_X1 MEM_stage_inst_dmem_U1462 ( .A1(MEM_stage_inst_dmem_n1296), .A2(MEM_stage_inst_dmem_n1295), .ZN(MEM_stage_inst_dmem_n1300) );
NAND2_X1 MEM_stage_inst_dmem_U1461 ( .A1(MEM_stage_inst_dmem_ram_946), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n1295) );
NAND2_X1 MEM_stage_inst_dmem_U1460 ( .A1(MEM_stage_inst_dmem_ram_626), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n1296) );
NOR2_X1 MEM_stage_inst_dmem_U1459 ( .A1(MEM_stage_inst_dmem_n1294), .A2(MEM_stage_inst_dmem_n1293), .ZN(MEM_stage_inst_dmem_n1302) );
NAND2_X1 MEM_stage_inst_dmem_U1458 ( .A1(MEM_stage_inst_dmem_n1292), .A2(MEM_stage_inst_dmem_n1291), .ZN(MEM_stage_inst_dmem_n1293) );
NAND2_X1 MEM_stage_inst_dmem_U1457 ( .A1(MEM_stage_inst_dmem_ram_466), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n1291) );
NAND2_X1 MEM_stage_inst_dmem_U1456 ( .A1(MEM_stage_inst_dmem_ram_738), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n1292) );
NAND2_X1 MEM_stage_inst_dmem_U1455 ( .A1(MEM_stage_inst_dmem_n1290), .A2(MEM_stage_inst_dmem_n1289), .ZN(MEM_stage_inst_dmem_n1294) );
NAND2_X1 MEM_stage_inst_dmem_U1454 ( .A1(MEM_stage_inst_dmem_ram_882), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n1289) );
NAND2_X1 MEM_stage_inst_dmem_U1453 ( .A1(MEM_stage_inst_dmem_ram_530), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n1290) );
NAND2_X1 MEM_stage_inst_dmem_U1452 ( .A1(MEM_stage_inst_dmem_n1288), .A2(MEM_stage_inst_dmem_n1287), .ZN(MEM_stage_inst_dmem_n1304) );
NOR2_X1 MEM_stage_inst_dmem_U1451 ( .A1(MEM_stage_inst_dmem_n1286), .A2(MEM_stage_inst_dmem_n1285), .ZN(MEM_stage_inst_dmem_n1287) );
NAND2_X1 MEM_stage_inst_dmem_U1450 ( .A1(MEM_stage_inst_dmem_n1284), .A2(MEM_stage_inst_dmem_n1283), .ZN(MEM_stage_inst_dmem_n1285) );
NAND2_X1 MEM_stage_inst_dmem_U1449 ( .A1(MEM_stage_inst_dmem_ram_834), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n1283) );
NAND2_X1 MEM_stage_inst_dmem_U1448 ( .A1(MEM_stage_inst_dmem_ram_18), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n1284) );
NAND2_X1 MEM_stage_inst_dmem_U1447 ( .A1(MEM_stage_inst_dmem_n1282), .A2(MEM_stage_inst_dmem_n1281), .ZN(MEM_stage_inst_dmem_n1286) );
NAND2_X1 MEM_stage_inst_dmem_U1446 ( .A1(MEM_stage_inst_dmem_ram_434), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n1281) );
NAND2_X1 MEM_stage_inst_dmem_U1445 ( .A1(MEM_stage_inst_dmem_ram_690), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n1282) );
NOR2_X1 MEM_stage_inst_dmem_U1444 ( .A1(MEM_stage_inst_dmem_n1280), .A2(MEM_stage_inst_dmem_n1279), .ZN(MEM_stage_inst_dmem_n1288) );
NAND2_X1 MEM_stage_inst_dmem_U1443 ( .A1(MEM_stage_inst_dmem_n1278), .A2(MEM_stage_inst_dmem_n1277), .ZN(MEM_stage_inst_dmem_n1279) );
NAND2_X1 MEM_stage_inst_dmem_U1442 ( .A1(MEM_stage_inst_dmem_ram_322), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n1277) );
NAND2_X1 MEM_stage_inst_dmem_U1441 ( .A1(MEM_stage_inst_dmem_ram_786), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n1278) );
NAND2_X1 MEM_stage_inst_dmem_U1440 ( .A1(MEM_stage_inst_dmem_n1276), .A2(MEM_stage_inst_dmem_n1275), .ZN(MEM_stage_inst_dmem_n1280) );
NAND2_X1 MEM_stage_inst_dmem_U1439 ( .A1(MEM_stage_inst_dmem_ram_706), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n1275) );
NAND2_X1 MEM_stage_inst_dmem_U1438 ( .A1(MEM_stage_inst_dmem_ram_578), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n1276) );
NAND2_X1 MEM_stage_inst_dmem_U1437 ( .A1(MEM_stage_inst_dmem_n1274), .A2(MEM_stage_inst_dmem_n1273), .ZN(MEM_stage_inst_mem_read_data_1) );
NOR2_X1 MEM_stage_inst_dmem_U1436 ( .A1(MEM_stage_inst_dmem_n1272), .A2(MEM_stage_inst_dmem_n1271), .ZN(MEM_stage_inst_dmem_n1273) );
NOR2_X1 MEM_stage_inst_dmem_U1435 ( .A1(MEM_stage_inst_dmem_n1270), .A2(MEM_stage_inst_dmem_n8286), .ZN(MEM_stage_inst_dmem_n1271) );
NOR2_X1 MEM_stage_inst_dmem_U1434 ( .A1(MEM_stage_inst_dmem_n1269), .A2(MEM_stage_inst_dmem_n1268), .ZN(MEM_stage_inst_dmem_n1270) );
NAND2_X1 MEM_stage_inst_dmem_U1433 ( .A1(MEM_stage_inst_dmem_n1267), .A2(MEM_stage_inst_dmem_n1266), .ZN(MEM_stage_inst_dmem_n1268) );
NOR2_X1 MEM_stage_inst_dmem_U1432 ( .A1(MEM_stage_inst_dmem_n1265), .A2(MEM_stage_inst_dmem_n1264), .ZN(MEM_stage_inst_dmem_n1266) );
NAND2_X1 MEM_stage_inst_dmem_U1431 ( .A1(MEM_stage_inst_dmem_n1263), .A2(MEM_stage_inst_dmem_n1262), .ZN(MEM_stage_inst_dmem_n1264) );
NOR2_X1 MEM_stage_inst_dmem_U1430 ( .A1(MEM_stage_inst_dmem_n1261), .A2(MEM_stage_inst_dmem_n1260), .ZN(MEM_stage_inst_dmem_n1262) );
NAND2_X1 MEM_stage_inst_dmem_U1429 ( .A1(MEM_stage_inst_dmem_n1259), .A2(MEM_stage_inst_dmem_n1258), .ZN(MEM_stage_inst_dmem_n1260) );
NAND2_X1 MEM_stage_inst_dmem_U1428 ( .A1(MEM_stage_inst_dmem_ram_2273), .A2(MEM_stage_inst_dmem_n3152), .ZN(MEM_stage_inst_dmem_n1258) );
NAND2_X1 MEM_stage_inst_dmem_U1427 ( .A1(MEM_stage_inst_dmem_ram_2977), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n1259) );
NAND2_X1 MEM_stage_inst_dmem_U1426 ( .A1(MEM_stage_inst_dmem_n1257), .A2(MEM_stage_inst_dmem_n1256), .ZN(MEM_stage_inst_dmem_n1261) );
NAND2_X1 MEM_stage_inst_dmem_U1425 ( .A1(MEM_stage_inst_dmem_ram_2897), .A2(MEM_stage_inst_dmem_n3141), .ZN(MEM_stage_inst_dmem_n1256) );
NAND2_X1 MEM_stage_inst_dmem_U1424 ( .A1(MEM_stage_inst_dmem_ram_2561), .A2(MEM_stage_inst_dmem_n3182), .ZN(MEM_stage_inst_dmem_n1257) );
NOR2_X1 MEM_stage_inst_dmem_U1423 ( .A1(MEM_stage_inst_dmem_n1255), .A2(MEM_stage_inst_dmem_n1254), .ZN(MEM_stage_inst_dmem_n1263) );
NAND2_X1 MEM_stage_inst_dmem_U1422 ( .A1(MEM_stage_inst_dmem_n1253), .A2(MEM_stage_inst_dmem_n1252), .ZN(MEM_stage_inst_dmem_n1254) );
NAND2_X1 MEM_stage_inst_dmem_U1421 ( .A1(MEM_stage_inst_dmem_ram_2161), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n1252) );
NAND2_X1 MEM_stage_inst_dmem_U1420 ( .A1(MEM_stage_inst_dmem_ram_2433), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n1253) );
NAND2_X1 MEM_stage_inst_dmem_U1419 ( .A1(MEM_stage_inst_dmem_n1251), .A2(MEM_stage_inst_dmem_n1250), .ZN(MEM_stage_inst_dmem_n1255) );
NAND2_X1 MEM_stage_inst_dmem_U1418 ( .A1(MEM_stage_inst_dmem_ram_3041), .A2(MEM_stage_inst_dmem_n3113), .ZN(MEM_stage_inst_dmem_n1250) );
NAND2_X1 MEM_stage_inst_dmem_U1417 ( .A1(MEM_stage_inst_dmem_ram_2193), .A2(MEM_stage_inst_dmem_n44), .ZN(MEM_stage_inst_dmem_n1251) );
NAND2_X1 MEM_stage_inst_dmem_U1416 ( .A1(MEM_stage_inst_dmem_n1249), .A2(MEM_stage_inst_dmem_n1248), .ZN(MEM_stage_inst_dmem_n1265) );
NOR2_X1 MEM_stage_inst_dmem_U1415 ( .A1(MEM_stage_inst_dmem_n1247), .A2(MEM_stage_inst_dmem_n1246), .ZN(MEM_stage_inst_dmem_n1248) );
NAND2_X1 MEM_stage_inst_dmem_U1414 ( .A1(MEM_stage_inst_dmem_n1245), .A2(MEM_stage_inst_dmem_n1244), .ZN(MEM_stage_inst_dmem_n1246) );
NAND2_X1 MEM_stage_inst_dmem_U1413 ( .A1(MEM_stage_inst_dmem_ram_2945), .A2(MEM_stage_inst_dmem_n3123), .ZN(MEM_stage_inst_dmem_n1244) );
NAND2_X1 MEM_stage_inst_dmem_U1412 ( .A1(MEM_stage_inst_dmem_ram_2145), .A2(MEM_stage_inst_dmem_n3179), .ZN(MEM_stage_inst_dmem_n1245) );
NAND2_X1 MEM_stage_inst_dmem_U1411 ( .A1(MEM_stage_inst_dmem_n1243), .A2(MEM_stage_inst_dmem_n1242), .ZN(MEM_stage_inst_dmem_n1247) );
NAND2_X1 MEM_stage_inst_dmem_U1410 ( .A1(MEM_stage_inst_dmem_ram_2529), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n1242) );
NAND2_X1 MEM_stage_inst_dmem_U1409 ( .A1(MEM_stage_inst_dmem_ram_2849), .A2(MEM_stage_inst_dmem_n3137), .ZN(MEM_stage_inst_dmem_n1243) );
NOR2_X1 MEM_stage_inst_dmem_U1408 ( .A1(MEM_stage_inst_dmem_n1241), .A2(MEM_stage_inst_dmem_n1240), .ZN(MEM_stage_inst_dmem_n1249) );
NAND2_X1 MEM_stage_inst_dmem_U1407 ( .A1(MEM_stage_inst_dmem_n1239), .A2(MEM_stage_inst_dmem_n1238), .ZN(MEM_stage_inst_dmem_n1240) );
NAND2_X1 MEM_stage_inst_dmem_U1406 ( .A1(MEM_stage_inst_dmem_ram_2545), .A2(MEM_stage_inst_dmem_n3170), .ZN(MEM_stage_inst_dmem_n1238) );
NAND2_X1 MEM_stage_inst_dmem_U1405 ( .A1(MEM_stage_inst_dmem_ram_2769), .A2(MEM_stage_inst_dmem_n3112), .ZN(MEM_stage_inst_dmem_n1239) );
NAND2_X1 MEM_stage_inst_dmem_U1404 ( .A1(MEM_stage_inst_dmem_n1237), .A2(MEM_stage_inst_dmem_n1236), .ZN(MEM_stage_inst_dmem_n1241) );
NAND2_X1 MEM_stage_inst_dmem_U1403 ( .A1(MEM_stage_inst_dmem_ram_2081), .A2(MEM_stage_inst_dmem_n3092), .ZN(MEM_stage_inst_dmem_n1236) );
NAND2_X1 MEM_stage_inst_dmem_U1402 ( .A1(MEM_stage_inst_dmem_ram_3025), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n1237) );
NOR2_X1 MEM_stage_inst_dmem_U1401 ( .A1(MEM_stage_inst_dmem_n1235), .A2(MEM_stage_inst_dmem_n1234), .ZN(MEM_stage_inst_dmem_n1267) );
NAND2_X1 MEM_stage_inst_dmem_U1400 ( .A1(MEM_stage_inst_dmem_n1233), .A2(MEM_stage_inst_dmem_n1232), .ZN(MEM_stage_inst_dmem_n1234) );
NOR2_X1 MEM_stage_inst_dmem_U1399 ( .A1(MEM_stage_inst_dmem_n1231), .A2(MEM_stage_inst_dmem_n1230), .ZN(MEM_stage_inst_dmem_n1232) );
NAND2_X1 MEM_stage_inst_dmem_U1398 ( .A1(MEM_stage_inst_dmem_n1229), .A2(MEM_stage_inst_dmem_n1228), .ZN(MEM_stage_inst_dmem_n1230) );
NAND2_X1 MEM_stage_inst_dmem_U1397 ( .A1(MEM_stage_inst_dmem_ram_2465), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n1228) );
NAND2_X1 MEM_stage_inst_dmem_U1396 ( .A1(MEM_stage_inst_dmem_ram_2833), .A2(MEM_stage_inst_dmem_n3191), .ZN(MEM_stage_inst_dmem_n1229) );
NAND2_X1 MEM_stage_inst_dmem_U1395 ( .A1(MEM_stage_inst_dmem_n1227), .A2(MEM_stage_inst_dmem_n1226), .ZN(MEM_stage_inst_dmem_n1231) );
NAND2_X1 MEM_stage_inst_dmem_U1394 ( .A1(MEM_stage_inst_dmem_ram_2321), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n1226) );
NAND2_X1 MEM_stage_inst_dmem_U1393 ( .A1(MEM_stage_inst_dmem_ram_2337), .A2(MEM_stage_inst_dmem_n3209), .ZN(MEM_stage_inst_dmem_n1227) );
NOR2_X1 MEM_stage_inst_dmem_U1392 ( .A1(MEM_stage_inst_dmem_n1225), .A2(MEM_stage_inst_dmem_n1224), .ZN(MEM_stage_inst_dmem_n1233) );
NAND2_X1 MEM_stage_inst_dmem_U1391 ( .A1(MEM_stage_inst_dmem_n1223), .A2(MEM_stage_inst_dmem_n1222), .ZN(MEM_stage_inst_dmem_n1224) );
NAND2_X1 MEM_stage_inst_dmem_U1390 ( .A1(MEM_stage_inst_dmem_ram_2513), .A2(MEM_stage_inst_dmem_n3174), .ZN(MEM_stage_inst_dmem_n1222) );
NAND2_X1 MEM_stage_inst_dmem_U1389 ( .A1(MEM_stage_inst_dmem_ram_2209), .A2(MEM_stage_inst_dmem_n3081), .ZN(MEM_stage_inst_dmem_n1223) );
NAND2_X1 MEM_stage_inst_dmem_U1388 ( .A1(MEM_stage_inst_dmem_n1221), .A2(MEM_stage_inst_dmem_n1220), .ZN(MEM_stage_inst_dmem_n1225) );
NAND2_X1 MEM_stage_inst_dmem_U1387 ( .A1(MEM_stage_inst_dmem_ram_2113), .A2(MEM_stage_inst_dmem_n3102), .ZN(MEM_stage_inst_dmem_n1220) );
NAND2_X1 MEM_stage_inst_dmem_U1386 ( .A1(MEM_stage_inst_dmem_ram_2673), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n1221) );
NAND2_X1 MEM_stage_inst_dmem_U1385 ( .A1(MEM_stage_inst_dmem_n1219), .A2(MEM_stage_inst_dmem_n1218), .ZN(MEM_stage_inst_dmem_n1235) );
NOR2_X1 MEM_stage_inst_dmem_U1384 ( .A1(MEM_stage_inst_dmem_n1217), .A2(MEM_stage_inst_dmem_n1216), .ZN(MEM_stage_inst_dmem_n1218) );
NAND2_X1 MEM_stage_inst_dmem_U1383 ( .A1(MEM_stage_inst_dmem_n1215), .A2(MEM_stage_inst_dmem_n1214), .ZN(MEM_stage_inst_dmem_n1216) );
NAND2_X1 MEM_stage_inst_dmem_U1382 ( .A1(MEM_stage_inst_dmem_ram_2865), .A2(MEM_stage_inst_dmem_n46), .ZN(MEM_stage_inst_dmem_n1214) );
NAND2_X1 MEM_stage_inst_dmem_U1381 ( .A1(MEM_stage_inst_dmem_ram_2497), .A2(MEM_stage_inst_dmem_n3173), .ZN(MEM_stage_inst_dmem_n1215) );
NAND2_X1 MEM_stage_inst_dmem_U1380 ( .A1(MEM_stage_inst_dmem_n1213), .A2(MEM_stage_inst_dmem_n1212), .ZN(MEM_stage_inst_dmem_n1217) );
NAND2_X1 MEM_stage_inst_dmem_U1379 ( .A1(MEM_stage_inst_dmem_ram_2753), .A2(MEM_stage_inst_dmem_n3192), .ZN(MEM_stage_inst_dmem_n1212) );
NAND2_X1 MEM_stage_inst_dmem_U1378 ( .A1(MEM_stage_inst_dmem_ram_2625), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n1213) );
NOR2_X1 MEM_stage_inst_dmem_U1377 ( .A1(MEM_stage_inst_dmem_n1211), .A2(MEM_stage_inst_dmem_n1210), .ZN(MEM_stage_inst_dmem_n1219) );
NAND2_X1 MEM_stage_inst_dmem_U1376 ( .A1(MEM_stage_inst_dmem_n1209), .A2(MEM_stage_inst_dmem_n1208), .ZN(MEM_stage_inst_dmem_n1210) );
NAND2_X1 MEM_stage_inst_dmem_U1375 ( .A1(MEM_stage_inst_dmem_ram_2241), .A2(MEM_stage_inst_dmem_n3082), .ZN(MEM_stage_inst_dmem_n1208) );
NAND2_X1 MEM_stage_inst_dmem_U1374 ( .A1(MEM_stage_inst_dmem_ram_2721), .A2(MEM_stage_inst_dmem_n3155), .ZN(MEM_stage_inst_dmem_n1209) );
NAND2_X1 MEM_stage_inst_dmem_U1373 ( .A1(MEM_stage_inst_dmem_n1207), .A2(MEM_stage_inst_dmem_n1206), .ZN(MEM_stage_inst_dmem_n1211) );
NAND2_X1 MEM_stage_inst_dmem_U1372 ( .A1(MEM_stage_inst_dmem_ram_2401), .A2(MEM_stage_inst_dmem_n3217), .ZN(MEM_stage_inst_dmem_n1206) );
NAND2_X1 MEM_stage_inst_dmem_U1371 ( .A1(MEM_stage_inst_dmem_ram_2961), .A2(MEM_stage_inst_dmem_n3073), .ZN(MEM_stage_inst_dmem_n1207) );
NAND2_X1 MEM_stage_inst_dmem_U1370 ( .A1(MEM_stage_inst_dmem_n1205), .A2(MEM_stage_inst_dmem_n1204), .ZN(MEM_stage_inst_dmem_n1269) );
NOR2_X1 MEM_stage_inst_dmem_U1369 ( .A1(MEM_stage_inst_dmem_n1203), .A2(MEM_stage_inst_dmem_n1202), .ZN(MEM_stage_inst_dmem_n1204) );
NAND2_X1 MEM_stage_inst_dmem_U1368 ( .A1(MEM_stage_inst_dmem_n1201), .A2(MEM_stage_inst_dmem_n1200), .ZN(MEM_stage_inst_dmem_n1202) );
NOR2_X1 MEM_stage_inst_dmem_U1367 ( .A1(MEM_stage_inst_dmem_n1199), .A2(MEM_stage_inst_dmem_n1198), .ZN(MEM_stage_inst_dmem_n1200) );
NAND2_X1 MEM_stage_inst_dmem_U1366 ( .A1(MEM_stage_inst_dmem_n1197), .A2(MEM_stage_inst_dmem_n1196), .ZN(MEM_stage_inst_dmem_n1198) );
NAND2_X1 MEM_stage_inst_dmem_U1365 ( .A1(MEM_stage_inst_dmem_ram_2353), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n1196) );
NAND2_X1 MEM_stage_inst_dmem_U1364 ( .A1(MEM_stage_inst_dmem_ram_2129), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n1197) );
NAND2_X1 MEM_stage_inst_dmem_U1363 ( .A1(MEM_stage_inst_dmem_n1195), .A2(MEM_stage_inst_dmem_n1194), .ZN(MEM_stage_inst_dmem_n1199) );
NAND2_X1 MEM_stage_inst_dmem_U1362 ( .A1(MEM_stage_inst_dmem_ram_2993), .A2(MEM_stage_inst_dmem_n3163), .ZN(MEM_stage_inst_dmem_n1194) );
NAND2_X1 MEM_stage_inst_dmem_U1361 ( .A1(MEM_stage_inst_dmem_ram_2225), .A2(MEM_stage_inst_dmem_n55), .ZN(MEM_stage_inst_dmem_n1195) );
NOR2_X1 MEM_stage_inst_dmem_U1360 ( .A1(MEM_stage_inst_dmem_n1193), .A2(MEM_stage_inst_dmem_n1192), .ZN(MEM_stage_inst_dmem_n1201) );
NAND2_X1 MEM_stage_inst_dmem_U1359 ( .A1(MEM_stage_inst_dmem_n1191), .A2(MEM_stage_inst_dmem_n1190), .ZN(MEM_stage_inst_dmem_n1192) );
NAND2_X1 MEM_stage_inst_dmem_U1358 ( .A1(MEM_stage_inst_dmem_ram_2177), .A2(MEM_stage_inst_dmem_n3130), .ZN(MEM_stage_inst_dmem_n1190) );
NAND2_X1 MEM_stage_inst_dmem_U1357 ( .A1(MEM_stage_inst_dmem_ram_2049), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n1191) );
NAND2_X1 MEM_stage_inst_dmem_U1356 ( .A1(MEM_stage_inst_dmem_n1189), .A2(MEM_stage_inst_dmem_n1188), .ZN(MEM_stage_inst_dmem_n1193) );
NAND2_X1 MEM_stage_inst_dmem_U1355 ( .A1(MEM_stage_inst_dmem_ram_2097), .A2(MEM_stage_inst_dmem_n3103), .ZN(MEM_stage_inst_dmem_n1188) );
NAND2_X1 MEM_stage_inst_dmem_U1354 ( .A1(MEM_stage_inst_dmem_ram_3057), .A2(MEM_stage_inst_dmem_n3199), .ZN(MEM_stage_inst_dmem_n1189) );
NAND2_X1 MEM_stage_inst_dmem_U1353 ( .A1(MEM_stage_inst_dmem_n1187), .A2(MEM_stage_inst_dmem_n1186), .ZN(MEM_stage_inst_dmem_n1203) );
NOR2_X1 MEM_stage_inst_dmem_U1352 ( .A1(MEM_stage_inst_dmem_n1185), .A2(MEM_stage_inst_dmem_n1184), .ZN(MEM_stage_inst_dmem_n1186) );
NAND2_X1 MEM_stage_inst_dmem_U1351 ( .A1(MEM_stage_inst_dmem_n1183), .A2(MEM_stage_inst_dmem_n1182), .ZN(MEM_stage_inst_dmem_n1184) );
NAND2_X1 MEM_stage_inst_dmem_U1350 ( .A1(MEM_stage_inst_dmem_ram_2817), .A2(MEM_stage_inst_dmem_n37), .ZN(MEM_stage_inst_dmem_n1182) );
NAND2_X1 MEM_stage_inst_dmem_U1349 ( .A1(MEM_stage_inst_dmem_ram_2801), .A2(MEM_stage_inst_dmem_n3202), .ZN(MEM_stage_inst_dmem_n1183) );
NAND2_X1 MEM_stage_inst_dmem_U1348 ( .A1(MEM_stage_inst_dmem_n1181), .A2(MEM_stage_inst_dmem_n1180), .ZN(MEM_stage_inst_dmem_n1185) );
NAND2_X1 MEM_stage_inst_dmem_U1347 ( .A1(MEM_stage_inst_dmem_ram_2289), .A2(MEM_stage_inst_dmem_n39), .ZN(MEM_stage_inst_dmem_n1180) );
NAND2_X1 MEM_stage_inst_dmem_U1346 ( .A1(MEM_stage_inst_dmem_ram_2593), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n1181) );
NOR2_X1 MEM_stage_inst_dmem_U1345 ( .A1(MEM_stage_inst_dmem_n1179), .A2(MEM_stage_inst_dmem_n1178), .ZN(MEM_stage_inst_dmem_n1187) );
NAND2_X1 MEM_stage_inst_dmem_U1344 ( .A1(MEM_stage_inst_dmem_n1177), .A2(MEM_stage_inst_dmem_n1176), .ZN(MEM_stage_inst_dmem_n1178) );
NAND2_X1 MEM_stage_inst_dmem_U1343 ( .A1(MEM_stage_inst_dmem_ram_2369), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n1176) );
NAND2_X1 MEM_stage_inst_dmem_U1342 ( .A1(MEM_stage_inst_dmem_ram_2577), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n1177) );
NAND2_X1 MEM_stage_inst_dmem_U1341 ( .A1(MEM_stage_inst_dmem_n1175), .A2(MEM_stage_inst_dmem_n1174), .ZN(MEM_stage_inst_dmem_n1179) );
NAND2_X1 MEM_stage_inst_dmem_U1340 ( .A1(MEM_stage_inst_dmem_ram_2641), .A2(MEM_stage_inst_dmem_n3140), .ZN(MEM_stage_inst_dmem_n1174) );
NAND2_X1 MEM_stage_inst_dmem_U1339 ( .A1(MEM_stage_inst_dmem_ram_2305), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n1175) );
NOR2_X1 MEM_stage_inst_dmem_U1338 ( .A1(MEM_stage_inst_dmem_n1173), .A2(MEM_stage_inst_dmem_n1172), .ZN(MEM_stage_inst_dmem_n1205) );
NAND2_X1 MEM_stage_inst_dmem_U1337 ( .A1(MEM_stage_inst_dmem_n1171), .A2(MEM_stage_inst_dmem_n1170), .ZN(MEM_stage_inst_dmem_n1172) );
NOR2_X1 MEM_stage_inst_dmem_U1336 ( .A1(MEM_stage_inst_dmem_n1169), .A2(MEM_stage_inst_dmem_n1168), .ZN(MEM_stage_inst_dmem_n1170) );
NAND2_X1 MEM_stage_inst_dmem_U1335 ( .A1(MEM_stage_inst_dmem_n1167), .A2(MEM_stage_inst_dmem_n1166), .ZN(MEM_stage_inst_dmem_n1168) );
NAND2_X1 MEM_stage_inst_dmem_U1334 ( .A1(MEM_stage_inst_dmem_ram_2065), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n1166) );
NAND2_X1 MEM_stage_inst_dmem_U1333 ( .A1(MEM_stage_inst_dmem_ram_2385), .A2(MEM_stage_inst_dmem_n3216), .ZN(MEM_stage_inst_dmem_n1167) );
NAND2_X1 MEM_stage_inst_dmem_U1332 ( .A1(MEM_stage_inst_dmem_n1165), .A2(MEM_stage_inst_dmem_n1164), .ZN(MEM_stage_inst_dmem_n1169) );
NAND2_X1 MEM_stage_inst_dmem_U1331 ( .A1(MEM_stage_inst_dmem_ram_2449), .A2(MEM_stage_inst_dmem_n3160), .ZN(MEM_stage_inst_dmem_n1164) );
NAND2_X1 MEM_stage_inst_dmem_U1330 ( .A1(MEM_stage_inst_dmem_ram_2657), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n1165) );
NOR2_X1 MEM_stage_inst_dmem_U1329 ( .A1(MEM_stage_inst_dmem_n1163), .A2(MEM_stage_inst_dmem_n1162), .ZN(MEM_stage_inst_dmem_n1171) );
NAND2_X1 MEM_stage_inst_dmem_U1328 ( .A1(MEM_stage_inst_dmem_n1161), .A2(MEM_stage_inst_dmem_n1160), .ZN(MEM_stage_inst_dmem_n1162) );
NAND2_X1 MEM_stage_inst_dmem_U1327 ( .A1(MEM_stage_inst_dmem_ram_2609), .A2(MEM_stage_inst_dmem_n3085), .ZN(MEM_stage_inst_dmem_n1160) );
NAND2_X1 MEM_stage_inst_dmem_U1326 ( .A1(MEM_stage_inst_dmem_ram_2785), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n1161) );
NAND2_X1 MEM_stage_inst_dmem_U1325 ( .A1(MEM_stage_inst_dmem_n1159), .A2(MEM_stage_inst_dmem_n1158), .ZN(MEM_stage_inst_dmem_n1163) );
NAND2_X1 MEM_stage_inst_dmem_U1324 ( .A1(MEM_stage_inst_dmem_ram_2913), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n1158) );
NAND2_X1 MEM_stage_inst_dmem_U1323 ( .A1(MEM_stage_inst_dmem_ram_2881), .A2(MEM_stage_inst_dmem_n3120), .ZN(MEM_stage_inst_dmem_n1159) );
NAND2_X1 MEM_stage_inst_dmem_U1322 ( .A1(MEM_stage_inst_dmem_n1157), .A2(MEM_stage_inst_dmem_n1156), .ZN(MEM_stage_inst_dmem_n1173) );
NOR2_X1 MEM_stage_inst_dmem_U1321 ( .A1(MEM_stage_inst_dmem_n1155), .A2(MEM_stage_inst_dmem_n1154), .ZN(MEM_stage_inst_dmem_n1156) );
NAND2_X1 MEM_stage_inst_dmem_U1320 ( .A1(MEM_stage_inst_dmem_n1153), .A2(MEM_stage_inst_dmem_n1152), .ZN(MEM_stage_inst_dmem_n1154) );
NAND2_X1 MEM_stage_inst_dmem_U1319 ( .A1(MEM_stage_inst_dmem_ram_2929), .A2(MEM_stage_inst_dmem_n3099), .ZN(MEM_stage_inst_dmem_n1152) );
NAND2_X1 MEM_stage_inst_dmem_U1318 ( .A1(MEM_stage_inst_dmem_ram_2689), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n1153) );
NAND2_X1 MEM_stage_inst_dmem_U1317 ( .A1(MEM_stage_inst_dmem_n1151), .A2(MEM_stage_inst_dmem_n1150), .ZN(MEM_stage_inst_dmem_n1155) );
NAND2_X1 MEM_stage_inst_dmem_U1316 ( .A1(MEM_stage_inst_dmem_ram_2481), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n1150) );
NAND2_X1 MEM_stage_inst_dmem_U1315 ( .A1(MEM_stage_inst_dmem_ram_2705), .A2(MEM_stage_inst_dmem_n3076), .ZN(MEM_stage_inst_dmem_n1151) );
NOR2_X1 MEM_stage_inst_dmem_U1314 ( .A1(MEM_stage_inst_dmem_n1149), .A2(MEM_stage_inst_dmem_n1148), .ZN(MEM_stage_inst_dmem_n1157) );
NAND2_X1 MEM_stage_inst_dmem_U1313 ( .A1(MEM_stage_inst_dmem_n1147), .A2(MEM_stage_inst_dmem_n1146), .ZN(MEM_stage_inst_dmem_n1148) );
NAND2_X1 MEM_stage_inst_dmem_U1312 ( .A1(MEM_stage_inst_dmem_ram_2257), .A2(MEM_stage_inst_dmem_n3220), .ZN(MEM_stage_inst_dmem_n1146) );
NAND2_X1 MEM_stage_inst_dmem_U1311 ( .A1(MEM_stage_inst_dmem_ram_2417), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n1147) );
NAND2_X1 MEM_stage_inst_dmem_U1310 ( .A1(MEM_stage_inst_dmem_n1145), .A2(MEM_stage_inst_dmem_n1144), .ZN(MEM_stage_inst_dmem_n1149) );
NAND2_X1 MEM_stage_inst_dmem_U1309 ( .A1(MEM_stage_inst_dmem_ram_3009), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n1144) );
NAND2_X1 MEM_stage_inst_dmem_U1308 ( .A1(MEM_stage_inst_dmem_ram_2737), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n1145) );
NOR2_X1 MEM_stage_inst_dmem_U1307 ( .A1(MEM_stage_inst_dmem_n1143), .A2(MEM_stage_inst_dmem_n8551), .ZN(MEM_stage_inst_dmem_n1272) );
NOR2_X1 MEM_stage_inst_dmem_U1306 ( .A1(MEM_stage_inst_dmem_n1142), .A2(MEM_stage_inst_dmem_n1141), .ZN(MEM_stage_inst_dmem_n1143) );
NAND2_X1 MEM_stage_inst_dmem_U1305 ( .A1(MEM_stage_inst_dmem_n1140), .A2(MEM_stage_inst_dmem_n1139), .ZN(MEM_stage_inst_dmem_n1141) );
NOR2_X1 MEM_stage_inst_dmem_U1304 ( .A1(MEM_stage_inst_dmem_n1138), .A2(MEM_stage_inst_dmem_n1137), .ZN(MEM_stage_inst_dmem_n1139) );
NAND2_X1 MEM_stage_inst_dmem_U1303 ( .A1(MEM_stage_inst_dmem_n1136), .A2(MEM_stage_inst_dmem_n1135), .ZN(MEM_stage_inst_dmem_n1137) );
NOR2_X1 MEM_stage_inst_dmem_U1302 ( .A1(MEM_stage_inst_dmem_n1134), .A2(MEM_stage_inst_dmem_n1133), .ZN(MEM_stage_inst_dmem_n1135) );
NAND2_X1 MEM_stage_inst_dmem_U1301 ( .A1(MEM_stage_inst_dmem_n1132), .A2(MEM_stage_inst_dmem_n1131), .ZN(MEM_stage_inst_dmem_n1133) );
NAND2_X1 MEM_stage_inst_dmem_U1300 ( .A1(MEM_stage_inst_dmem_ram_129), .A2(MEM_stage_inst_dmem_n61), .ZN(MEM_stage_inst_dmem_n1131) );
NAND2_X1 MEM_stage_inst_dmem_U1299 ( .A1(MEM_stage_inst_dmem_ram_529), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n1132) );
NAND2_X1 MEM_stage_inst_dmem_U1298 ( .A1(MEM_stage_inst_dmem_n1130), .A2(MEM_stage_inst_dmem_n1129), .ZN(MEM_stage_inst_dmem_n1134) );
NAND2_X1 MEM_stage_inst_dmem_U1297 ( .A1(MEM_stage_inst_dmem_ram_929), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n1129) );
NAND2_X1 MEM_stage_inst_dmem_U1296 ( .A1(MEM_stage_inst_dmem_ram_657), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n1130) );
NOR2_X1 MEM_stage_inst_dmem_U1295 ( .A1(MEM_stage_inst_dmem_n1128), .A2(MEM_stage_inst_dmem_n1127), .ZN(MEM_stage_inst_dmem_n1136) );
NAND2_X1 MEM_stage_inst_dmem_U1294 ( .A1(MEM_stage_inst_dmem_n1126), .A2(MEM_stage_inst_dmem_n1125), .ZN(MEM_stage_inst_dmem_n1127) );
NAND2_X1 MEM_stage_inst_dmem_U1293 ( .A1(MEM_stage_inst_dmem_ram_817), .A2(MEM_stage_inst_dmem_n8005), .ZN(MEM_stage_inst_dmem_n1125) );
NAND2_X1 MEM_stage_inst_dmem_U1292 ( .A1(MEM_stage_inst_dmem_ram_177), .A2(MEM_stage_inst_dmem_n55), .ZN(MEM_stage_inst_dmem_n1126) );
NAND2_X1 MEM_stage_inst_dmem_U1291 ( .A1(MEM_stage_inst_dmem_n1124), .A2(MEM_stage_inst_dmem_n1123), .ZN(MEM_stage_inst_dmem_n1128) );
NAND2_X1 MEM_stage_inst_dmem_U1290 ( .A1(MEM_stage_inst_dmem_ram_401), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n1123) );
NAND2_X1 MEM_stage_inst_dmem_U1289 ( .A1(MEM_stage_inst_dmem_ram_513), .A2(MEM_stage_inst_dmem_n71), .ZN(MEM_stage_inst_dmem_n1124) );
NAND2_X1 MEM_stage_inst_dmem_U1288 ( .A1(MEM_stage_inst_dmem_n1122), .A2(MEM_stage_inst_dmem_n1121), .ZN(MEM_stage_inst_dmem_n1138) );
NOR2_X1 MEM_stage_inst_dmem_U1287 ( .A1(MEM_stage_inst_dmem_n1120), .A2(MEM_stage_inst_dmem_n1119), .ZN(MEM_stage_inst_dmem_n1121) );
NAND2_X1 MEM_stage_inst_dmem_U1286 ( .A1(MEM_stage_inst_dmem_n1118), .A2(MEM_stage_inst_dmem_n1117), .ZN(MEM_stage_inst_dmem_n1119) );
NAND2_X1 MEM_stage_inst_dmem_U1285 ( .A1(MEM_stage_inst_dmem_ram_753), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n1117) );
NAND2_X1 MEM_stage_inst_dmem_U1284 ( .A1(MEM_stage_inst_dmem_ram_465), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n1118) );
NAND2_X1 MEM_stage_inst_dmem_U1283 ( .A1(MEM_stage_inst_dmem_n1116), .A2(MEM_stage_inst_dmem_n1115), .ZN(MEM_stage_inst_dmem_n1120) );
NAND2_X1 MEM_stage_inst_dmem_U1282 ( .A1(MEM_stage_inst_dmem_ram_561), .A2(MEM_stage_inst_dmem_n41), .ZN(MEM_stage_inst_dmem_n1115) );
NAND2_X1 MEM_stage_inst_dmem_U1281 ( .A1(MEM_stage_inst_dmem_ram_545), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n1116) );
NOR2_X1 MEM_stage_inst_dmem_U1280 ( .A1(MEM_stage_inst_dmem_n1114), .A2(MEM_stage_inst_dmem_n1113), .ZN(MEM_stage_inst_dmem_n1122) );
NAND2_X1 MEM_stage_inst_dmem_U1279 ( .A1(MEM_stage_inst_dmem_n1112), .A2(MEM_stage_inst_dmem_n1111), .ZN(MEM_stage_inst_dmem_n1113) );
NAND2_X1 MEM_stage_inst_dmem_U1278 ( .A1(MEM_stage_inst_dmem_ram_273), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n1111) );
NAND2_X1 MEM_stage_inst_dmem_U1277 ( .A1(MEM_stage_inst_dmem_ram_369), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n1112) );
NAND2_X1 MEM_stage_inst_dmem_U1276 ( .A1(MEM_stage_inst_dmem_n1110), .A2(MEM_stage_inst_dmem_n1109), .ZN(MEM_stage_inst_dmem_n1114) );
NAND2_X1 MEM_stage_inst_dmem_U1275 ( .A1(MEM_stage_inst_dmem_ram_993), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n1109) );
NAND2_X1 MEM_stage_inst_dmem_U1274 ( .A1(MEM_stage_inst_dmem_ram_977), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n1110) );
NOR2_X1 MEM_stage_inst_dmem_U1273 ( .A1(MEM_stage_inst_dmem_n1108), .A2(MEM_stage_inst_dmem_n1107), .ZN(MEM_stage_inst_dmem_n1140) );
NAND2_X1 MEM_stage_inst_dmem_U1272 ( .A1(MEM_stage_inst_dmem_n1106), .A2(MEM_stage_inst_dmem_n1105), .ZN(MEM_stage_inst_dmem_n1107) );
NOR2_X1 MEM_stage_inst_dmem_U1271 ( .A1(MEM_stage_inst_dmem_n1104), .A2(MEM_stage_inst_dmem_n1103), .ZN(MEM_stage_inst_dmem_n1105) );
NAND2_X1 MEM_stage_inst_dmem_U1270 ( .A1(MEM_stage_inst_dmem_n1102), .A2(MEM_stage_inst_dmem_n1101), .ZN(MEM_stage_inst_dmem_n1103) );
NAND2_X1 MEM_stage_inst_dmem_U1269 ( .A1(MEM_stage_inst_dmem_ram_913), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n1101) );
NAND2_X1 MEM_stage_inst_dmem_U1268 ( .A1(MEM_stage_inst_dmem_ram_241), .A2(MEM_stage_inst_dmem_n7914), .ZN(MEM_stage_inst_dmem_n1102) );
NAND2_X1 MEM_stage_inst_dmem_U1267 ( .A1(MEM_stage_inst_dmem_n1100), .A2(MEM_stage_inst_dmem_n1099), .ZN(MEM_stage_inst_dmem_n1104) );
NAND2_X1 MEM_stage_inst_dmem_U1266 ( .A1(MEM_stage_inst_dmem_ram_865), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n1099) );
NAND2_X1 MEM_stage_inst_dmem_U1265 ( .A1(MEM_stage_inst_dmem_ram_209), .A2(MEM_stage_inst_dmem_n51), .ZN(MEM_stage_inst_dmem_n1100) );
NOR2_X1 MEM_stage_inst_dmem_U1264 ( .A1(MEM_stage_inst_dmem_n1098), .A2(MEM_stage_inst_dmem_n1097), .ZN(MEM_stage_inst_dmem_n1106) );
NAND2_X1 MEM_stage_inst_dmem_U1263 ( .A1(MEM_stage_inst_dmem_n1096), .A2(MEM_stage_inst_dmem_n1095), .ZN(MEM_stage_inst_dmem_n1097) );
NAND2_X1 MEM_stage_inst_dmem_U1262 ( .A1(MEM_stage_inst_dmem_ram_385), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n1095) );
NAND2_X1 MEM_stage_inst_dmem_U1261 ( .A1(MEM_stage_inst_dmem_ram_721), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n1096) );
NAND2_X1 MEM_stage_inst_dmem_U1260 ( .A1(MEM_stage_inst_dmem_n1094), .A2(MEM_stage_inst_dmem_n1093), .ZN(MEM_stage_inst_dmem_n1098) );
NAND2_X1 MEM_stage_inst_dmem_U1259 ( .A1(MEM_stage_inst_dmem_ram_17), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n1093) );
NAND2_X1 MEM_stage_inst_dmem_U1258 ( .A1(MEM_stage_inst_dmem_ram_289), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n1094) );
NAND2_X1 MEM_stage_inst_dmem_U1257 ( .A1(MEM_stage_inst_dmem_n1092), .A2(MEM_stage_inst_dmem_n1091), .ZN(MEM_stage_inst_dmem_n1108) );
NOR2_X1 MEM_stage_inst_dmem_U1256 ( .A1(MEM_stage_inst_dmem_n1090), .A2(MEM_stage_inst_dmem_n1089), .ZN(MEM_stage_inst_dmem_n1091) );
NAND2_X1 MEM_stage_inst_dmem_U1255 ( .A1(MEM_stage_inst_dmem_n1088), .A2(MEM_stage_inst_dmem_n1087), .ZN(MEM_stage_inst_dmem_n1089) );
NAND2_X1 MEM_stage_inst_dmem_U1254 ( .A1(MEM_stage_inst_dmem_ram_225), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n1087) );
NAND2_X1 MEM_stage_inst_dmem_U1253 ( .A1(MEM_stage_inst_dmem_ram_449), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n1088) );
NAND2_X1 MEM_stage_inst_dmem_U1252 ( .A1(MEM_stage_inst_dmem_n1086), .A2(MEM_stage_inst_dmem_n1085), .ZN(MEM_stage_inst_dmem_n1090) );
NAND2_X1 MEM_stage_inst_dmem_U1251 ( .A1(MEM_stage_inst_dmem_ram_881), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n1085) );
NAND2_X1 MEM_stage_inst_dmem_U1250 ( .A1(MEM_stage_inst_dmem_ram_609), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n1086) );
NOR2_X1 MEM_stage_inst_dmem_U1249 ( .A1(MEM_stage_inst_dmem_n1084), .A2(MEM_stage_inst_dmem_n1083), .ZN(MEM_stage_inst_dmem_n1092) );
NAND2_X1 MEM_stage_inst_dmem_U1248 ( .A1(MEM_stage_inst_dmem_n1082), .A2(MEM_stage_inst_dmem_n1081), .ZN(MEM_stage_inst_dmem_n1083) );
NAND2_X1 MEM_stage_inst_dmem_U1247 ( .A1(MEM_stage_inst_dmem_ram_849), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n1081) );
NAND2_X1 MEM_stage_inst_dmem_U1246 ( .A1(MEM_stage_inst_dmem_ram_417), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n1082) );
NAND2_X1 MEM_stage_inst_dmem_U1245 ( .A1(MEM_stage_inst_dmem_n1080), .A2(MEM_stage_inst_dmem_n1079), .ZN(MEM_stage_inst_dmem_n1084) );
NAND2_X1 MEM_stage_inst_dmem_U1244 ( .A1(MEM_stage_inst_dmem_ram_145), .A2(MEM_stage_inst_dmem_n5807), .ZN(MEM_stage_inst_dmem_n1079) );
NAND2_X1 MEM_stage_inst_dmem_U1243 ( .A1(MEM_stage_inst_dmem_ram_257), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n1080) );
NAND2_X1 MEM_stage_inst_dmem_U1242 ( .A1(MEM_stage_inst_dmem_n1078), .A2(MEM_stage_inst_dmem_n1077), .ZN(MEM_stage_inst_dmem_n1142) );
NOR2_X1 MEM_stage_inst_dmem_U1241 ( .A1(MEM_stage_inst_dmem_n1076), .A2(MEM_stage_inst_dmem_n1075), .ZN(MEM_stage_inst_dmem_n1077) );
NAND2_X1 MEM_stage_inst_dmem_U1240 ( .A1(MEM_stage_inst_dmem_n1074), .A2(MEM_stage_inst_dmem_n1073), .ZN(MEM_stage_inst_dmem_n1075) );
NOR2_X1 MEM_stage_inst_dmem_U1239 ( .A1(MEM_stage_inst_dmem_n1072), .A2(MEM_stage_inst_dmem_n1071), .ZN(MEM_stage_inst_dmem_n1073) );
NAND2_X1 MEM_stage_inst_dmem_U1238 ( .A1(MEM_stage_inst_dmem_n1070), .A2(MEM_stage_inst_dmem_n1069), .ZN(MEM_stage_inst_dmem_n1071) );
NAND2_X1 MEM_stage_inst_dmem_U1237 ( .A1(MEM_stage_inst_dmem_ram_673), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n1069) );
NAND2_X1 MEM_stage_inst_dmem_U1236 ( .A1(MEM_stage_inst_dmem_ram_81), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n1070) );
NAND2_X1 MEM_stage_inst_dmem_U1235 ( .A1(MEM_stage_inst_dmem_n1068), .A2(MEM_stage_inst_dmem_n1067), .ZN(MEM_stage_inst_dmem_n1072) );
NAND2_X1 MEM_stage_inst_dmem_U1234 ( .A1(MEM_stage_inst_dmem_ram_321), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n1067) );
NAND2_X1 MEM_stage_inst_dmem_U1233 ( .A1(MEM_stage_inst_dmem_ram_785), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n1068) );
NOR2_X1 MEM_stage_inst_dmem_U1232 ( .A1(MEM_stage_inst_dmem_n1066), .A2(MEM_stage_inst_dmem_n1065), .ZN(MEM_stage_inst_dmem_n1074) );
NAND2_X1 MEM_stage_inst_dmem_U1231 ( .A1(MEM_stage_inst_dmem_n1064), .A2(MEM_stage_inst_dmem_n1063), .ZN(MEM_stage_inst_dmem_n1065) );
NAND2_X1 MEM_stage_inst_dmem_U1230 ( .A1(MEM_stage_inst_dmem_ram_961), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n1063) );
NAND2_X1 MEM_stage_inst_dmem_U1229 ( .A1(MEM_stage_inst_dmem_ram_737), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n1064) );
NAND2_X1 MEM_stage_inst_dmem_U1228 ( .A1(MEM_stage_inst_dmem_n1062), .A2(MEM_stage_inst_dmem_n1061), .ZN(MEM_stage_inst_dmem_n1066) );
NAND2_X1 MEM_stage_inst_dmem_U1227 ( .A1(MEM_stage_inst_dmem_ram_65), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n1061) );
NAND2_X1 MEM_stage_inst_dmem_U1226 ( .A1(MEM_stage_inst_dmem_ram_625), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n1062) );
NAND2_X1 MEM_stage_inst_dmem_U1225 ( .A1(MEM_stage_inst_dmem_n1060), .A2(MEM_stage_inst_dmem_n1059), .ZN(MEM_stage_inst_dmem_n1076) );
NOR2_X1 MEM_stage_inst_dmem_U1224 ( .A1(MEM_stage_inst_dmem_n1058), .A2(MEM_stage_inst_dmem_n1057), .ZN(MEM_stage_inst_dmem_n1059) );
NAND2_X1 MEM_stage_inst_dmem_U1223 ( .A1(MEM_stage_inst_dmem_n1056), .A2(MEM_stage_inst_dmem_n1055), .ZN(MEM_stage_inst_dmem_n1057) );
NAND2_X1 MEM_stage_inst_dmem_U1222 ( .A1(MEM_stage_inst_dmem_ram_897), .A2(MEM_stage_inst_dmem_n72), .ZN(MEM_stage_inst_dmem_n1055) );
NAND2_X1 MEM_stage_inst_dmem_U1221 ( .A1(MEM_stage_inst_dmem_ram_161), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n1056) );
NAND2_X1 MEM_stage_inst_dmem_U1220 ( .A1(MEM_stage_inst_dmem_n1054), .A2(MEM_stage_inst_dmem_n1053), .ZN(MEM_stage_inst_dmem_n1058) );
NAND2_X1 MEM_stage_inst_dmem_U1219 ( .A1(MEM_stage_inst_dmem_ram_945), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n1053) );
NAND2_X1 MEM_stage_inst_dmem_U1218 ( .A1(MEM_stage_inst_dmem_ram_641), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n1054) );
NOR2_X1 MEM_stage_inst_dmem_U1217 ( .A1(MEM_stage_inst_dmem_n1052), .A2(MEM_stage_inst_dmem_n1051), .ZN(MEM_stage_inst_dmem_n1060) );
NAND2_X1 MEM_stage_inst_dmem_U1216 ( .A1(MEM_stage_inst_dmem_n1050), .A2(MEM_stage_inst_dmem_n1049), .ZN(MEM_stage_inst_dmem_n1051) );
NAND2_X1 MEM_stage_inst_dmem_U1215 ( .A1(MEM_stage_inst_dmem_ram_433), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n1049) );
NAND2_X1 MEM_stage_inst_dmem_U1214 ( .A1(MEM_stage_inst_dmem_ram_481), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n1050) );
NAND2_X1 MEM_stage_inst_dmem_U1213 ( .A1(MEM_stage_inst_dmem_n1048), .A2(MEM_stage_inst_dmem_n1047), .ZN(MEM_stage_inst_dmem_n1052) );
NAND2_X1 MEM_stage_inst_dmem_U1212 ( .A1(MEM_stage_inst_dmem_ram_1009), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n1047) );
NAND2_X1 MEM_stage_inst_dmem_U1211 ( .A1(MEM_stage_inst_dmem_ram_593), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n1048) );
NOR2_X1 MEM_stage_inst_dmem_U1210 ( .A1(MEM_stage_inst_dmem_n1046), .A2(MEM_stage_inst_dmem_n1045), .ZN(MEM_stage_inst_dmem_n1078) );
NAND2_X1 MEM_stage_inst_dmem_U1209 ( .A1(MEM_stage_inst_dmem_n1044), .A2(MEM_stage_inst_dmem_n1043), .ZN(MEM_stage_inst_dmem_n1045) );
NOR2_X1 MEM_stage_inst_dmem_U1208 ( .A1(MEM_stage_inst_dmem_n1042), .A2(MEM_stage_inst_dmem_n1041), .ZN(MEM_stage_inst_dmem_n1043) );
NAND2_X1 MEM_stage_inst_dmem_U1207 ( .A1(MEM_stage_inst_dmem_n1040), .A2(MEM_stage_inst_dmem_n1039), .ZN(MEM_stage_inst_dmem_n1041) );
NAND2_X1 MEM_stage_inst_dmem_U1206 ( .A1(MEM_stage_inst_dmem_ram_801), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n1039) );
NAND2_X1 MEM_stage_inst_dmem_U1205 ( .A1(MEM_stage_inst_dmem_ram_689), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n1040) );
NAND2_X1 MEM_stage_inst_dmem_U1204 ( .A1(MEM_stage_inst_dmem_n1038), .A2(MEM_stage_inst_dmem_n1037), .ZN(MEM_stage_inst_dmem_n1042) );
NAND2_X1 MEM_stage_inst_dmem_U1203 ( .A1(MEM_stage_inst_dmem_ram_497), .A2(MEM_stage_inst_dmem_n8535), .ZN(MEM_stage_inst_dmem_n1037) );
NAND2_X1 MEM_stage_inst_dmem_U1202 ( .A1(MEM_stage_inst_dmem_ram_833), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n1038) );
NOR2_X1 MEM_stage_inst_dmem_U1201 ( .A1(MEM_stage_inst_dmem_n1036), .A2(MEM_stage_inst_dmem_n1035), .ZN(MEM_stage_inst_dmem_n1044) );
NAND2_X1 MEM_stage_inst_dmem_U1200 ( .A1(MEM_stage_inst_dmem_n1034), .A2(MEM_stage_inst_dmem_n1033), .ZN(MEM_stage_inst_dmem_n1035) );
NAND2_X1 MEM_stage_inst_dmem_U1199 ( .A1(MEM_stage_inst_dmem_ram_337), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n1033) );
NAND2_X1 MEM_stage_inst_dmem_U1198 ( .A1(MEM_stage_inst_dmem_ram_1), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n1034) );
NAND2_X1 MEM_stage_inst_dmem_U1197 ( .A1(MEM_stage_inst_dmem_n1032), .A2(MEM_stage_inst_dmem_n1031), .ZN(MEM_stage_inst_dmem_n1036) );
NAND2_X1 MEM_stage_inst_dmem_U1196 ( .A1(MEM_stage_inst_dmem_ram_193), .A2(MEM_stage_inst_dmem_n36), .ZN(MEM_stage_inst_dmem_n1031) );
NAND2_X1 MEM_stage_inst_dmem_U1195 ( .A1(MEM_stage_inst_dmem_ram_113), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n1032) );
NAND2_X1 MEM_stage_inst_dmem_U1194 ( .A1(MEM_stage_inst_dmem_n1030), .A2(MEM_stage_inst_dmem_n1029), .ZN(MEM_stage_inst_dmem_n1046) );
NOR2_X1 MEM_stage_inst_dmem_U1193 ( .A1(MEM_stage_inst_dmem_n1028), .A2(MEM_stage_inst_dmem_n1027), .ZN(MEM_stage_inst_dmem_n1029) );
NAND2_X1 MEM_stage_inst_dmem_U1192 ( .A1(MEM_stage_inst_dmem_n1026), .A2(MEM_stage_inst_dmem_n1025), .ZN(MEM_stage_inst_dmem_n1027) );
NAND2_X1 MEM_stage_inst_dmem_U1191 ( .A1(MEM_stage_inst_dmem_ram_769), .A2(MEM_stage_inst_dmem_n37), .ZN(MEM_stage_inst_dmem_n1025) );
NAND2_X1 MEM_stage_inst_dmem_U1190 ( .A1(MEM_stage_inst_dmem_ram_33), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n1026) );
NAND2_X1 MEM_stage_inst_dmem_U1189 ( .A1(MEM_stage_inst_dmem_n1024), .A2(MEM_stage_inst_dmem_n1023), .ZN(MEM_stage_inst_dmem_n1028) );
NAND2_X1 MEM_stage_inst_dmem_U1188 ( .A1(MEM_stage_inst_dmem_ram_353), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n1023) );
NAND2_X1 MEM_stage_inst_dmem_U1187 ( .A1(MEM_stage_inst_dmem_ram_577), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n1024) );
NOR2_X1 MEM_stage_inst_dmem_U1186 ( .A1(MEM_stage_inst_dmem_n1022), .A2(MEM_stage_inst_dmem_n1021), .ZN(MEM_stage_inst_dmem_n1030) );
NAND2_X1 MEM_stage_inst_dmem_U1185 ( .A1(MEM_stage_inst_dmem_n1020), .A2(MEM_stage_inst_dmem_n1019), .ZN(MEM_stage_inst_dmem_n1021) );
NAND2_X1 MEM_stage_inst_dmem_U1184 ( .A1(MEM_stage_inst_dmem_ram_305), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n1019) );
NAND2_X1 MEM_stage_inst_dmem_U1183 ( .A1(MEM_stage_inst_dmem_ram_49), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n1020) );
NAND2_X1 MEM_stage_inst_dmem_U1182 ( .A1(MEM_stage_inst_dmem_n1018), .A2(MEM_stage_inst_dmem_n1017), .ZN(MEM_stage_inst_dmem_n1022) );
NAND2_X1 MEM_stage_inst_dmem_U1181 ( .A1(MEM_stage_inst_dmem_ram_705), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n1017) );
NAND2_X1 MEM_stage_inst_dmem_U1180 ( .A1(MEM_stage_inst_dmem_ram_97), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n1018) );
NOR2_X1 MEM_stage_inst_dmem_U1179 ( .A1(MEM_stage_inst_dmem_n1016), .A2(MEM_stage_inst_dmem_n1015), .ZN(MEM_stage_inst_dmem_n1274) );
NOR2_X1 MEM_stage_inst_dmem_U1178 ( .A1(MEM_stage_inst_dmem_n1014), .A2(MEM_stage_inst_dmem_n8417), .ZN(MEM_stage_inst_dmem_n1015) );
NOR2_X1 MEM_stage_inst_dmem_U1177 ( .A1(MEM_stage_inst_dmem_n1013), .A2(MEM_stage_inst_dmem_n1012), .ZN(MEM_stage_inst_dmem_n1014) );
NAND2_X1 MEM_stage_inst_dmem_U1176 ( .A1(MEM_stage_inst_dmem_n1011), .A2(MEM_stage_inst_dmem_n1010), .ZN(MEM_stage_inst_dmem_n1012) );
NOR2_X1 MEM_stage_inst_dmem_U1175 ( .A1(MEM_stage_inst_dmem_n1009), .A2(MEM_stage_inst_dmem_n1008), .ZN(MEM_stage_inst_dmem_n1010) );
NAND2_X1 MEM_stage_inst_dmem_U1174 ( .A1(MEM_stage_inst_dmem_n1007), .A2(MEM_stage_inst_dmem_n1006), .ZN(MEM_stage_inst_dmem_n1008) );
NOR2_X1 MEM_stage_inst_dmem_U1173 ( .A1(MEM_stage_inst_dmem_n1005), .A2(MEM_stage_inst_dmem_n1004), .ZN(MEM_stage_inst_dmem_n1006) );
NAND2_X1 MEM_stage_inst_dmem_U1172 ( .A1(MEM_stage_inst_dmem_n1003), .A2(MEM_stage_inst_dmem_n1002), .ZN(MEM_stage_inst_dmem_n1004) );
NAND2_X1 MEM_stage_inst_dmem_U1171 ( .A1(MEM_stage_inst_dmem_ram_3569), .A2(MEM_stage_inst_dmem_n3170), .ZN(MEM_stage_inst_dmem_n1002) );
NAND2_X1 MEM_stage_inst_dmem_U1170 ( .A1(MEM_stage_inst_dmem_ram_4001), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n1003) );
NAND2_X1 MEM_stage_inst_dmem_U1169 ( .A1(MEM_stage_inst_dmem_n1001), .A2(MEM_stage_inst_dmem_n1000), .ZN(MEM_stage_inst_dmem_n1005) );
NAND2_X1 MEM_stage_inst_dmem_U1168 ( .A1(MEM_stage_inst_dmem_ram_3345), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n1000) );
NAND2_X1 MEM_stage_inst_dmem_U1167 ( .A1(MEM_stage_inst_dmem_ram_3457), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n1001) );
NOR2_X1 MEM_stage_inst_dmem_U1166 ( .A1(MEM_stage_inst_dmem_n999), .A2(MEM_stage_inst_dmem_n998), .ZN(MEM_stage_inst_dmem_n1007) );
NAND2_X1 MEM_stage_inst_dmem_U1165 ( .A1(MEM_stage_inst_dmem_n997), .A2(MEM_stage_inst_dmem_n996), .ZN(MEM_stage_inst_dmem_n998) );
NAND2_X1 MEM_stage_inst_dmem_U1164 ( .A1(MEM_stage_inst_dmem_ram_3121), .A2(MEM_stage_inst_dmem_n3103), .ZN(MEM_stage_inst_dmem_n996) );
NAND2_X1 MEM_stage_inst_dmem_U1163 ( .A1(MEM_stage_inst_dmem_ram_3073), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n997) );
NAND2_X1 MEM_stage_inst_dmem_U1162 ( .A1(MEM_stage_inst_dmem_n995), .A2(MEM_stage_inst_dmem_n994), .ZN(MEM_stage_inst_dmem_n999) );
NAND2_X1 MEM_stage_inst_dmem_U1161 ( .A1(MEM_stage_inst_dmem_ram_3953), .A2(MEM_stage_inst_dmem_n3099), .ZN(MEM_stage_inst_dmem_n994) );
NAND2_X1 MEM_stage_inst_dmem_U1160 ( .A1(MEM_stage_inst_dmem_ram_3681), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n995) );
NAND2_X1 MEM_stage_inst_dmem_U1159 ( .A1(MEM_stage_inst_dmem_n993), .A2(MEM_stage_inst_dmem_n992), .ZN(MEM_stage_inst_dmem_n1009) );
NOR2_X1 MEM_stage_inst_dmem_U1158 ( .A1(MEM_stage_inst_dmem_n991), .A2(MEM_stage_inst_dmem_n990), .ZN(MEM_stage_inst_dmem_n992) );
NAND2_X1 MEM_stage_inst_dmem_U1157 ( .A1(MEM_stage_inst_dmem_n989), .A2(MEM_stage_inst_dmem_n988), .ZN(MEM_stage_inst_dmem_n990) );
NAND2_X1 MEM_stage_inst_dmem_U1156 ( .A1(MEM_stage_inst_dmem_ram_3329), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n988) );
NAND2_X1 MEM_stage_inst_dmem_U1155 ( .A1(MEM_stage_inst_dmem_ram_3649), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n989) );
NAND2_X1 MEM_stage_inst_dmem_U1154 ( .A1(MEM_stage_inst_dmem_n987), .A2(MEM_stage_inst_dmem_n986), .ZN(MEM_stage_inst_dmem_n991) );
NAND2_X1 MEM_stage_inst_dmem_U1153 ( .A1(MEM_stage_inst_dmem_ram_3137), .A2(MEM_stage_inst_dmem_n3102), .ZN(MEM_stage_inst_dmem_n986) );
NAND2_X1 MEM_stage_inst_dmem_U1152 ( .A1(MEM_stage_inst_dmem_ram_3441), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n987) );
NOR2_X1 MEM_stage_inst_dmem_U1151 ( .A1(MEM_stage_inst_dmem_n985), .A2(MEM_stage_inst_dmem_n984), .ZN(MEM_stage_inst_dmem_n993) );
NAND2_X1 MEM_stage_inst_dmem_U1150 ( .A1(MEM_stage_inst_dmem_n983), .A2(MEM_stage_inst_dmem_n982), .ZN(MEM_stage_inst_dmem_n984) );
NAND2_X1 MEM_stage_inst_dmem_U1149 ( .A1(MEM_stage_inst_dmem_ram_3281), .A2(MEM_stage_inst_dmem_n3220), .ZN(MEM_stage_inst_dmem_n982) );
NAND2_X1 MEM_stage_inst_dmem_U1148 ( .A1(MEM_stage_inst_dmem_ram_3793), .A2(MEM_stage_inst_dmem_n3112), .ZN(MEM_stage_inst_dmem_n983) );
NAND2_X1 MEM_stage_inst_dmem_U1147 ( .A1(MEM_stage_inst_dmem_n981), .A2(MEM_stage_inst_dmem_n980), .ZN(MEM_stage_inst_dmem_n985) );
NAND2_X1 MEM_stage_inst_dmem_U1146 ( .A1(MEM_stage_inst_dmem_ram_3553), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n980) );
NAND2_X1 MEM_stage_inst_dmem_U1145 ( .A1(MEM_stage_inst_dmem_ram_3713), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n981) );
NOR2_X1 MEM_stage_inst_dmem_U1144 ( .A1(MEM_stage_inst_dmem_n979), .A2(MEM_stage_inst_dmem_n978), .ZN(MEM_stage_inst_dmem_n1011) );
NAND2_X1 MEM_stage_inst_dmem_U1143 ( .A1(MEM_stage_inst_dmem_n977), .A2(MEM_stage_inst_dmem_n976), .ZN(MEM_stage_inst_dmem_n978) );
NOR2_X1 MEM_stage_inst_dmem_U1142 ( .A1(MEM_stage_inst_dmem_n975), .A2(MEM_stage_inst_dmem_n974), .ZN(MEM_stage_inst_dmem_n976) );
NAND2_X1 MEM_stage_inst_dmem_U1141 ( .A1(MEM_stage_inst_dmem_n973), .A2(MEM_stage_inst_dmem_n972), .ZN(MEM_stage_inst_dmem_n974) );
NAND2_X1 MEM_stage_inst_dmem_U1140 ( .A1(MEM_stage_inst_dmem_ram_3489), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n972) );
NAND2_X1 MEM_stage_inst_dmem_U1139 ( .A1(MEM_stage_inst_dmem_ram_3745), .A2(MEM_stage_inst_dmem_n3155), .ZN(MEM_stage_inst_dmem_n973) );
NAND2_X1 MEM_stage_inst_dmem_U1138 ( .A1(MEM_stage_inst_dmem_n971), .A2(MEM_stage_inst_dmem_n970), .ZN(MEM_stage_inst_dmem_n975) );
NAND2_X1 MEM_stage_inst_dmem_U1137 ( .A1(MEM_stage_inst_dmem_ram_3153), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n970) );
NAND2_X1 MEM_stage_inst_dmem_U1136 ( .A1(MEM_stage_inst_dmem_ram_3665), .A2(MEM_stage_inst_dmem_n3140), .ZN(MEM_stage_inst_dmem_n971) );
NOR2_X1 MEM_stage_inst_dmem_U1135 ( .A1(MEM_stage_inst_dmem_n969), .A2(MEM_stage_inst_dmem_n968), .ZN(MEM_stage_inst_dmem_n977) );
NAND2_X1 MEM_stage_inst_dmem_U1134 ( .A1(MEM_stage_inst_dmem_n967), .A2(MEM_stage_inst_dmem_n966), .ZN(MEM_stage_inst_dmem_n968) );
NAND2_X1 MEM_stage_inst_dmem_U1133 ( .A1(MEM_stage_inst_dmem_ram_3265), .A2(MEM_stage_inst_dmem_n3082), .ZN(MEM_stage_inst_dmem_n966) );
NAND2_X1 MEM_stage_inst_dmem_U1132 ( .A1(MEM_stage_inst_dmem_ram_3201), .A2(MEM_stage_inst_dmem_n3130), .ZN(MEM_stage_inst_dmem_n967) );
NAND2_X1 MEM_stage_inst_dmem_U1131 ( .A1(MEM_stage_inst_dmem_n965), .A2(MEM_stage_inst_dmem_n964), .ZN(MEM_stage_inst_dmem_n969) );
NAND2_X1 MEM_stage_inst_dmem_U1130 ( .A1(MEM_stage_inst_dmem_ram_3889), .A2(MEM_stage_inst_dmem_n46), .ZN(MEM_stage_inst_dmem_n964) );
NAND2_X1 MEM_stage_inst_dmem_U1129 ( .A1(MEM_stage_inst_dmem_ram_3361), .A2(MEM_stage_inst_dmem_n3209), .ZN(MEM_stage_inst_dmem_n965) );
NAND2_X1 MEM_stage_inst_dmem_U1128 ( .A1(MEM_stage_inst_dmem_n963), .A2(MEM_stage_inst_dmem_n962), .ZN(MEM_stage_inst_dmem_n979) );
NOR2_X1 MEM_stage_inst_dmem_U1127 ( .A1(MEM_stage_inst_dmem_n961), .A2(MEM_stage_inst_dmem_n960), .ZN(MEM_stage_inst_dmem_n962) );
NAND2_X1 MEM_stage_inst_dmem_U1126 ( .A1(MEM_stage_inst_dmem_n959), .A2(MEM_stage_inst_dmem_n958), .ZN(MEM_stage_inst_dmem_n960) );
NAND2_X1 MEM_stage_inst_dmem_U1125 ( .A1(MEM_stage_inst_dmem_ram_3905), .A2(MEM_stage_inst_dmem_n3120), .ZN(MEM_stage_inst_dmem_n958) );
NAND2_X1 MEM_stage_inst_dmem_U1124 ( .A1(MEM_stage_inst_dmem_ram_3729), .A2(MEM_stage_inst_dmem_n3076), .ZN(MEM_stage_inst_dmem_n959) );
NAND2_X1 MEM_stage_inst_dmem_U1123 ( .A1(MEM_stage_inst_dmem_n957), .A2(MEM_stage_inst_dmem_n956), .ZN(MEM_stage_inst_dmem_n961) );
NAND2_X1 MEM_stage_inst_dmem_U1122 ( .A1(MEM_stage_inst_dmem_ram_3601), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n956) );
NAND2_X1 MEM_stage_inst_dmem_U1121 ( .A1(MEM_stage_inst_dmem_ram_3585), .A2(MEM_stage_inst_dmem_n3182), .ZN(MEM_stage_inst_dmem_n957) );
NOR2_X1 MEM_stage_inst_dmem_U1120 ( .A1(MEM_stage_inst_dmem_n955), .A2(MEM_stage_inst_dmem_n954), .ZN(MEM_stage_inst_dmem_n963) );
NAND2_X1 MEM_stage_inst_dmem_U1119 ( .A1(MEM_stage_inst_dmem_n953), .A2(MEM_stage_inst_dmem_n952), .ZN(MEM_stage_inst_dmem_n954) );
NAND2_X1 MEM_stage_inst_dmem_U1118 ( .A1(MEM_stage_inst_dmem_ram_3921), .A2(MEM_stage_inst_dmem_n3141), .ZN(MEM_stage_inst_dmem_n952) );
NAND2_X1 MEM_stage_inst_dmem_U1117 ( .A1(MEM_stage_inst_dmem_ram_4049), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n953) );
NAND2_X1 MEM_stage_inst_dmem_U1116 ( .A1(MEM_stage_inst_dmem_n951), .A2(MEM_stage_inst_dmem_n950), .ZN(MEM_stage_inst_dmem_n955) );
NAND2_X1 MEM_stage_inst_dmem_U1115 ( .A1(MEM_stage_inst_dmem_ram_4033), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n950) );
NAND2_X1 MEM_stage_inst_dmem_U1114 ( .A1(MEM_stage_inst_dmem_ram_3169), .A2(MEM_stage_inst_dmem_n3179), .ZN(MEM_stage_inst_dmem_n951) );
NAND2_X1 MEM_stage_inst_dmem_U1113 ( .A1(MEM_stage_inst_dmem_n949), .A2(MEM_stage_inst_dmem_n948), .ZN(MEM_stage_inst_dmem_n1013) );
NOR2_X1 MEM_stage_inst_dmem_U1112 ( .A1(MEM_stage_inst_dmem_n947), .A2(MEM_stage_inst_dmem_n946), .ZN(MEM_stage_inst_dmem_n948) );
NAND2_X1 MEM_stage_inst_dmem_U1111 ( .A1(MEM_stage_inst_dmem_n945), .A2(MEM_stage_inst_dmem_n944), .ZN(MEM_stage_inst_dmem_n946) );
NOR2_X1 MEM_stage_inst_dmem_U1110 ( .A1(MEM_stage_inst_dmem_n943), .A2(MEM_stage_inst_dmem_n942), .ZN(MEM_stage_inst_dmem_n944) );
NAND2_X1 MEM_stage_inst_dmem_U1109 ( .A1(MEM_stage_inst_dmem_n941), .A2(MEM_stage_inst_dmem_n940), .ZN(MEM_stage_inst_dmem_n942) );
NAND2_X1 MEM_stage_inst_dmem_U1108 ( .A1(MEM_stage_inst_dmem_ram_3505), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n940) );
NAND2_X1 MEM_stage_inst_dmem_U1107 ( .A1(MEM_stage_inst_dmem_ram_3249), .A2(MEM_stage_inst_dmem_n8434), .ZN(MEM_stage_inst_dmem_n941) );
NAND2_X1 MEM_stage_inst_dmem_U1106 ( .A1(MEM_stage_inst_dmem_n939), .A2(MEM_stage_inst_dmem_n938), .ZN(MEM_stage_inst_dmem_n943) );
NAND2_X1 MEM_stage_inst_dmem_U1105 ( .A1(MEM_stage_inst_dmem_ram_3393), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n938) );
NAND2_X1 MEM_stage_inst_dmem_U1104 ( .A1(MEM_stage_inst_dmem_ram_3825), .A2(MEM_stage_inst_dmem_n3202), .ZN(MEM_stage_inst_dmem_n939) );
NOR2_X1 MEM_stage_inst_dmem_U1103 ( .A1(MEM_stage_inst_dmem_n937), .A2(MEM_stage_inst_dmem_n936), .ZN(MEM_stage_inst_dmem_n945) );
NAND2_X1 MEM_stage_inst_dmem_U1102 ( .A1(MEM_stage_inst_dmem_n935), .A2(MEM_stage_inst_dmem_n934), .ZN(MEM_stage_inst_dmem_n936) );
NAND2_X1 MEM_stage_inst_dmem_U1101 ( .A1(MEM_stage_inst_dmem_ram_3937), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n934) );
NAND2_X1 MEM_stage_inst_dmem_U1100 ( .A1(MEM_stage_inst_dmem_ram_4017), .A2(MEM_stage_inst_dmem_n3163), .ZN(MEM_stage_inst_dmem_n935) );
NAND2_X1 MEM_stage_inst_dmem_U1099 ( .A1(MEM_stage_inst_dmem_n933), .A2(MEM_stage_inst_dmem_n932), .ZN(MEM_stage_inst_dmem_n937) );
NAND2_X1 MEM_stage_inst_dmem_U1098 ( .A1(MEM_stage_inst_dmem_ram_3297), .A2(MEM_stage_inst_dmem_n3152), .ZN(MEM_stage_inst_dmem_n932) );
NAND2_X1 MEM_stage_inst_dmem_U1097 ( .A1(MEM_stage_inst_dmem_ram_3217), .A2(MEM_stage_inst_dmem_n44), .ZN(MEM_stage_inst_dmem_n933) );
NAND2_X1 MEM_stage_inst_dmem_U1096 ( .A1(MEM_stage_inst_dmem_n931), .A2(MEM_stage_inst_dmem_n930), .ZN(MEM_stage_inst_dmem_n947) );
NOR2_X1 MEM_stage_inst_dmem_U1095 ( .A1(MEM_stage_inst_dmem_n929), .A2(MEM_stage_inst_dmem_n928), .ZN(MEM_stage_inst_dmem_n930) );
NAND2_X1 MEM_stage_inst_dmem_U1094 ( .A1(MEM_stage_inst_dmem_n927), .A2(MEM_stage_inst_dmem_n926), .ZN(MEM_stage_inst_dmem_n928) );
NAND2_X1 MEM_stage_inst_dmem_U1093 ( .A1(MEM_stage_inst_dmem_ram_3985), .A2(MEM_stage_inst_dmem_n3073), .ZN(MEM_stage_inst_dmem_n926) );
NAND2_X1 MEM_stage_inst_dmem_U1092 ( .A1(MEM_stage_inst_dmem_ram_3697), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n927) );
NAND2_X1 MEM_stage_inst_dmem_U1091 ( .A1(MEM_stage_inst_dmem_n925), .A2(MEM_stage_inst_dmem_n924), .ZN(MEM_stage_inst_dmem_n929) );
NAND2_X1 MEM_stage_inst_dmem_U1090 ( .A1(MEM_stage_inst_dmem_ram_3313), .A2(MEM_stage_inst_dmem_n39), .ZN(MEM_stage_inst_dmem_n924) );
NAND2_X1 MEM_stage_inst_dmem_U1089 ( .A1(MEM_stage_inst_dmem_ram_3873), .A2(MEM_stage_inst_dmem_n3137), .ZN(MEM_stage_inst_dmem_n925) );
NOR2_X1 MEM_stage_inst_dmem_U1088 ( .A1(MEM_stage_inst_dmem_n923), .A2(MEM_stage_inst_dmem_n922), .ZN(MEM_stage_inst_dmem_n931) );
NAND2_X1 MEM_stage_inst_dmem_U1087 ( .A1(MEM_stage_inst_dmem_n921), .A2(MEM_stage_inst_dmem_n920), .ZN(MEM_stage_inst_dmem_n922) );
NAND2_X1 MEM_stage_inst_dmem_U1086 ( .A1(MEM_stage_inst_dmem_ram_3089), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n920) );
NAND2_X1 MEM_stage_inst_dmem_U1085 ( .A1(MEM_stage_inst_dmem_ram_3409), .A2(MEM_stage_inst_dmem_n3216), .ZN(MEM_stage_inst_dmem_n921) );
NAND2_X1 MEM_stage_inst_dmem_U1084 ( .A1(MEM_stage_inst_dmem_n919), .A2(MEM_stage_inst_dmem_n918), .ZN(MEM_stage_inst_dmem_n923) );
NAND2_X1 MEM_stage_inst_dmem_U1083 ( .A1(MEM_stage_inst_dmem_ram_3425), .A2(MEM_stage_inst_dmem_n3217), .ZN(MEM_stage_inst_dmem_n918) );
NAND2_X1 MEM_stage_inst_dmem_U1082 ( .A1(MEM_stage_inst_dmem_ram_3633), .A2(MEM_stage_inst_dmem_n3085), .ZN(MEM_stage_inst_dmem_n919) );
NOR2_X1 MEM_stage_inst_dmem_U1081 ( .A1(MEM_stage_inst_dmem_n917), .A2(MEM_stage_inst_dmem_n916), .ZN(MEM_stage_inst_dmem_n949) );
NAND2_X1 MEM_stage_inst_dmem_U1080 ( .A1(MEM_stage_inst_dmem_n915), .A2(MEM_stage_inst_dmem_n914), .ZN(MEM_stage_inst_dmem_n916) );
NOR2_X1 MEM_stage_inst_dmem_U1079 ( .A1(MEM_stage_inst_dmem_n913), .A2(MEM_stage_inst_dmem_n912), .ZN(MEM_stage_inst_dmem_n914) );
NAND2_X1 MEM_stage_inst_dmem_U1078 ( .A1(MEM_stage_inst_dmem_n911), .A2(MEM_stage_inst_dmem_n910), .ZN(MEM_stage_inst_dmem_n912) );
NAND2_X1 MEM_stage_inst_dmem_U1077 ( .A1(MEM_stage_inst_dmem_ram_3473), .A2(MEM_stage_inst_dmem_n3160), .ZN(MEM_stage_inst_dmem_n910) );
NAND2_X1 MEM_stage_inst_dmem_U1076 ( .A1(MEM_stage_inst_dmem_ram_3537), .A2(MEM_stage_inst_dmem_n3174), .ZN(MEM_stage_inst_dmem_n911) );
NAND2_X1 MEM_stage_inst_dmem_U1075 ( .A1(MEM_stage_inst_dmem_n909), .A2(MEM_stage_inst_dmem_n908), .ZN(MEM_stage_inst_dmem_n913) );
NAND2_X1 MEM_stage_inst_dmem_U1074 ( .A1(MEM_stage_inst_dmem_ram_4065), .A2(MEM_stage_inst_dmem_n3113), .ZN(MEM_stage_inst_dmem_n908) );
NAND2_X1 MEM_stage_inst_dmem_U1073 ( .A1(MEM_stage_inst_dmem_ram_3809), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n909) );
NOR2_X1 MEM_stage_inst_dmem_U1072 ( .A1(MEM_stage_inst_dmem_n907), .A2(MEM_stage_inst_dmem_n906), .ZN(MEM_stage_inst_dmem_n915) );
NAND2_X1 MEM_stage_inst_dmem_U1071 ( .A1(MEM_stage_inst_dmem_n905), .A2(MEM_stage_inst_dmem_n904), .ZN(MEM_stage_inst_dmem_n906) );
NAND2_X1 MEM_stage_inst_dmem_U1070 ( .A1(MEM_stage_inst_dmem_ram_3969), .A2(MEM_stage_inst_dmem_n3123), .ZN(MEM_stage_inst_dmem_n904) );
NAND2_X1 MEM_stage_inst_dmem_U1069 ( .A1(MEM_stage_inst_dmem_ram_3105), .A2(MEM_stage_inst_dmem_n3092), .ZN(MEM_stage_inst_dmem_n905) );
NAND2_X1 MEM_stage_inst_dmem_U1068 ( .A1(MEM_stage_inst_dmem_n903), .A2(MEM_stage_inst_dmem_n902), .ZN(MEM_stage_inst_dmem_n907) );
NAND2_X1 MEM_stage_inst_dmem_U1067 ( .A1(MEM_stage_inst_dmem_ram_3185), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n902) );
NAND2_X1 MEM_stage_inst_dmem_U1066 ( .A1(MEM_stage_inst_dmem_ram_3233), .A2(MEM_stage_inst_dmem_n3081), .ZN(MEM_stage_inst_dmem_n903) );
NAND2_X1 MEM_stage_inst_dmem_U1065 ( .A1(MEM_stage_inst_dmem_n901), .A2(MEM_stage_inst_dmem_n900), .ZN(MEM_stage_inst_dmem_n917) );
NOR2_X1 MEM_stage_inst_dmem_U1064 ( .A1(MEM_stage_inst_dmem_n899), .A2(MEM_stage_inst_dmem_n898), .ZN(MEM_stage_inst_dmem_n900) );
NAND2_X1 MEM_stage_inst_dmem_U1063 ( .A1(MEM_stage_inst_dmem_n897), .A2(MEM_stage_inst_dmem_n896), .ZN(MEM_stage_inst_dmem_n898) );
NAND2_X1 MEM_stage_inst_dmem_U1062 ( .A1(MEM_stage_inst_dmem_ram_3377), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n896) );
NAND2_X1 MEM_stage_inst_dmem_U1061 ( .A1(MEM_stage_inst_dmem_ram_3761), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n897) );
NAND2_X1 MEM_stage_inst_dmem_U1060 ( .A1(MEM_stage_inst_dmem_n895), .A2(MEM_stage_inst_dmem_n894), .ZN(MEM_stage_inst_dmem_n899) );
NAND2_X1 MEM_stage_inst_dmem_U1059 ( .A1(MEM_stage_inst_dmem_ram_4081), .A2(MEM_stage_inst_dmem_n3199), .ZN(MEM_stage_inst_dmem_n894) );
NAND2_X1 MEM_stage_inst_dmem_U1058 ( .A1(MEM_stage_inst_dmem_ram_3857), .A2(MEM_stage_inst_dmem_n3191), .ZN(MEM_stage_inst_dmem_n895) );
NOR2_X1 MEM_stage_inst_dmem_U1057 ( .A1(MEM_stage_inst_dmem_n893), .A2(MEM_stage_inst_dmem_n892), .ZN(MEM_stage_inst_dmem_n901) );
NAND2_X1 MEM_stage_inst_dmem_U1056 ( .A1(MEM_stage_inst_dmem_n891), .A2(MEM_stage_inst_dmem_n890), .ZN(MEM_stage_inst_dmem_n892) );
NAND2_X1 MEM_stage_inst_dmem_U1055 ( .A1(MEM_stage_inst_dmem_ram_3617), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n890) );
NAND2_X1 MEM_stage_inst_dmem_U1054 ( .A1(MEM_stage_inst_dmem_ram_3521), .A2(MEM_stage_inst_dmem_n3173), .ZN(MEM_stage_inst_dmem_n891) );
NAND2_X1 MEM_stage_inst_dmem_U1053 ( .A1(MEM_stage_inst_dmem_n889), .A2(MEM_stage_inst_dmem_n888), .ZN(MEM_stage_inst_dmem_n893) );
NAND2_X1 MEM_stage_inst_dmem_U1052 ( .A1(MEM_stage_inst_dmem_ram_3841), .A2(MEM_stage_inst_dmem_n8472), .ZN(MEM_stage_inst_dmem_n888) );
NAND2_X1 MEM_stage_inst_dmem_U1051 ( .A1(MEM_stage_inst_dmem_ram_3777), .A2(MEM_stage_inst_dmem_n3192), .ZN(MEM_stage_inst_dmem_n889) );
NOR2_X1 MEM_stage_inst_dmem_U1050 ( .A1(MEM_stage_inst_dmem_n887), .A2(MEM_stage_inst_dmem_n8152), .ZN(MEM_stage_inst_dmem_n1016) );
NOR2_X1 MEM_stage_inst_dmem_U1049 ( .A1(MEM_stage_inst_dmem_n886), .A2(MEM_stage_inst_dmem_n885), .ZN(MEM_stage_inst_dmem_n887) );
NAND2_X1 MEM_stage_inst_dmem_U1048 ( .A1(MEM_stage_inst_dmem_n884), .A2(MEM_stage_inst_dmem_n883), .ZN(MEM_stage_inst_dmem_n885) );
NOR2_X1 MEM_stage_inst_dmem_U1047 ( .A1(MEM_stage_inst_dmem_n882), .A2(MEM_stage_inst_dmem_n881), .ZN(MEM_stage_inst_dmem_n883) );
NAND2_X1 MEM_stage_inst_dmem_U1046 ( .A1(MEM_stage_inst_dmem_n880), .A2(MEM_stage_inst_dmem_n879), .ZN(MEM_stage_inst_dmem_n881) );
NOR2_X1 MEM_stage_inst_dmem_U1045 ( .A1(MEM_stage_inst_dmem_n878), .A2(MEM_stage_inst_dmem_n877), .ZN(MEM_stage_inst_dmem_n879) );
NAND2_X1 MEM_stage_inst_dmem_U1044 ( .A1(MEM_stage_inst_dmem_n876), .A2(MEM_stage_inst_dmem_n875), .ZN(MEM_stage_inst_dmem_n877) );
NAND2_X1 MEM_stage_inst_dmem_U1043 ( .A1(MEM_stage_inst_dmem_ram_1313), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n875) );
NAND2_X1 MEM_stage_inst_dmem_U1042 ( .A1(MEM_stage_inst_dmem_ram_1361), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n876) );
NAND2_X1 MEM_stage_inst_dmem_U1041 ( .A1(MEM_stage_inst_dmem_n874), .A2(MEM_stage_inst_dmem_n873), .ZN(MEM_stage_inst_dmem_n878) );
NAND2_X1 MEM_stage_inst_dmem_U1040 ( .A1(MEM_stage_inst_dmem_ram_1521), .A2(MEM_stage_inst_dmem_n8535), .ZN(MEM_stage_inst_dmem_n873) );
NAND2_X1 MEM_stage_inst_dmem_U1039 ( .A1(MEM_stage_inst_dmem_ram_1121), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n874) );
NOR2_X1 MEM_stage_inst_dmem_U1038 ( .A1(MEM_stage_inst_dmem_n872), .A2(MEM_stage_inst_dmem_n871), .ZN(MEM_stage_inst_dmem_n880) );
NAND2_X1 MEM_stage_inst_dmem_U1037 ( .A1(MEM_stage_inst_dmem_n870), .A2(MEM_stage_inst_dmem_n869), .ZN(MEM_stage_inst_dmem_n871) );
NAND2_X1 MEM_stage_inst_dmem_U1036 ( .A1(MEM_stage_inst_dmem_ram_1697), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n869) );
NAND2_X1 MEM_stage_inst_dmem_U1035 ( .A1(MEM_stage_inst_dmem_ram_1025), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n870) );
NAND2_X1 MEM_stage_inst_dmem_U1034 ( .A1(MEM_stage_inst_dmem_n868), .A2(MEM_stage_inst_dmem_n867), .ZN(MEM_stage_inst_dmem_n872) );
NAND2_X1 MEM_stage_inst_dmem_U1033 ( .A1(MEM_stage_inst_dmem_ram_1297), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n867) );
NAND2_X1 MEM_stage_inst_dmem_U1032 ( .A1(MEM_stage_inst_dmem_ram_1473), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n868) );
NAND2_X1 MEM_stage_inst_dmem_U1031 ( .A1(MEM_stage_inst_dmem_n866), .A2(MEM_stage_inst_dmem_n865), .ZN(MEM_stage_inst_dmem_n882) );
NOR2_X1 MEM_stage_inst_dmem_U1030 ( .A1(MEM_stage_inst_dmem_n864), .A2(MEM_stage_inst_dmem_n863), .ZN(MEM_stage_inst_dmem_n865) );
NAND2_X1 MEM_stage_inst_dmem_U1029 ( .A1(MEM_stage_inst_dmem_n862), .A2(MEM_stage_inst_dmem_n861), .ZN(MEM_stage_inst_dmem_n863) );
NAND2_X1 MEM_stage_inst_dmem_U1028 ( .A1(MEM_stage_inst_dmem_ram_1105), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n861) );
NAND2_X1 MEM_stage_inst_dmem_U1027 ( .A1(MEM_stage_inst_dmem_ram_1681), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n862) );
NAND2_X1 MEM_stage_inst_dmem_U1026 ( .A1(MEM_stage_inst_dmem_n860), .A2(MEM_stage_inst_dmem_n859), .ZN(MEM_stage_inst_dmem_n864) );
NAND2_X1 MEM_stage_inst_dmem_U1025 ( .A1(MEM_stage_inst_dmem_ram_1713), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n859) );
NAND2_X1 MEM_stage_inst_dmem_U1024 ( .A1(MEM_stage_inst_dmem_ram_1953), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n860) );
NOR2_X1 MEM_stage_inst_dmem_U1023 ( .A1(MEM_stage_inst_dmem_n858), .A2(MEM_stage_inst_dmem_n857), .ZN(MEM_stage_inst_dmem_n866) );
NAND2_X1 MEM_stage_inst_dmem_U1022 ( .A1(MEM_stage_inst_dmem_n856), .A2(MEM_stage_inst_dmem_n855), .ZN(MEM_stage_inst_dmem_n857) );
NAND2_X1 MEM_stage_inst_dmem_U1021 ( .A1(MEM_stage_inst_dmem_ram_1825), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n855) );
NAND2_X1 MEM_stage_inst_dmem_U1020 ( .A1(MEM_stage_inst_dmem_ram_1393), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n856) );
NAND2_X1 MEM_stage_inst_dmem_U1019 ( .A1(MEM_stage_inst_dmem_n854), .A2(MEM_stage_inst_dmem_n853), .ZN(MEM_stage_inst_dmem_n858) );
NAND2_X1 MEM_stage_inst_dmem_U1018 ( .A1(MEM_stage_inst_dmem_ram_2033), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n853) );
NAND2_X1 MEM_stage_inst_dmem_U1017 ( .A1(MEM_stage_inst_dmem_ram_1201), .A2(MEM_stage_inst_dmem_n55), .ZN(MEM_stage_inst_dmem_n854) );
NOR2_X1 MEM_stage_inst_dmem_U1016 ( .A1(MEM_stage_inst_dmem_n852), .A2(MEM_stage_inst_dmem_n851), .ZN(MEM_stage_inst_dmem_n884) );
NAND2_X1 MEM_stage_inst_dmem_U1015 ( .A1(MEM_stage_inst_dmem_n850), .A2(MEM_stage_inst_dmem_n849), .ZN(MEM_stage_inst_dmem_n851) );
NOR2_X1 MEM_stage_inst_dmem_U1014 ( .A1(MEM_stage_inst_dmem_n848), .A2(MEM_stage_inst_dmem_n847), .ZN(MEM_stage_inst_dmem_n849) );
NAND2_X1 MEM_stage_inst_dmem_U1013 ( .A1(MEM_stage_inst_dmem_n846), .A2(MEM_stage_inst_dmem_n845), .ZN(MEM_stage_inst_dmem_n847) );
NAND2_X1 MEM_stage_inst_dmem_U1012 ( .A1(MEM_stage_inst_dmem_ram_1793), .A2(MEM_stage_inst_dmem_n37), .ZN(MEM_stage_inst_dmem_n845) );
NAND2_X1 MEM_stage_inst_dmem_U1011 ( .A1(MEM_stage_inst_dmem_ram_1185), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n846) );
NAND2_X1 MEM_stage_inst_dmem_U1010 ( .A1(MEM_stage_inst_dmem_n844), .A2(MEM_stage_inst_dmem_n843), .ZN(MEM_stage_inst_dmem_n848) );
NAND2_X1 MEM_stage_inst_dmem_U1009 ( .A1(MEM_stage_inst_dmem_ram_1873), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n843) );
NAND2_X1 MEM_stage_inst_dmem_U1008 ( .A1(MEM_stage_inst_dmem_ram_1969), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n844) );
NOR2_X1 MEM_stage_inst_dmem_U1007 ( .A1(MEM_stage_inst_dmem_n842), .A2(MEM_stage_inst_dmem_n841), .ZN(MEM_stage_inst_dmem_n850) );
NAND2_X1 MEM_stage_inst_dmem_U1006 ( .A1(MEM_stage_inst_dmem_n840), .A2(MEM_stage_inst_dmem_n839), .ZN(MEM_stage_inst_dmem_n841) );
NAND2_X1 MEM_stage_inst_dmem_U1005 ( .A1(MEM_stage_inst_dmem_ram_1249), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n839) );
NAND2_X1 MEM_stage_inst_dmem_U1004 ( .A1(MEM_stage_inst_dmem_ram_1425), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n840) );
NAND2_X1 MEM_stage_inst_dmem_U1003 ( .A1(MEM_stage_inst_dmem_n838), .A2(MEM_stage_inst_dmem_n837), .ZN(MEM_stage_inst_dmem_n842) );
NAND2_X1 MEM_stage_inst_dmem_U1002 ( .A1(MEM_stage_inst_dmem_ram_1457), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n837) );
NAND2_X1 MEM_stage_inst_dmem_U1001 ( .A1(MEM_stage_inst_dmem_ram_1585), .A2(MEM_stage_inst_dmem_n41), .ZN(MEM_stage_inst_dmem_n838) );
NAND2_X1 MEM_stage_inst_dmem_U1000 ( .A1(MEM_stage_inst_dmem_n836), .A2(MEM_stage_inst_dmem_n835), .ZN(MEM_stage_inst_dmem_n852) );
NOR2_X1 MEM_stage_inst_dmem_U999 ( .A1(MEM_stage_inst_dmem_n834), .A2(MEM_stage_inst_dmem_n833), .ZN(MEM_stage_inst_dmem_n835) );
NAND2_X1 MEM_stage_inst_dmem_U998 ( .A1(MEM_stage_inst_dmem_n832), .A2(MEM_stage_inst_dmem_n831), .ZN(MEM_stage_inst_dmem_n833) );
NAND2_X1 MEM_stage_inst_dmem_U997 ( .A1(MEM_stage_inst_dmem_ram_1889), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n831) );
NAND2_X1 MEM_stage_inst_dmem_U996 ( .A1(MEM_stage_inst_dmem_ram_1553), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n832) );
NAND2_X1 MEM_stage_inst_dmem_U995 ( .A1(MEM_stage_inst_dmem_n830), .A2(MEM_stage_inst_dmem_n829), .ZN(MEM_stage_inst_dmem_n834) );
NAND2_X1 MEM_stage_inst_dmem_U994 ( .A1(MEM_stage_inst_dmem_ram_1633), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n829) );
NAND2_X1 MEM_stage_inst_dmem_U993 ( .A1(MEM_stage_inst_dmem_ram_1809), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n830) );
NOR2_X1 MEM_stage_inst_dmem_U992 ( .A1(MEM_stage_inst_dmem_n828), .A2(MEM_stage_inst_dmem_n827), .ZN(MEM_stage_inst_dmem_n836) );
NAND2_X1 MEM_stage_inst_dmem_U991 ( .A1(MEM_stage_inst_dmem_n826), .A2(MEM_stage_inst_dmem_n825), .ZN(MEM_stage_inst_dmem_n827) );
NAND2_X1 MEM_stage_inst_dmem_U990 ( .A1(MEM_stage_inst_dmem_ram_1937), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n825) );
NAND2_X1 MEM_stage_inst_dmem_U989 ( .A1(MEM_stage_inst_dmem_ram_1921), .A2(MEM_stage_inst_dmem_n72), .ZN(MEM_stage_inst_dmem_n826) );
NAND2_X1 MEM_stage_inst_dmem_U988 ( .A1(MEM_stage_inst_dmem_n824), .A2(MEM_stage_inst_dmem_n823), .ZN(MEM_stage_inst_dmem_n828) );
NAND2_X1 MEM_stage_inst_dmem_U987 ( .A1(MEM_stage_inst_dmem_ram_1041), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n823) );
NAND2_X1 MEM_stage_inst_dmem_U986 ( .A1(MEM_stage_inst_dmem_ram_1649), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n824) );
NAND2_X1 MEM_stage_inst_dmem_U985 ( .A1(MEM_stage_inst_dmem_n822), .A2(MEM_stage_inst_dmem_n821), .ZN(MEM_stage_inst_dmem_n886) );
NOR2_X1 MEM_stage_inst_dmem_U984 ( .A1(MEM_stage_inst_dmem_n820), .A2(MEM_stage_inst_dmem_n819), .ZN(MEM_stage_inst_dmem_n821) );
NAND2_X1 MEM_stage_inst_dmem_U983 ( .A1(MEM_stage_inst_dmem_n818), .A2(MEM_stage_inst_dmem_n817), .ZN(MEM_stage_inst_dmem_n819) );
NOR2_X1 MEM_stage_inst_dmem_U982 ( .A1(MEM_stage_inst_dmem_n816), .A2(MEM_stage_inst_dmem_n815), .ZN(MEM_stage_inst_dmem_n817) );
NAND2_X1 MEM_stage_inst_dmem_U981 ( .A1(MEM_stage_inst_dmem_n814), .A2(MEM_stage_inst_dmem_n813), .ZN(MEM_stage_inst_dmem_n815) );
NAND2_X1 MEM_stage_inst_dmem_U980 ( .A1(MEM_stage_inst_dmem_ram_1857), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n813) );
NAND2_X1 MEM_stage_inst_dmem_U979 ( .A1(MEM_stage_inst_dmem_ram_1265), .A2(MEM_stage_inst_dmem_n39), .ZN(MEM_stage_inst_dmem_n814) );
NAND2_X1 MEM_stage_inst_dmem_U978 ( .A1(MEM_stage_inst_dmem_n812), .A2(MEM_stage_inst_dmem_n811), .ZN(MEM_stage_inst_dmem_n816) );
NAND2_X1 MEM_stage_inst_dmem_U977 ( .A1(MEM_stage_inst_dmem_ram_1985), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n811) );
NAND2_X1 MEM_stage_inst_dmem_U976 ( .A1(MEM_stage_inst_dmem_ram_1761), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n812) );
NOR2_X1 MEM_stage_inst_dmem_U975 ( .A1(MEM_stage_inst_dmem_n810), .A2(MEM_stage_inst_dmem_n809), .ZN(MEM_stage_inst_dmem_n818) );
NAND2_X1 MEM_stage_inst_dmem_U974 ( .A1(MEM_stage_inst_dmem_n808), .A2(MEM_stage_inst_dmem_n807), .ZN(MEM_stage_inst_dmem_n809) );
NAND2_X1 MEM_stage_inst_dmem_U973 ( .A1(MEM_stage_inst_dmem_ram_1905), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n807) );
NAND2_X1 MEM_stage_inst_dmem_U972 ( .A1(MEM_stage_inst_dmem_ram_1777), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n808) );
NAND2_X1 MEM_stage_inst_dmem_U971 ( .A1(MEM_stage_inst_dmem_n806), .A2(MEM_stage_inst_dmem_n805), .ZN(MEM_stage_inst_dmem_n810) );
NAND2_X1 MEM_stage_inst_dmem_U970 ( .A1(MEM_stage_inst_dmem_ram_2017), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n805) );
NAND2_X1 MEM_stage_inst_dmem_U969 ( .A1(MEM_stage_inst_dmem_ram_1569), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n806) );
NAND2_X1 MEM_stage_inst_dmem_U968 ( .A1(MEM_stage_inst_dmem_n804), .A2(MEM_stage_inst_dmem_n803), .ZN(MEM_stage_inst_dmem_n820) );
NOR2_X1 MEM_stage_inst_dmem_U967 ( .A1(MEM_stage_inst_dmem_n802), .A2(MEM_stage_inst_dmem_n801), .ZN(MEM_stage_inst_dmem_n803) );
NAND2_X1 MEM_stage_inst_dmem_U966 ( .A1(MEM_stage_inst_dmem_n800), .A2(MEM_stage_inst_dmem_n799), .ZN(MEM_stage_inst_dmem_n801) );
NAND2_X1 MEM_stage_inst_dmem_U965 ( .A1(MEM_stage_inst_dmem_ram_1841), .A2(MEM_stage_inst_dmem_n46), .ZN(MEM_stage_inst_dmem_n799) );
NAND2_X1 MEM_stage_inst_dmem_U964 ( .A1(MEM_stage_inst_dmem_ram_1233), .A2(MEM_stage_inst_dmem_n51), .ZN(MEM_stage_inst_dmem_n800) );
NAND2_X1 MEM_stage_inst_dmem_U963 ( .A1(MEM_stage_inst_dmem_n798), .A2(MEM_stage_inst_dmem_n797), .ZN(MEM_stage_inst_dmem_n802) );
NAND2_X1 MEM_stage_inst_dmem_U962 ( .A1(MEM_stage_inst_dmem_ram_1345), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n797) );
NAND2_X1 MEM_stage_inst_dmem_U961 ( .A1(MEM_stage_inst_dmem_ram_1505), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n798) );
NOR2_X1 MEM_stage_inst_dmem_U960 ( .A1(MEM_stage_inst_dmem_n796), .A2(MEM_stage_inst_dmem_n795), .ZN(MEM_stage_inst_dmem_n804) );
NAND2_X1 MEM_stage_inst_dmem_U959 ( .A1(MEM_stage_inst_dmem_n794), .A2(MEM_stage_inst_dmem_n793), .ZN(MEM_stage_inst_dmem_n795) );
NAND2_X1 MEM_stage_inst_dmem_U958 ( .A1(MEM_stage_inst_dmem_ram_2001), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n793) );
NAND2_X1 MEM_stage_inst_dmem_U957 ( .A1(MEM_stage_inst_dmem_ram_1169), .A2(MEM_stage_inst_dmem_n44), .ZN(MEM_stage_inst_dmem_n794) );
NAND2_X1 MEM_stage_inst_dmem_U956 ( .A1(MEM_stage_inst_dmem_n792), .A2(MEM_stage_inst_dmem_n791), .ZN(MEM_stage_inst_dmem_n796) );
NAND2_X1 MEM_stage_inst_dmem_U955 ( .A1(MEM_stage_inst_dmem_ram_1057), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n791) );
NAND2_X1 MEM_stage_inst_dmem_U954 ( .A1(MEM_stage_inst_dmem_ram_1409), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n792) );
NOR2_X1 MEM_stage_inst_dmem_U953 ( .A1(MEM_stage_inst_dmem_n790), .A2(MEM_stage_inst_dmem_n789), .ZN(MEM_stage_inst_dmem_n822) );
NAND2_X1 MEM_stage_inst_dmem_U952 ( .A1(MEM_stage_inst_dmem_n788), .A2(MEM_stage_inst_dmem_n787), .ZN(MEM_stage_inst_dmem_n789) );
NOR2_X1 MEM_stage_inst_dmem_U951 ( .A1(MEM_stage_inst_dmem_n786), .A2(MEM_stage_inst_dmem_n785), .ZN(MEM_stage_inst_dmem_n787) );
NAND2_X1 MEM_stage_inst_dmem_U950 ( .A1(MEM_stage_inst_dmem_n784), .A2(MEM_stage_inst_dmem_n783), .ZN(MEM_stage_inst_dmem_n785) );
NAND2_X1 MEM_stage_inst_dmem_U949 ( .A1(MEM_stage_inst_dmem_ram_1073), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n783) );
NAND2_X1 MEM_stage_inst_dmem_U948 ( .A1(MEM_stage_inst_dmem_ram_1489), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n784) );
NAND2_X1 MEM_stage_inst_dmem_U947 ( .A1(MEM_stage_inst_dmem_n782), .A2(MEM_stage_inst_dmem_n781), .ZN(MEM_stage_inst_dmem_n786) );
NAND2_X1 MEM_stage_inst_dmem_U946 ( .A1(MEM_stage_inst_dmem_ram_1377), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n781) );
NAND2_X1 MEM_stage_inst_dmem_U945 ( .A1(MEM_stage_inst_dmem_ram_1537), .A2(MEM_stage_inst_dmem_n71), .ZN(MEM_stage_inst_dmem_n782) );
NOR2_X1 MEM_stage_inst_dmem_U944 ( .A1(MEM_stage_inst_dmem_n780), .A2(MEM_stage_inst_dmem_n779), .ZN(MEM_stage_inst_dmem_n788) );
NAND2_X1 MEM_stage_inst_dmem_U943 ( .A1(MEM_stage_inst_dmem_n778), .A2(MEM_stage_inst_dmem_n777), .ZN(MEM_stage_inst_dmem_n779) );
NAND2_X1 MEM_stage_inst_dmem_U942 ( .A1(MEM_stage_inst_dmem_ram_1329), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n777) );
NAND2_X1 MEM_stage_inst_dmem_U941 ( .A1(MEM_stage_inst_dmem_ram_1281), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n778) );
NAND2_X1 MEM_stage_inst_dmem_U940 ( .A1(MEM_stage_inst_dmem_n776), .A2(MEM_stage_inst_dmem_n775), .ZN(MEM_stage_inst_dmem_n780) );
NAND2_X1 MEM_stage_inst_dmem_U939 ( .A1(MEM_stage_inst_dmem_ram_1153), .A2(MEM_stage_inst_dmem_n61), .ZN(MEM_stage_inst_dmem_n775) );
NAND2_X1 MEM_stage_inst_dmem_U938 ( .A1(MEM_stage_inst_dmem_ram_1617), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n776) );
NAND2_X1 MEM_stage_inst_dmem_U937 ( .A1(MEM_stage_inst_dmem_n774), .A2(MEM_stage_inst_dmem_n773), .ZN(MEM_stage_inst_dmem_n790) );
NOR2_X1 MEM_stage_inst_dmem_U936 ( .A1(MEM_stage_inst_dmem_n772), .A2(MEM_stage_inst_dmem_n771), .ZN(MEM_stage_inst_dmem_n773) );
NAND2_X1 MEM_stage_inst_dmem_U935 ( .A1(MEM_stage_inst_dmem_n770), .A2(MEM_stage_inst_dmem_n769), .ZN(MEM_stage_inst_dmem_n771) );
NAND2_X1 MEM_stage_inst_dmem_U934 ( .A1(MEM_stage_inst_dmem_ram_1217), .A2(MEM_stage_inst_dmem_n36), .ZN(MEM_stage_inst_dmem_n769) );
NAND2_X1 MEM_stage_inst_dmem_U933 ( .A1(MEM_stage_inst_dmem_ram_1089), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n770) );
NAND2_X1 MEM_stage_inst_dmem_U932 ( .A1(MEM_stage_inst_dmem_n768), .A2(MEM_stage_inst_dmem_n767), .ZN(MEM_stage_inst_dmem_n772) );
NAND2_X1 MEM_stage_inst_dmem_U931 ( .A1(MEM_stage_inst_dmem_ram_1729), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n767) );
NAND2_X1 MEM_stage_inst_dmem_U930 ( .A1(MEM_stage_inst_dmem_ram_1601), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n768) );
NOR2_X1 MEM_stage_inst_dmem_U929 ( .A1(MEM_stage_inst_dmem_n766), .A2(MEM_stage_inst_dmem_n765), .ZN(MEM_stage_inst_dmem_n774) );
NAND2_X1 MEM_stage_inst_dmem_U928 ( .A1(MEM_stage_inst_dmem_n764), .A2(MEM_stage_inst_dmem_n763), .ZN(MEM_stage_inst_dmem_n765) );
NAND2_X1 MEM_stage_inst_dmem_U927 ( .A1(MEM_stage_inst_dmem_ram_1665), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n763) );
NAND2_X1 MEM_stage_inst_dmem_U926 ( .A1(MEM_stage_inst_dmem_ram_1745), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n764) );
NAND2_X1 MEM_stage_inst_dmem_U925 ( .A1(MEM_stage_inst_dmem_n762), .A2(MEM_stage_inst_dmem_n761), .ZN(MEM_stage_inst_dmem_n766) );
NAND2_X1 MEM_stage_inst_dmem_U924 ( .A1(MEM_stage_inst_dmem_ram_1441), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n761) );
NAND2_X1 MEM_stage_inst_dmem_U923 ( .A1(MEM_stage_inst_dmem_ram_1137), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n762) );
NAND2_X1 MEM_stage_inst_dmem_U922 ( .A1(MEM_stage_inst_dmem_n760), .A2(MEM_stage_inst_dmem_n759), .ZN(MEM_stage_inst_mem_read_data_0) );
NOR2_X1 MEM_stage_inst_dmem_U921 ( .A1(MEM_stage_inst_dmem_n758), .A2(MEM_stage_inst_dmem_n757), .ZN(MEM_stage_inst_dmem_n759) );
NOR2_X1 MEM_stage_inst_dmem_U920 ( .A1(MEM_stage_inst_dmem_n756), .A2(MEM_stage_inst_dmem_n8417), .ZN(MEM_stage_inst_dmem_n757) );
OR2_X1 MEM_stage_inst_dmem_U919 ( .A1(EX_pipeline_reg_out_28), .A2(EX_pipeline_reg_out_29), .ZN(MEM_stage_inst_dmem_n8417) );
NOR2_X1 MEM_stage_inst_dmem_U918 ( .A1(MEM_stage_inst_dmem_n755), .A2(MEM_stage_inst_dmem_n754), .ZN(MEM_stage_inst_dmem_n756) );
NAND2_X1 MEM_stage_inst_dmem_U917 ( .A1(MEM_stage_inst_dmem_n753), .A2(MEM_stage_inst_dmem_n752), .ZN(MEM_stage_inst_dmem_n754) );
NOR2_X1 MEM_stage_inst_dmem_U916 ( .A1(MEM_stage_inst_dmem_n751), .A2(MEM_stage_inst_dmem_n750), .ZN(MEM_stage_inst_dmem_n752) );
NAND2_X1 MEM_stage_inst_dmem_U915 ( .A1(MEM_stage_inst_dmem_n749), .A2(MEM_stage_inst_dmem_n748), .ZN(MEM_stage_inst_dmem_n750) );
NOR2_X1 MEM_stage_inst_dmem_U914 ( .A1(MEM_stage_inst_dmem_n747), .A2(MEM_stage_inst_dmem_n746), .ZN(MEM_stage_inst_dmem_n748) );
NAND2_X1 MEM_stage_inst_dmem_U913 ( .A1(MEM_stage_inst_dmem_n745), .A2(MEM_stage_inst_dmem_n744), .ZN(MEM_stage_inst_dmem_n746) );
NAND2_X1 MEM_stage_inst_dmem_U912 ( .A1(MEM_stage_inst_dmem_ram_3088), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n744) );
NAND2_X1 MEM_stage_inst_dmem_U911 ( .A1(MEM_stage_inst_dmem_ram_3520), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n745) );
NAND2_X1 MEM_stage_inst_dmem_U910 ( .A1(MEM_stage_inst_dmem_n743), .A2(MEM_stage_inst_dmem_n742), .ZN(MEM_stage_inst_dmem_n747) );
NAND2_X1 MEM_stage_inst_dmem_U909 ( .A1(MEM_stage_inst_dmem_ram_3920), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n742) );
NAND2_X1 MEM_stage_inst_dmem_U908 ( .A1(MEM_stage_inst_dmem_ram_3712), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n743) );
NOR2_X1 MEM_stage_inst_dmem_U907 ( .A1(MEM_stage_inst_dmem_n741), .A2(MEM_stage_inst_dmem_n740), .ZN(MEM_stage_inst_dmem_n749) );
NAND2_X1 MEM_stage_inst_dmem_U906 ( .A1(MEM_stage_inst_dmem_n739), .A2(MEM_stage_inst_dmem_n738), .ZN(MEM_stage_inst_dmem_n740) );
NAND2_X1 MEM_stage_inst_dmem_U905 ( .A1(MEM_stage_inst_dmem_ram_3760), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n738) );
NAND2_X1 MEM_stage_inst_dmem_U904 ( .A1(MEM_stage_inst_dmem_ram_3280), .A2(MEM_stage_inst_dmem_n51), .ZN(MEM_stage_inst_dmem_n739) );
NAND2_X1 MEM_stage_inst_dmem_U903 ( .A1(MEM_stage_inst_dmem_n737), .A2(MEM_stage_inst_dmem_n736), .ZN(MEM_stage_inst_dmem_n741) );
NAND2_X1 MEM_stage_inst_dmem_U902 ( .A1(MEM_stage_inst_dmem_ram_3184), .A2(MEM_stage_inst_dmem_n4710), .ZN(MEM_stage_inst_dmem_n736) );
NAND2_X1 MEM_stage_inst_dmem_U901 ( .A1(MEM_stage_inst_dmem_ram_3664), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n737) );
NAND2_X1 MEM_stage_inst_dmem_U900 ( .A1(MEM_stage_inst_dmem_n735), .A2(MEM_stage_inst_dmem_n734), .ZN(MEM_stage_inst_dmem_n751) );
NOR2_X1 MEM_stage_inst_dmem_U899 ( .A1(MEM_stage_inst_dmem_n733), .A2(MEM_stage_inst_dmem_n732), .ZN(MEM_stage_inst_dmem_n734) );
NAND2_X1 MEM_stage_inst_dmem_U898 ( .A1(MEM_stage_inst_dmem_n731), .A2(MEM_stage_inst_dmem_n730), .ZN(MEM_stage_inst_dmem_n732) );
NAND2_X1 MEM_stage_inst_dmem_U897 ( .A1(MEM_stage_inst_dmem_ram_3376), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n730) );
NAND2_X1 MEM_stage_inst_dmem_U896 ( .A1(MEM_stage_inst_dmem_ram_3408), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n731) );
NAND2_X1 MEM_stage_inst_dmem_U895 ( .A1(MEM_stage_inst_dmem_n729), .A2(MEM_stage_inst_dmem_n728), .ZN(MEM_stage_inst_dmem_n733) );
NAND2_X1 MEM_stage_inst_dmem_U894 ( .A1(MEM_stage_inst_dmem_ram_3248), .A2(MEM_stage_inst_dmem_n55), .ZN(MEM_stage_inst_dmem_n728) );
NAND2_X1 MEM_stage_inst_dmem_U893 ( .A1(MEM_stage_inst_dmem_ram_3168), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n729) );
NOR2_X1 MEM_stage_inst_dmem_U892 ( .A1(MEM_stage_inst_dmem_n727), .A2(MEM_stage_inst_dmem_n726), .ZN(MEM_stage_inst_dmem_n735) );
NAND2_X1 MEM_stage_inst_dmem_U891 ( .A1(MEM_stage_inst_dmem_n725), .A2(MEM_stage_inst_dmem_n724), .ZN(MEM_stage_inst_dmem_n726) );
NAND2_X1 MEM_stage_inst_dmem_U890 ( .A1(MEM_stage_inst_dmem_ram_3904), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n724) );
NAND2_X1 MEM_stage_inst_dmem_U889 ( .A1(MEM_stage_inst_dmem_ram_3744), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n725) );
NAND2_X1 MEM_stage_inst_dmem_U888 ( .A1(MEM_stage_inst_dmem_n723), .A2(MEM_stage_inst_dmem_n722), .ZN(MEM_stage_inst_dmem_n727) );
NAND2_X1 MEM_stage_inst_dmem_U887 ( .A1(MEM_stage_inst_dmem_ram_3776), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n722) );
NAND2_X1 MEM_stage_inst_dmem_U886 ( .A1(MEM_stage_inst_dmem_ram_4080), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n723) );
NOR2_X1 MEM_stage_inst_dmem_U885 ( .A1(MEM_stage_inst_dmem_n721), .A2(MEM_stage_inst_dmem_n720), .ZN(MEM_stage_inst_dmem_n753) );
NAND2_X1 MEM_stage_inst_dmem_U884 ( .A1(MEM_stage_inst_dmem_n719), .A2(MEM_stage_inst_dmem_n718), .ZN(MEM_stage_inst_dmem_n720) );
NOR2_X1 MEM_stage_inst_dmem_U883 ( .A1(MEM_stage_inst_dmem_n717), .A2(MEM_stage_inst_dmem_n716), .ZN(MEM_stage_inst_dmem_n718) );
NAND2_X1 MEM_stage_inst_dmem_U882 ( .A1(MEM_stage_inst_dmem_n715), .A2(MEM_stage_inst_dmem_n714), .ZN(MEM_stage_inst_dmem_n716) );
NAND2_X1 MEM_stage_inst_dmem_U881 ( .A1(MEM_stage_inst_dmem_ram_3200), .A2(MEM_stage_inst_dmem_n61), .ZN(MEM_stage_inst_dmem_n714) );
NAND2_X1 MEM_stage_inst_dmem_U880 ( .A1(MEM_stage_inst_dmem_ram_3344), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n715) );
NAND2_X1 MEM_stage_inst_dmem_U879 ( .A1(MEM_stage_inst_dmem_n713), .A2(MEM_stage_inst_dmem_n712), .ZN(MEM_stage_inst_dmem_n717) );
NAND2_X1 MEM_stage_inst_dmem_U878 ( .A1(MEM_stage_inst_dmem_ram_3936), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n712) );
NAND2_X1 MEM_stage_inst_dmem_U877 ( .A1(MEM_stage_inst_dmem_ram_4000), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n713) );
NOR2_X1 MEM_stage_inst_dmem_U876 ( .A1(MEM_stage_inst_dmem_n711), .A2(MEM_stage_inst_dmem_n710), .ZN(MEM_stage_inst_dmem_n719) );
NAND2_X1 MEM_stage_inst_dmem_U875 ( .A1(MEM_stage_inst_dmem_n709), .A2(MEM_stage_inst_dmem_n708), .ZN(MEM_stage_inst_dmem_n710) );
NAND2_X1 MEM_stage_inst_dmem_U874 ( .A1(MEM_stage_inst_dmem_ram_3568), .A2(MEM_stage_inst_dmem_n8535), .ZN(MEM_stage_inst_dmem_n708) );
NAND2_X1 MEM_stage_inst_dmem_U873 ( .A1(MEM_stage_inst_dmem_ram_3536), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n709) );
NAND2_X1 MEM_stage_inst_dmem_U872 ( .A1(MEM_stage_inst_dmem_n707), .A2(MEM_stage_inst_dmem_n706), .ZN(MEM_stage_inst_dmem_n711) );
NAND2_X1 MEM_stage_inst_dmem_U871 ( .A1(MEM_stage_inst_dmem_ram_3392), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n706) );
NAND2_X1 MEM_stage_inst_dmem_U870 ( .A1(MEM_stage_inst_dmem_ram_3360), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n707) );
NAND2_X1 MEM_stage_inst_dmem_U869 ( .A1(MEM_stage_inst_dmem_n705), .A2(MEM_stage_inst_dmem_n704), .ZN(MEM_stage_inst_dmem_n721) );
NOR2_X1 MEM_stage_inst_dmem_U868 ( .A1(MEM_stage_inst_dmem_n703), .A2(MEM_stage_inst_dmem_n702), .ZN(MEM_stage_inst_dmem_n704) );
NAND2_X1 MEM_stage_inst_dmem_U867 ( .A1(MEM_stage_inst_dmem_n701), .A2(MEM_stage_inst_dmem_n700), .ZN(MEM_stage_inst_dmem_n702) );
NAND2_X1 MEM_stage_inst_dmem_U866 ( .A1(MEM_stage_inst_dmem_ram_3120), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n700) );
NAND2_X1 MEM_stage_inst_dmem_U865 ( .A1(MEM_stage_inst_dmem_ram_3968), .A2(MEM_stage_inst_dmem_n72), .ZN(MEM_stage_inst_dmem_n701) );
NAND2_X1 MEM_stage_inst_dmem_U864 ( .A1(MEM_stage_inst_dmem_n699), .A2(MEM_stage_inst_dmem_n698), .ZN(MEM_stage_inst_dmem_n703) );
NAND2_X1 MEM_stage_inst_dmem_U863 ( .A1(MEM_stage_inst_dmem_ram_3232), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n698) );
NAND2_X1 MEM_stage_inst_dmem_U862 ( .A1(MEM_stage_inst_dmem_ram_3584), .A2(MEM_stage_inst_dmem_n71), .ZN(MEM_stage_inst_dmem_n699) );
NOR2_X1 MEM_stage_inst_dmem_U861 ( .A1(MEM_stage_inst_dmem_n697), .A2(MEM_stage_inst_dmem_n696), .ZN(MEM_stage_inst_dmem_n705) );
NAND2_X1 MEM_stage_inst_dmem_U860 ( .A1(MEM_stage_inst_dmem_n695), .A2(MEM_stage_inst_dmem_n694), .ZN(MEM_stage_inst_dmem_n696) );
NAND2_X1 MEM_stage_inst_dmem_U859 ( .A1(MEM_stage_inst_dmem_ram_3296), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n694) );
NAND2_X1 MEM_stage_inst_dmem_U858 ( .A1(MEM_stage_inst_dmem_ram_3136), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n695) );
NAND2_X1 MEM_stage_inst_dmem_U857 ( .A1(MEM_stage_inst_dmem_n693), .A2(MEM_stage_inst_dmem_n692), .ZN(MEM_stage_inst_dmem_n697) );
NAND2_X1 MEM_stage_inst_dmem_U856 ( .A1(MEM_stage_inst_dmem_ram_3680), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n692) );
NAND2_X1 MEM_stage_inst_dmem_U855 ( .A1(MEM_stage_inst_dmem_ram_3792), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n693) );
NAND2_X1 MEM_stage_inst_dmem_U854 ( .A1(MEM_stage_inst_dmem_n691), .A2(MEM_stage_inst_dmem_n690), .ZN(MEM_stage_inst_dmem_n755) );
NOR2_X1 MEM_stage_inst_dmem_U853 ( .A1(MEM_stage_inst_dmem_n689), .A2(MEM_stage_inst_dmem_n688), .ZN(MEM_stage_inst_dmem_n690) );
NAND2_X1 MEM_stage_inst_dmem_U852 ( .A1(MEM_stage_inst_dmem_n687), .A2(MEM_stage_inst_dmem_n686), .ZN(MEM_stage_inst_dmem_n688) );
NOR2_X1 MEM_stage_inst_dmem_U851 ( .A1(MEM_stage_inst_dmem_n685), .A2(MEM_stage_inst_dmem_n684), .ZN(MEM_stage_inst_dmem_n686) );
NAND2_X1 MEM_stage_inst_dmem_U850 ( .A1(MEM_stage_inst_dmem_n683), .A2(MEM_stage_inst_dmem_n682), .ZN(MEM_stage_inst_dmem_n684) );
NAND2_X1 MEM_stage_inst_dmem_U849 ( .A1(MEM_stage_inst_dmem_ram_3696), .A2(MEM_stage_inst_dmem_n4652), .ZN(MEM_stage_inst_dmem_n682) );
NAND2_X1 MEM_stage_inst_dmem_U848 ( .A1(MEM_stage_inst_dmem_ram_3440), .A2(MEM_stage_inst_dmem_n4721), .ZN(MEM_stage_inst_dmem_n683) );
NAND2_X1 MEM_stage_inst_dmem_U847 ( .A1(MEM_stage_inst_dmem_n681), .A2(MEM_stage_inst_dmem_n680), .ZN(MEM_stage_inst_dmem_n685) );
NAND2_X1 MEM_stage_inst_dmem_U846 ( .A1(MEM_stage_inst_dmem_ram_4016), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n680) );
NAND2_X1 MEM_stage_inst_dmem_U845 ( .A1(MEM_stage_inst_dmem_ram_4048), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n681) );
NOR2_X1 MEM_stage_inst_dmem_U844 ( .A1(MEM_stage_inst_dmem_n679), .A2(MEM_stage_inst_dmem_n678), .ZN(MEM_stage_inst_dmem_n687) );
NAND2_X1 MEM_stage_inst_dmem_U843 ( .A1(MEM_stage_inst_dmem_n677), .A2(MEM_stage_inst_dmem_n676), .ZN(MEM_stage_inst_dmem_n678) );
NAND2_X1 MEM_stage_inst_dmem_U842 ( .A1(MEM_stage_inst_dmem_ram_3264), .A2(MEM_stage_inst_dmem_n36), .ZN(MEM_stage_inst_dmem_n676) );
NAND2_X1 MEM_stage_inst_dmem_U841 ( .A1(MEM_stage_inst_dmem_ram_3840), .A2(MEM_stage_inst_dmem_n37), .ZN(MEM_stage_inst_dmem_n677) );
NAND2_X1 MEM_stage_inst_dmem_U840 ( .A1(MEM_stage_inst_dmem_n675), .A2(MEM_stage_inst_dmem_n674), .ZN(MEM_stage_inst_dmem_n679) );
NAND2_X1 MEM_stage_inst_dmem_U839 ( .A1(MEM_stage_inst_dmem_ram_3856), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n674) );
NAND2_X1 MEM_stage_inst_dmem_U838 ( .A1(MEM_stage_inst_dmem_ram_3328), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n675) );
NAND2_X1 MEM_stage_inst_dmem_U837 ( .A1(MEM_stage_inst_dmem_n673), .A2(MEM_stage_inst_dmem_n672), .ZN(MEM_stage_inst_dmem_n689) );
NOR2_X1 MEM_stage_inst_dmem_U836 ( .A1(MEM_stage_inst_dmem_n671), .A2(MEM_stage_inst_dmem_n670), .ZN(MEM_stage_inst_dmem_n672) );
NAND2_X1 MEM_stage_inst_dmem_U835 ( .A1(MEM_stage_inst_dmem_n669), .A2(MEM_stage_inst_dmem_n668), .ZN(MEM_stage_inst_dmem_n670) );
NAND2_X1 MEM_stage_inst_dmem_U834 ( .A1(MEM_stage_inst_dmem_ram_3312), .A2(MEM_stage_inst_dmem_n39), .ZN(MEM_stage_inst_dmem_n668) );
NAND2_X1 MEM_stage_inst_dmem_U833 ( .A1(MEM_stage_inst_dmem_ram_3152), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n669) );
NAND2_X1 MEM_stage_inst_dmem_U832 ( .A1(MEM_stage_inst_dmem_n667), .A2(MEM_stage_inst_dmem_n666), .ZN(MEM_stage_inst_dmem_n671) );
NAND2_X1 MEM_stage_inst_dmem_U831 ( .A1(MEM_stage_inst_dmem_ram_3632), .A2(MEM_stage_inst_dmem_n41), .ZN(MEM_stage_inst_dmem_n666) );
NAND2_X1 MEM_stage_inst_dmem_U830 ( .A1(MEM_stage_inst_dmem_ram_4032), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n667) );
NOR2_X1 MEM_stage_inst_dmem_U829 ( .A1(MEM_stage_inst_dmem_n665), .A2(MEM_stage_inst_dmem_n664), .ZN(MEM_stage_inst_dmem_n673) );
NAND2_X1 MEM_stage_inst_dmem_U828 ( .A1(MEM_stage_inst_dmem_n663), .A2(MEM_stage_inst_dmem_n662), .ZN(MEM_stage_inst_dmem_n664) );
NAND2_X1 MEM_stage_inst_dmem_U827 ( .A1(MEM_stage_inst_dmem_ram_3504), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n662) );
NAND2_X1 MEM_stage_inst_dmem_U826 ( .A1(MEM_stage_inst_dmem_ram_3216), .A2(MEM_stage_inst_dmem_n5807), .ZN(MEM_stage_inst_dmem_n663) );
NAND2_X1 MEM_stage_inst_dmem_U825 ( .A1(MEM_stage_inst_dmem_n661), .A2(MEM_stage_inst_dmem_n660), .ZN(MEM_stage_inst_dmem_n665) );
NAND2_X1 MEM_stage_inst_dmem_U824 ( .A1(MEM_stage_inst_dmem_ram_3104), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n660) );
NAND2_X1 MEM_stage_inst_dmem_U823 ( .A1(MEM_stage_inst_dmem_ram_3600), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n661) );
NOR2_X1 MEM_stage_inst_dmem_U822 ( .A1(MEM_stage_inst_dmem_n659), .A2(MEM_stage_inst_dmem_n658), .ZN(MEM_stage_inst_dmem_n691) );
NAND2_X1 MEM_stage_inst_dmem_U821 ( .A1(MEM_stage_inst_dmem_n657), .A2(MEM_stage_inst_dmem_n656), .ZN(MEM_stage_inst_dmem_n658) );
NOR2_X1 MEM_stage_inst_dmem_U820 ( .A1(MEM_stage_inst_dmem_n655), .A2(MEM_stage_inst_dmem_n654), .ZN(MEM_stage_inst_dmem_n656) );
NAND2_X1 MEM_stage_inst_dmem_U819 ( .A1(MEM_stage_inst_dmem_n653), .A2(MEM_stage_inst_dmem_n652), .ZN(MEM_stage_inst_dmem_n654) );
NAND2_X1 MEM_stage_inst_dmem_U818 ( .A1(MEM_stage_inst_dmem_ram_3616), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n652) );
NAND2_X1 MEM_stage_inst_dmem_U817 ( .A1(MEM_stage_inst_dmem_ram_3456), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n653) );
NAND2_X1 MEM_stage_inst_dmem_U816 ( .A1(MEM_stage_inst_dmem_n651), .A2(MEM_stage_inst_dmem_n650), .ZN(MEM_stage_inst_dmem_n655) );
NAND2_X1 MEM_stage_inst_dmem_U815 ( .A1(MEM_stage_inst_dmem_ram_3888), .A2(MEM_stage_inst_dmem_n46), .ZN(MEM_stage_inst_dmem_n650) );
NAND2_X1 MEM_stage_inst_dmem_U814 ( .A1(MEM_stage_inst_dmem_ram_3728), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n651) );
NOR2_X1 MEM_stage_inst_dmem_U813 ( .A1(MEM_stage_inst_dmem_n649), .A2(MEM_stage_inst_dmem_n648), .ZN(MEM_stage_inst_dmem_n657) );
NAND2_X1 MEM_stage_inst_dmem_U812 ( .A1(MEM_stage_inst_dmem_n647), .A2(MEM_stage_inst_dmem_n646), .ZN(MEM_stage_inst_dmem_n648) );
NAND2_X1 MEM_stage_inst_dmem_U811 ( .A1(MEM_stage_inst_dmem_ram_4064), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n646) );
NAND2_X1 MEM_stage_inst_dmem_U810 ( .A1(MEM_stage_inst_dmem_ram_3488), .A2(MEM_stage_inst_dmem_n4772), .ZN(MEM_stage_inst_dmem_n647) );
NAND2_X1 MEM_stage_inst_dmem_U809 ( .A1(MEM_stage_inst_dmem_n645), .A2(MEM_stage_inst_dmem_n644), .ZN(MEM_stage_inst_dmem_n649) );
NAND2_X1 MEM_stage_inst_dmem_U808 ( .A1(MEM_stage_inst_dmem_ram_3552), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n644) );
NAND2_X1 MEM_stage_inst_dmem_U807 ( .A1(MEM_stage_inst_dmem_ram_3824), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n645) );
NAND2_X1 MEM_stage_inst_dmem_U806 ( .A1(MEM_stage_inst_dmem_n643), .A2(MEM_stage_inst_dmem_n642), .ZN(MEM_stage_inst_dmem_n659) );
NOR2_X1 MEM_stage_inst_dmem_U805 ( .A1(MEM_stage_inst_dmem_n641), .A2(MEM_stage_inst_dmem_n640), .ZN(MEM_stage_inst_dmem_n642) );
NAND2_X1 MEM_stage_inst_dmem_U804 ( .A1(MEM_stage_inst_dmem_n639), .A2(MEM_stage_inst_dmem_n638), .ZN(MEM_stage_inst_dmem_n640) );
NAND2_X1 MEM_stage_inst_dmem_U803 ( .A1(MEM_stage_inst_dmem_ram_3952), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n638) );
NAND2_X1 MEM_stage_inst_dmem_U802 ( .A1(MEM_stage_inst_dmem_ram_3808), .A2(MEM_stage_inst_dmem_n4769), .ZN(MEM_stage_inst_dmem_n639) );
NAND2_X1 MEM_stage_inst_dmem_U801 ( .A1(MEM_stage_inst_dmem_n637), .A2(MEM_stage_inst_dmem_n636), .ZN(MEM_stage_inst_dmem_n641) );
NAND2_X1 MEM_stage_inst_dmem_U800 ( .A1(MEM_stage_inst_dmem_ram_3472), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n636) );
NAND2_X1 MEM_stage_inst_dmem_U799 ( .A1(MEM_stage_inst_dmem_ram_3984), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n637) );
NOR2_X1 MEM_stage_inst_dmem_U798 ( .A1(MEM_stage_inst_dmem_n635), .A2(MEM_stage_inst_dmem_n634), .ZN(MEM_stage_inst_dmem_n643) );
NAND2_X1 MEM_stage_inst_dmem_U797 ( .A1(MEM_stage_inst_dmem_n633), .A2(MEM_stage_inst_dmem_n632), .ZN(MEM_stage_inst_dmem_n634) );
NAND2_X1 MEM_stage_inst_dmem_U796 ( .A1(MEM_stage_inst_dmem_ram_3424), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n632) );
NAND2_X1 MEM_stage_inst_dmem_U795 ( .A1(MEM_stage_inst_dmem_ram_3072), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n633) );
NAND2_X1 MEM_stage_inst_dmem_U794 ( .A1(MEM_stage_inst_dmem_n631), .A2(MEM_stage_inst_dmem_n630), .ZN(MEM_stage_inst_dmem_n635) );
NAND2_X1 MEM_stage_inst_dmem_U793 ( .A1(MEM_stage_inst_dmem_ram_3872), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n630) );
NAND2_X1 MEM_stage_inst_dmem_U792 ( .A1(MEM_stage_inst_dmem_ram_3648), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n631) );
NOR2_X1 MEM_stage_inst_dmem_U791 ( .A1(MEM_stage_inst_dmem_n629), .A2(MEM_stage_inst_dmem_n8152), .ZN(MEM_stage_inst_dmem_n758) );
NAND2_X1 MEM_stage_inst_dmem_U790 ( .A1(EX_pipeline_reg_out_29), .A2(MEM_stage_inst_dmem_n15967), .ZN(MEM_stage_inst_dmem_n8152) );
NOR2_X1 MEM_stage_inst_dmem_U789 ( .A1(MEM_stage_inst_dmem_n628), .A2(MEM_stage_inst_dmem_n627), .ZN(MEM_stage_inst_dmem_n629) );
NAND2_X1 MEM_stage_inst_dmem_U788 ( .A1(MEM_stage_inst_dmem_n626), .A2(MEM_stage_inst_dmem_n625), .ZN(MEM_stage_inst_dmem_n627) );
NOR2_X1 MEM_stage_inst_dmem_U787 ( .A1(MEM_stage_inst_dmem_n624), .A2(MEM_stage_inst_dmem_n623), .ZN(MEM_stage_inst_dmem_n625) );
NAND2_X1 MEM_stage_inst_dmem_U786 ( .A1(MEM_stage_inst_dmem_n622), .A2(MEM_stage_inst_dmem_n621), .ZN(MEM_stage_inst_dmem_n623) );
NOR2_X1 MEM_stage_inst_dmem_U785 ( .A1(MEM_stage_inst_dmem_n620), .A2(MEM_stage_inst_dmem_n619), .ZN(MEM_stage_inst_dmem_n621) );
NAND2_X1 MEM_stage_inst_dmem_U784 ( .A1(MEM_stage_inst_dmem_n618), .A2(MEM_stage_inst_dmem_n617), .ZN(MEM_stage_inst_dmem_n619) );
NAND2_X1 MEM_stage_inst_dmem_U783 ( .A1(MEM_stage_inst_dmem_ram_1968), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n617) );
NAND2_X1 MEM_stage_inst_dmem_U782 ( .A1(MEM_stage_inst_dmem_ram_1280), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n618) );
NAND2_X1 MEM_stage_inst_dmem_U781 ( .A1(MEM_stage_inst_dmem_n616), .A2(MEM_stage_inst_dmem_n615), .ZN(MEM_stage_inst_dmem_n620) );
NAND2_X1 MEM_stage_inst_dmem_U780 ( .A1(MEM_stage_inst_dmem_ram_1904), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n615) );
NAND2_X1 MEM_stage_inst_dmem_U779 ( .A1(MEM_stage_inst_dmem_ram_1040), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n616) );
NOR2_X1 MEM_stage_inst_dmem_U778 ( .A1(MEM_stage_inst_dmem_n614), .A2(MEM_stage_inst_dmem_n613), .ZN(MEM_stage_inst_dmem_n622) );
NAND2_X1 MEM_stage_inst_dmem_U777 ( .A1(MEM_stage_inst_dmem_n612), .A2(MEM_stage_inst_dmem_n611), .ZN(MEM_stage_inst_dmem_n613) );
NAND2_X1 MEM_stage_inst_dmem_U776 ( .A1(MEM_stage_inst_dmem_ram_1424), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n611) );
NAND2_X1 MEM_stage_inst_dmem_U775 ( .A1(MEM_stage_inst_dmem_ram_1712), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n612) );
NAND2_X1 MEM_stage_inst_dmem_U774 ( .A1(MEM_stage_inst_dmem_n610), .A2(MEM_stage_inst_dmem_n609), .ZN(MEM_stage_inst_dmem_n614) );
NAND2_X1 MEM_stage_inst_dmem_U773 ( .A1(MEM_stage_inst_dmem_ram_1152), .A2(MEM_stage_inst_dmem_n61), .ZN(MEM_stage_inst_dmem_n609) );
NAND2_X1 MEM_stage_inst_dmem_U772 ( .A1(MEM_stage_inst_dmem_ram_1488), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n610) );
NAND2_X1 MEM_stage_inst_dmem_U771 ( .A1(MEM_stage_inst_dmem_n608), .A2(MEM_stage_inst_dmem_n607), .ZN(MEM_stage_inst_dmem_n624) );
NOR2_X1 MEM_stage_inst_dmem_U770 ( .A1(MEM_stage_inst_dmem_n606), .A2(MEM_stage_inst_dmem_n605), .ZN(MEM_stage_inst_dmem_n607) );
NAND2_X1 MEM_stage_inst_dmem_U769 ( .A1(MEM_stage_inst_dmem_n604), .A2(MEM_stage_inst_dmem_n603), .ZN(MEM_stage_inst_dmem_n605) );
NAND2_X1 MEM_stage_inst_dmem_U768 ( .A1(MEM_stage_inst_dmem_ram_1728), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n603) );
NAND2_X1 MEM_stage_inst_dmem_U767 ( .A1(MEM_stage_inst_dmem_ram_1760), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n604) );
NAND2_X1 MEM_stage_inst_dmem_U766 ( .A1(MEM_stage_inst_dmem_n602), .A2(MEM_stage_inst_dmem_n601), .ZN(MEM_stage_inst_dmem_n606) );
NAND2_X1 MEM_stage_inst_dmem_U765 ( .A1(MEM_stage_inst_dmem_ram_1584), .A2(MEM_stage_inst_dmem_n41), .ZN(MEM_stage_inst_dmem_n601) );
NAND2_X1 MEM_stage_inst_dmem_U764 ( .A1(MEM_stage_inst_dmem_ram_1776), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n602) );
NOR2_X1 MEM_stage_inst_dmem_U763 ( .A1(MEM_stage_inst_dmem_n600), .A2(MEM_stage_inst_dmem_n599), .ZN(MEM_stage_inst_dmem_n608) );
NAND2_X1 MEM_stage_inst_dmem_U762 ( .A1(MEM_stage_inst_dmem_n598), .A2(MEM_stage_inst_dmem_n597), .ZN(MEM_stage_inst_dmem_n599) );
NAND2_X1 MEM_stage_inst_dmem_U761 ( .A1(MEM_stage_inst_dmem_ram_1216), .A2(MEM_stage_inst_dmem_n36), .ZN(MEM_stage_inst_dmem_n597) );
NAND2_X1 MEM_stage_inst_dmem_U760 ( .A1(MEM_stage_inst_dmem_ram_1536), .A2(MEM_stage_inst_dmem_n71), .ZN(MEM_stage_inst_dmem_n598) );
NAND2_X1 MEM_stage_inst_dmem_U759 ( .A1(MEM_stage_inst_dmem_n596), .A2(MEM_stage_inst_dmem_n595), .ZN(MEM_stage_inst_dmem_n600) );
NAND2_X1 MEM_stage_inst_dmem_U758 ( .A1(MEM_stage_inst_dmem_ram_1792), .A2(MEM_stage_inst_dmem_n37), .ZN(MEM_stage_inst_dmem_n595) );
NAND2_X1 MEM_stage_inst_dmem_U757 ( .A1(MEM_stage_inst_dmem_ram_1600), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n596) );
NOR2_X1 MEM_stage_inst_dmem_U756 ( .A1(MEM_stage_inst_dmem_n594), .A2(MEM_stage_inst_dmem_n593), .ZN(MEM_stage_inst_dmem_n626) );
NAND2_X1 MEM_stage_inst_dmem_U755 ( .A1(MEM_stage_inst_dmem_n592), .A2(MEM_stage_inst_dmem_n591), .ZN(MEM_stage_inst_dmem_n593) );
NOR2_X1 MEM_stage_inst_dmem_U754 ( .A1(MEM_stage_inst_dmem_n590), .A2(MEM_stage_inst_dmem_n589), .ZN(MEM_stage_inst_dmem_n591) );
NAND2_X1 MEM_stage_inst_dmem_U753 ( .A1(MEM_stage_inst_dmem_n588), .A2(MEM_stage_inst_dmem_n587), .ZN(MEM_stage_inst_dmem_n589) );
NAND2_X1 MEM_stage_inst_dmem_U752 ( .A1(MEM_stage_inst_dmem_ram_1168), .A2(MEM_stage_inst_dmem_n44), .ZN(MEM_stage_inst_dmem_n587) );
NAND2_X1 MEM_stage_inst_dmem_U751 ( .A1(MEM_stage_inst_dmem_ram_1024), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n588) );
NAND2_X1 MEM_stage_inst_dmem_U750 ( .A1(MEM_stage_inst_dmem_n586), .A2(MEM_stage_inst_dmem_n585), .ZN(MEM_stage_inst_dmem_n590) );
NAND2_X1 MEM_stage_inst_dmem_U749 ( .A1(MEM_stage_inst_dmem_ram_1696), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n585) );
NAND2_X1 MEM_stage_inst_dmem_U748 ( .A1(MEM_stage_inst_dmem_ram_1184), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n586) );
NOR2_X1 MEM_stage_inst_dmem_U747 ( .A1(MEM_stage_inst_dmem_n584), .A2(MEM_stage_inst_dmem_n583), .ZN(MEM_stage_inst_dmem_n592) );
NAND2_X1 MEM_stage_inst_dmem_U746 ( .A1(MEM_stage_inst_dmem_n582), .A2(MEM_stage_inst_dmem_n581), .ZN(MEM_stage_inst_dmem_n583) );
NAND2_X1 MEM_stage_inst_dmem_U745 ( .A1(MEM_stage_inst_dmem_ram_1264), .A2(MEM_stage_inst_dmem_n39), .ZN(MEM_stage_inst_dmem_n581) );
NAND2_X1 MEM_stage_inst_dmem_U744 ( .A1(MEM_stage_inst_dmem_ram_2032), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n582) );
NAND2_X1 MEM_stage_inst_dmem_U743 ( .A1(MEM_stage_inst_dmem_n580), .A2(MEM_stage_inst_dmem_n579), .ZN(MEM_stage_inst_dmem_n584) );
NAND2_X1 MEM_stage_inst_dmem_U742 ( .A1(MEM_stage_inst_dmem_ram_1520), .A2(MEM_stage_inst_dmem_n8535), .ZN(MEM_stage_inst_dmem_n579) );
NAND2_X1 MEM_stage_inst_dmem_U741 ( .A1(MEM_stage_inst_dmem_ram_1312), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n580) );
NAND2_X1 MEM_stage_inst_dmem_U740 ( .A1(MEM_stage_inst_dmem_n578), .A2(MEM_stage_inst_dmem_n577), .ZN(MEM_stage_inst_dmem_n594) );
NOR2_X1 MEM_stage_inst_dmem_U739 ( .A1(MEM_stage_inst_dmem_n576), .A2(MEM_stage_inst_dmem_n575), .ZN(MEM_stage_inst_dmem_n577) );
NAND2_X1 MEM_stage_inst_dmem_U738 ( .A1(MEM_stage_inst_dmem_n574), .A2(MEM_stage_inst_dmem_n573), .ZN(MEM_stage_inst_dmem_n575) );
NAND2_X1 MEM_stage_inst_dmem_U737 ( .A1(MEM_stage_inst_dmem_ram_1664), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n573) );
NAND2_X1 MEM_stage_inst_dmem_U736 ( .A1(MEM_stage_inst_dmem_ram_1056), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n574) );
NAND2_X1 MEM_stage_inst_dmem_U735 ( .A1(MEM_stage_inst_dmem_n572), .A2(MEM_stage_inst_dmem_n571), .ZN(MEM_stage_inst_dmem_n576) );
NAND2_X1 MEM_stage_inst_dmem_U734 ( .A1(MEM_stage_inst_dmem_ram_1632), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n571) );
NAND2_X1 MEM_stage_inst_dmem_U733 ( .A1(MEM_stage_inst_dmem_ram_1680), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n572) );
NOR2_X1 MEM_stage_inst_dmem_U732 ( .A1(MEM_stage_inst_dmem_n570), .A2(MEM_stage_inst_dmem_n569), .ZN(MEM_stage_inst_dmem_n578) );
NAND2_X1 MEM_stage_inst_dmem_U731 ( .A1(MEM_stage_inst_dmem_n568), .A2(MEM_stage_inst_dmem_n567), .ZN(MEM_stage_inst_dmem_n569) );
NAND2_X1 MEM_stage_inst_dmem_U730 ( .A1(MEM_stage_inst_dmem_ram_1328), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n567) );
NAND2_X1 MEM_stage_inst_dmem_U729 ( .A1(MEM_stage_inst_dmem_ram_1552), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n568) );
NAND2_X1 MEM_stage_inst_dmem_U728 ( .A1(MEM_stage_inst_dmem_n566), .A2(MEM_stage_inst_dmem_n565), .ZN(MEM_stage_inst_dmem_n570) );
NAND2_X1 MEM_stage_inst_dmem_U727 ( .A1(MEM_stage_inst_dmem_ram_2000), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n565) );
NAND2_X1 MEM_stage_inst_dmem_U726 ( .A1(MEM_stage_inst_dmem_ram_1808), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n566) );
NAND2_X1 MEM_stage_inst_dmem_U725 ( .A1(MEM_stage_inst_dmem_n564), .A2(MEM_stage_inst_dmem_n563), .ZN(MEM_stage_inst_dmem_n628) );
NOR2_X1 MEM_stage_inst_dmem_U724 ( .A1(MEM_stage_inst_dmem_n562), .A2(MEM_stage_inst_dmem_n561), .ZN(MEM_stage_inst_dmem_n563) );
NAND2_X1 MEM_stage_inst_dmem_U723 ( .A1(MEM_stage_inst_dmem_n560), .A2(MEM_stage_inst_dmem_n559), .ZN(MEM_stage_inst_dmem_n561) );
NOR2_X1 MEM_stage_inst_dmem_U722 ( .A1(MEM_stage_inst_dmem_n558), .A2(MEM_stage_inst_dmem_n557), .ZN(MEM_stage_inst_dmem_n559) );
NAND2_X1 MEM_stage_inst_dmem_U721 ( .A1(MEM_stage_inst_dmem_n556), .A2(MEM_stage_inst_dmem_n555), .ZN(MEM_stage_inst_dmem_n557) );
NAND2_X1 MEM_stage_inst_dmem_U720 ( .A1(MEM_stage_inst_dmem_ram_1568), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n555) );
NAND2_X1 MEM_stage_inst_dmem_U719 ( .A1(MEM_stage_inst_dmem_ram_1408), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n556) );
NAND2_X1 MEM_stage_inst_dmem_U718 ( .A1(MEM_stage_inst_dmem_n554), .A2(MEM_stage_inst_dmem_n553), .ZN(MEM_stage_inst_dmem_n558) );
NAND2_X1 MEM_stage_inst_dmem_U717 ( .A1(MEM_stage_inst_dmem_ram_1232), .A2(MEM_stage_inst_dmem_n51), .ZN(MEM_stage_inst_dmem_n553) );
NAND2_X1 MEM_stage_inst_dmem_U716 ( .A1(MEM_stage_inst_dmem_ram_1360), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n554) );
NOR2_X1 MEM_stage_inst_dmem_U715 ( .A1(MEM_stage_inst_dmem_n552), .A2(MEM_stage_inst_dmem_n551), .ZN(MEM_stage_inst_dmem_n560) );
NAND2_X1 MEM_stage_inst_dmem_U714 ( .A1(MEM_stage_inst_dmem_n550), .A2(MEM_stage_inst_dmem_n549), .ZN(MEM_stage_inst_dmem_n551) );
NAND2_X1 MEM_stage_inst_dmem_U713 ( .A1(MEM_stage_inst_dmem_ram_1344), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n549) );
NAND2_X1 MEM_stage_inst_dmem_U712 ( .A1(MEM_stage_inst_dmem_ram_1248), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n550) );
NAND2_X1 MEM_stage_inst_dmem_U711 ( .A1(MEM_stage_inst_dmem_n548), .A2(MEM_stage_inst_dmem_n547), .ZN(MEM_stage_inst_dmem_n552) );
NAND2_X1 MEM_stage_inst_dmem_U710 ( .A1(MEM_stage_inst_dmem_ram_1104), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n547) );
NAND2_X1 MEM_stage_inst_dmem_U709 ( .A1(MEM_stage_inst_dmem_ram_1200), .A2(MEM_stage_inst_dmem_n55), .ZN(MEM_stage_inst_dmem_n548) );
NAND2_X1 MEM_stage_inst_dmem_U708 ( .A1(MEM_stage_inst_dmem_n546), .A2(MEM_stage_inst_dmem_n545), .ZN(MEM_stage_inst_dmem_n562) );
NOR2_X1 MEM_stage_inst_dmem_U707 ( .A1(MEM_stage_inst_dmem_n544), .A2(MEM_stage_inst_dmem_n543), .ZN(MEM_stage_inst_dmem_n545) );
NAND2_X1 MEM_stage_inst_dmem_U706 ( .A1(MEM_stage_inst_dmem_n542), .A2(MEM_stage_inst_dmem_n541), .ZN(MEM_stage_inst_dmem_n543) );
NAND2_X1 MEM_stage_inst_dmem_U705 ( .A1(MEM_stage_inst_dmem_ram_1440), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n541) );
NAND2_X1 MEM_stage_inst_dmem_U704 ( .A1(MEM_stage_inst_dmem_ram_1840), .A2(MEM_stage_inst_dmem_n46), .ZN(MEM_stage_inst_dmem_n542) );
NAND2_X1 MEM_stage_inst_dmem_U703 ( .A1(MEM_stage_inst_dmem_n540), .A2(MEM_stage_inst_dmem_n539), .ZN(MEM_stage_inst_dmem_n544) );
NAND2_X1 MEM_stage_inst_dmem_U702 ( .A1(MEM_stage_inst_dmem_ram_1296), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n539) );
NAND2_X1 MEM_stage_inst_dmem_U701 ( .A1(MEM_stage_inst_dmem_ram_1744), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n540) );
NOR2_X1 MEM_stage_inst_dmem_U700 ( .A1(MEM_stage_inst_dmem_n538), .A2(MEM_stage_inst_dmem_n537), .ZN(MEM_stage_inst_dmem_n546) );
NAND2_X1 MEM_stage_inst_dmem_U699 ( .A1(MEM_stage_inst_dmem_n536), .A2(MEM_stage_inst_dmem_n535), .ZN(MEM_stage_inst_dmem_n537) );
NAND2_X1 MEM_stage_inst_dmem_U698 ( .A1(MEM_stage_inst_dmem_ram_1888), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n535) );
NAND2_X1 MEM_stage_inst_dmem_U697 ( .A1(MEM_stage_inst_dmem_ram_1648), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n536) );
NAND2_X1 MEM_stage_inst_dmem_U696 ( .A1(MEM_stage_inst_dmem_n534), .A2(MEM_stage_inst_dmem_n533), .ZN(MEM_stage_inst_dmem_n538) );
NAND2_X1 MEM_stage_inst_dmem_U695 ( .A1(MEM_stage_inst_dmem_ram_1472), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n533) );
NAND2_X1 MEM_stage_inst_dmem_U694 ( .A1(MEM_stage_inst_dmem_ram_1952), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n534) );
NOR2_X1 MEM_stage_inst_dmem_U693 ( .A1(MEM_stage_inst_dmem_n532), .A2(MEM_stage_inst_dmem_n531), .ZN(MEM_stage_inst_dmem_n564) );
NAND2_X1 MEM_stage_inst_dmem_U692 ( .A1(MEM_stage_inst_dmem_n530), .A2(MEM_stage_inst_dmem_n529), .ZN(MEM_stage_inst_dmem_n531) );
NOR2_X1 MEM_stage_inst_dmem_U691 ( .A1(MEM_stage_inst_dmem_n528), .A2(MEM_stage_inst_dmem_n527), .ZN(MEM_stage_inst_dmem_n529) );
NAND2_X1 MEM_stage_inst_dmem_U690 ( .A1(MEM_stage_inst_dmem_n526), .A2(MEM_stage_inst_dmem_n525), .ZN(MEM_stage_inst_dmem_n527) );
NAND2_X1 MEM_stage_inst_dmem_U689 ( .A1(MEM_stage_inst_dmem_ram_1856), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n525) );
NAND2_X1 MEM_stage_inst_dmem_U688 ( .A1(MEM_stage_inst_dmem_ram_1120), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n526) );
NAND2_X1 MEM_stage_inst_dmem_U687 ( .A1(MEM_stage_inst_dmem_n524), .A2(MEM_stage_inst_dmem_n523), .ZN(MEM_stage_inst_dmem_n528) );
NAND2_X1 MEM_stage_inst_dmem_U686 ( .A1(MEM_stage_inst_dmem_ram_1088), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n523) );
NAND2_X1 MEM_stage_inst_dmem_U685 ( .A1(MEM_stage_inst_dmem_ram_1392), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n524) );
NOR2_X1 MEM_stage_inst_dmem_U684 ( .A1(MEM_stage_inst_dmem_n522), .A2(MEM_stage_inst_dmem_n521), .ZN(MEM_stage_inst_dmem_n530) );
NAND2_X1 MEM_stage_inst_dmem_U683 ( .A1(MEM_stage_inst_dmem_n520), .A2(MEM_stage_inst_dmem_n519), .ZN(MEM_stage_inst_dmem_n521) );
NAND2_X1 MEM_stage_inst_dmem_U682 ( .A1(MEM_stage_inst_dmem_ram_1504), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n519) );
NAND2_X1 MEM_stage_inst_dmem_U681 ( .A1(MEM_stage_inst_dmem_ram_1824), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n520) );
NAND2_X1 MEM_stage_inst_dmem_U680 ( .A1(MEM_stage_inst_dmem_n518), .A2(MEM_stage_inst_dmem_n517), .ZN(MEM_stage_inst_dmem_n522) );
NAND2_X1 MEM_stage_inst_dmem_U679 ( .A1(MEM_stage_inst_dmem_ram_1984), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n517) );
NAND2_X1 MEM_stage_inst_dmem_U678 ( .A1(MEM_stage_inst_dmem_ram_1920), .A2(MEM_stage_inst_dmem_n72), .ZN(MEM_stage_inst_dmem_n518) );
NAND2_X1 MEM_stage_inst_dmem_U677 ( .A1(MEM_stage_inst_dmem_n516), .A2(MEM_stage_inst_dmem_n515), .ZN(MEM_stage_inst_dmem_n532) );
NOR2_X1 MEM_stage_inst_dmem_U676 ( .A1(MEM_stage_inst_dmem_n514), .A2(MEM_stage_inst_dmem_n513), .ZN(MEM_stage_inst_dmem_n515) );
NAND2_X1 MEM_stage_inst_dmem_U675 ( .A1(MEM_stage_inst_dmem_n512), .A2(MEM_stage_inst_dmem_n511), .ZN(MEM_stage_inst_dmem_n513) );
NAND2_X1 MEM_stage_inst_dmem_U674 ( .A1(MEM_stage_inst_dmem_ram_1072), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n511) );
NAND2_X1 MEM_stage_inst_dmem_U673 ( .A1(MEM_stage_inst_dmem_ram_1936), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n512) );
NAND2_X1 MEM_stage_inst_dmem_U672 ( .A1(MEM_stage_inst_dmem_n510), .A2(MEM_stage_inst_dmem_n509), .ZN(MEM_stage_inst_dmem_n514) );
NAND2_X1 MEM_stage_inst_dmem_U671 ( .A1(MEM_stage_inst_dmem_ram_1376), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n509) );
NAND2_X1 MEM_stage_inst_dmem_U670 ( .A1(MEM_stage_inst_dmem_ram_1136), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n510) );
NOR2_X1 MEM_stage_inst_dmem_U669 ( .A1(MEM_stage_inst_dmem_n508), .A2(MEM_stage_inst_dmem_n507), .ZN(MEM_stage_inst_dmem_n516) );
NAND2_X1 MEM_stage_inst_dmem_U668 ( .A1(MEM_stage_inst_dmem_n506), .A2(MEM_stage_inst_dmem_n505), .ZN(MEM_stage_inst_dmem_n507) );
NAND2_X1 MEM_stage_inst_dmem_U667 ( .A1(MEM_stage_inst_dmem_ram_1872), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n505) );
NAND2_X1 MEM_stage_inst_dmem_U666 ( .A1(MEM_stage_inst_dmem_ram_1616), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n506) );
NAND2_X1 MEM_stage_inst_dmem_U665 ( .A1(MEM_stage_inst_dmem_n504), .A2(MEM_stage_inst_dmem_n503), .ZN(MEM_stage_inst_dmem_n508) );
NAND2_X1 MEM_stage_inst_dmem_U664 ( .A1(MEM_stage_inst_dmem_ram_1456), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n503) );
NAND2_X1 MEM_stage_inst_dmem_U663 ( .A1(MEM_stage_inst_dmem_ram_2016), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n504) );
NOR2_X1 MEM_stage_inst_dmem_U662 ( .A1(MEM_stage_inst_dmem_n502), .A2(MEM_stage_inst_dmem_n501), .ZN(MEM_stage_inst_dmem_n760) );
NOR2_X1 MEM_stage_inst_dmem_U661 ( .A1(MEM_stage_inst_dmem_n500), .A2(MEM_stage_inst_dmem_n8286), .ZN(MEM_stage_inst_dmem_n501) );
OR2_X1 MEM_stage_inst_dmem_U660 ( .A1(MEM_stage_inst_dmem_n15967), .A2(EX_pipeline_reg_out_29), .ZN(MEM_stage_inst_dmem_n8286) );
INV_X1 MEM_stage_inst_dmem_U659 ( .A(EX_pipeline_reg_out_28), .ZN(MEM_stage_inst_dmem_n15967) );
NOR2_X1 MEM_stage_inst_dmem_U658 ( .A1(MEM_stage_inst_dmem_n499), .A2(MEM_stage_inst_dmem_n498), .ZN(MEM_stage_inst_dmem_n500) );
NAND2_X1 MEM_stage_inst_dmem_U657 ( .A1(MEM_stage_inst_dmem_n497), .A2(MEM_stage_inst_dmem_n496), .ZN(MEM_stage_inst_dmem_n498) );
NOR2_X1 MEM_stage_inst_dmem_U656 ( .A1(MEM_stage_inst_dmem_n495), .A2(MEM_stage_inst_dmem_n494), .ZN(MEM_stage_inst_dmem_n496) );
NAND2_X1 MEM_stage_inst_dmem_U655 ( .A1(MEM_stage_inst_dmem_n493), .A2(MEM_stage_inst_dmem_n492), .ZN(MEM_stage_inst_dmem_n494) );
NOR2_X1 MEM_stage_inst_dmem_U654 ( .A1(MEM_stage_inst_dmem_n491), .A2(MEM_stage_inst_dmem_n490), .ZN(MEM_stage_inst_dmem_n492) );
NAND2_X1 MEM_stage_inst_dmem_U653 ( .A1(MEM_stage_inst_dmem_n489), .A2(MEM_stage_inst_dmem_n488), .ZN(MEM_stage_inst_dmem_n490) );
NAND2_X1 MEM_stage_inst_dmem_U652 ( .A1(MEM_stage_inst_dmem_ram_2768), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n488) );
NAND2_X1 MEM_stage_inst_dmem_U651 ( .A1(MEM_stage_inst_dmem_ram_2704), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n489) );
NAND2_X1 MEM_stage_inst_dmem_U650 ( .A1(MEM_stage_inst_dmem_n487), .A2(MEM_stage_inst_dmem_n486), .ZN(MEM_stage_inst_dmem_n491) );
NAND2_X1 MEM_stage_inst_dmem_U649 ( .A1(MEM_stage_inst_dmem_ram_2544), .A2(MEM_stage_inst_dmem_n8535), .ZN(MEM_stage_inst_dmem_n486) );
NAND2_X1 MEM_stage_inst_dmem_U648 ( .A1(MEM_stage_inst_dmem_ram_2592), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n487) );
NOR2_X1 MEM_stage_inst_dmem_U647 ( .A1(MEM_stage_inst_dmem_n485), .A2(MEM_stage_inst_dmem_n484), .ZN(MEM_stage_inst_dmem_n493) );
NAND2_X1 MEM_stage_inst_dmem_U646 ( .A1(MEM_stage_inst_dmem_n483), .A2(MEM_stage_inst_dmem_n482), .ZN(MEM_stage_inst_dmem_n484) );
NAND2_X1 MEM_stage_inst_dmem_U645 ( .A1(MEM_stage_inst_dmem_ram_2608), .A2(MEM_stage_inst_dmem_n41), .ZN(MEM_stage_inst_dmem_n482) );
NAND2_X1 MEM_stage_inst_dmem_U644 ( .A1(MEM_stage_inst_dmem_ram_2192), .A2(MEM_stage_inst_dmem_n5807), .ZN(MEM_stage_inst_dmem_n483) );
BUF_X1 MEM_stage_inst_dmem_U643 ( .A(MEM_stage_inst_dmem_n7903), .Z(MEM_stage_inst_dmem_n5807) );
NAND2_X1 MEM_stage_inst_dmem_U642 ( .A1(MEM_stage_inst_dmem_n481), .A2(MEM_stage_inst_dmem_n480), .ZN(MEM_stage_inst_dmem_n485) );
NAND2_X1 MEM_stage_inst_dmem_U641 ( .A1(MEM_stage_inst_dmem_ram_2448), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n480) );
NAND2_X1 MEM_stage_inst_dmem_U640 ( .A1(MEM_stage_inst_dmem_ram_3056), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n481) );
NAND2_X1 MEM_stage_inst_dmem_U639 ( .A1(MEM_stage_inst_dmem_n479), .A2(MEM_stage_inst_dmem_n478), .ZN(MEM_stage_inst_dmem_n495) );
NOR2_X1 MEM_stage_inst_dmem_U638 ( .A1(MEM_stage_inst_dmem_n477), .A2(MEM_stage_inst_dmem_n476), .ZN(MEM_stage_inst_dmem_n478) );
NAND2_X1 MEM_stage_inst_dmem_U637 ( .A1(MEM_stage_inst_dmem_n475), .A2(MEM_stage_inst_dmem_n474), .ZN(MEM_stage_inst_dmem_n476) );
NAND2_X1 MEM_stage_inst_dmem_U636 ( .A1(MEM_stage_inst_dmem_ram_2736), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n474) );
NAND2_X1 MEM_stage_inst_dmem_U635 ( .A1(MEM_stage_inst_dmem_ram_2832), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n475) );
NAND2_X1 MEM_stage_inst_dmem_U634 ( .A1(MEM_stage_inst_dmem_n473), .A2(MEM_stage_inst_dmem_n472), .ZN(MEM_stage_inst_dmem_n477) );
NAND2_X1 MEM_stage_inst_dmem_U633 ( .A1(MEM_stage_inst_dmem_ram_2976), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n472) );
NAND2_X1 MEM_stage_inst_dmem_U632 ( .A1(MEM_stage_inst_dmem_ram_2224), .A2(MEM_stage_inst_dmem_n55), .ZN(MEM_stage_inst_dmem_n473) );
NOR2_X1 MEM_stage_inst_dmem_U631 ( .A1(MEM_stage_inst_dmem_n471), .A2(MEM_stage_inst_dmem_n470), .ZN(MEM_stage_inst_dmem_n479) );
NAND2_X1 MEM_stage_inst_dmem_U630 ( .A1(MEM_stage_inst_dmem_n469), .A2(MEM_stage_inst_dmem_n468), .ZN(MEM_stage_inst_dmem_n470) );
NAND2_X1 MEM_stage_inst_dmem_U629 ( .A1(MEM_stage_inst_dmem_ram_2992), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n468) );
NAND2_X1 MEM_stage_inst_dmem_U628 ( .A1(MEM_stage_inst_dmem_ram_2112), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n469) );
NAND2_X1 MEM_stage_inst_dmem_U627 ( .A1(MEM_stage_inst_dmem_n467), .A2(MEM_stage_inst_dmem_n466), .ZN(MEM_stage_inst_dmem_n471) );
NAND2_X1 MEM_stage_inst_dmem_U626 ( .A1(MEM_stage_inst_dmem_ram_2176), .A2(MEM_stage_inst_dmem_n61), .ZN(MEM_stage_inst_dmem_n466) );
NAND2_X1 MEM_stage_inst_dmem_U625 ( .A1(MEM_stage_inst_dmem_ram_2512), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n467) );
NOR2_X1 MEM_stage_inst_dmem_U624 ( .A1(MEM_stage_inst_dmem_n465), .A2(MEM_stage_inst_dmem_n464), .ZN(MEM_stage_inst_dmem_n497) );
NAND2_X1 MEM_stage_inst_dmem_U623 ( .A1(MEM_stage_inst_dmem_n463), .A2(MEM_stage_inst_dmem_n462), .ZN(MEM_stage_inst_dmem_n464) );
NOR2_X1 MEM_stage_inst_dmem_U622 ( .A1(MEM_stage_inst_dmem_n461), .A2(MEM_stage_inst_dmem_n460), .ZN(MEM_stage_inst_dmem_n462) );
NAND2_X1 MEM_stage_inst_dmem_U621 ( .A1(MEM_stage_inst_dmem_n459), .A2(MEM_stage_inst_dmem_n458), .ZN(MEM_stage_inst_dmem_n460) );
NAND2_X1 MEM_stage_inst_dmem_U620 ( .A1(MEM_stage_inst_dmem_ram_2800), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n458) );
NAND2_X1 MEM_stage_inst_dmem_U619 ( .A1(MEM_stage_inst_dmem_ram_2496), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n459) );
NAND2_X1 MEM_stage_inst_dmem_U618 ( .A1(MEM_stage_inst_dmem_n457), .A2(MEM_stage_inst_dmem_n456), .ZN(MEM_stage_inst_dmem_n461) );
NAND2_X1 MEM_stage_inst_dmem_U617 ( .A1(MEM_stage_inst_dmem_ram_2960), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n456) );
NAND2_X1 MEM_stage_inst_dmem_U616 ( .A1(MEM_stage_inst_dmem_ram_2208), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n457) );
NOR2_X1 MEM_stage_inst_dmem_U615 ( .A1(MEM_stage_inst_dmem_n455), .A2(MEM_stage_inst_dmem_n454), .ZN(MEM_stage_inst_dmem_n463) );
NAND2_X1 MEM_stage_inst_dmem_U614 ( .A1(MEM_stage_inst_dmem_n453), .A2(MEM_stage_inst_dmem_n452), .ZN(MEM_stage_inst_dmem_n454) );
NAND2_X1 MEM_stage_inst_dmem_U613 ( .A1(MEM_stage_inst_dmem_ram_2464), .A2(MEM_stage_inst_dmem_n4772), .ZN(MEM_stage_inst_dmem_n452) );
NAND2_X1 MEM_stage_inst_dmem_U612 ( .A1(MEM_stage_inst_dmem_ram_2640), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n453) );
NAND2_X1 MEM_stage_inst_dmem_U611 ( .A1(MEM_stage_inst_dmem_n451), .A2(MEM_stage_inst_dmem_n450), .ZN(MEM_stage_inst_dmem_n455) );
NAND2_X1 MEM_stage_inst_dmem_U610 ( .A1(MEM_stage_inst_dmem_ram_2880), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n450) );
NAND2_X1 MEM_stage_inst_dmem_U609 ( .A1(MEM_stage_inst_dmem_ram_2416), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n451) );
NAND2_X1 MEM_stage_inst_dmem_U608 ( .A1(MEM_stage_inst_dmem_n449), .A2(MEM_stage_inst_dmem_n448), .ZN(MEM_stage_inst_dmem_n465) );
NOR2_X1 MEM_stage_inst_dmem_U607 ( .A1(MEM_stage_inst_dmem_n447), .A2(MEM_stage_inst_dmem_n446), .ZN(MEM_stage_inst_dmem_n448) );
NAND2_X1 MEM_stage_inst_dmem_U606 ( .A1(MEM_stage_inst_dmem_n445), .A2(MEM_stage_inst_dmem_n444), .ZN(MEM_stage_inst_dmem_n446) );
NAND2_X1 MEM_stage_inst_dmem_U605 ( .A1(MEM_stage_inst_dmem_ram_2256), .A2(MEM_stage_inst_dmem_n51), .ZN(MEM_stage_inst_dmem_n444) );
NAND2_X1 MEM_stage_inst_dmem_U604 ( .A1(MEM_stage_inst_dmem_ram_2048), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n445) );
NAND2_X1 MEM_stage_inst_dmem_U603 ( .A1(MEM_stage_inst_dmem_n443), .A2(MEM_stage_inst_dmem_n442), .ZN(MEM_stage_inst_dmem_n447) );
NAND2_X1 MEM_stage_inst_dmem_U602 ( .A1(MEM_stage_inst_dmem_ram_2576), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n442) );
NAND2_X1 MEM_stage_inst_dmem_U601 ( .A1(MEM_stage_inst_dmem_ram_2304), .A2(MEM_stage_inst_dmem_n5857), .ZN(MEM_stage_inst_dmem_n443) );
NOR2_X1 MEM_stage_inst_dmem_U600 ( .A1(MEM_stage_inst_dmem_n441), .A2(MEM_stage_inst_dmem_n440), .ZN(MEM_stage_inst_dmem_n449) );
NAND2_X1 MEM_stage_inst_dmem_U599 ( .A1(MEM_stage_inst_dmem_n439), .A2(MEM_stage_inst_dmem_n438), .ZN(MEM_stage_inst_dmem_n440) );
NAND2_X1 MEM_stage_inst_dmem_U598 ( .A1(MEM_stage_inst_dmem_ram_2368), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n438) );
NAND2_X1 MEM_stage_inst_dmem_U597 ( .A1(MEM_stage_inst_dmem_ram_2272), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n439) );
NAND2_X1 MEM_stage_inst_dmem_U596 ( .A1(MEM_stage_inst_dmem_n437), .A2(MEM_stage_inst_dmem_n436), .ZN(MEM_stage_inst_dmem_n441) );
NAND2_X1 MEM_stage_inst_dmem_U595 ( .A1(MEM_stage_inst_dmem_ram_2080), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n436) );
NAND2_X1 MEM_stage_inst_dmem_U594 ( .A1(MEM_stage_inst_dmem_ram_2384), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n437) );
NAND2_X1 MEM_stage_inst_dmem_U593 ( .A1(MEM_stage_inst_dmem_n435), .A2(MEM_stage_inst_dmem_n434), .ZN(MEM_stage_inst_dmem_n499) );
NOR2_X1 MEM_stage_inst_dmem_U592 ( .A1(MEM_stage_inst_dmem_n433), .A2(MEM_stage_inst_dmem_n432), .ZN(MEM_stage_inst_dmem_n434) );
NAND2_X1 MEM_stage_inst_dmem_U591 ( .A1(MEM_stage_inst_dmem_n431), .A2(MEM_stage_inst_dmem_n430), .ZN(MEM_stage_inst_dmem_n432) );
NOR2_X1 MEM_stage_inst_dmem_U590 ( .A1(MEM_stage_inst_dmem_n429), .A2(MEM_stage_inst_dmem_n428), .ZN(MEM_stage_inst_dmem_n430) );
NAND2_X1 MEM_stage_inst_dmem_U589 ( .A1(MEM_stage_inst_dmem_n427), .A2(MEM_stage_inst_dmem_n426), .ZN(MEM_stage_inst_dmem_n428) );
NAND2_X1 MEM_stage_inst_dmem_U588 ( .A1(MEM_stage_inst_dmem_ram_2480), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n426) );
NAND2_X1 MEM_stage_inst_dmem_U587 ( .A1(MEM_stage_inst_dmem_ram_2144), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n427) );
NAND2_X1 MEM_stage_inst_dmem_U586 ( .A1(MEM_stage_inst_dmem_n425), .A2(MEM_stage_inst_dmem_n424), .ZN(MEM_stage_inst_dmem_n429) );
NAND2_X1 MEM_stage_inst_dmem_U585 ( .A1(MEM_stage_inst_dmem_ram_2912), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n424) );
NAND2_X1 MEM_stage_inst_dmem_U584 ( .A1(MEM_stage_inst_dmem_ram_2752), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n425) );
NOR2_X1 MEM_stage_inst_dmem_U583 ( .A1(MEM_stage_inst_dmem_n423), .A2(MEM_stage_inst_dmem_n422), .ZN(MEM_stage_inst_dmem_n431) );
NAND2_X1 MEM_stage_inst_dmem_U582 ( .A1(MEM_stage_inst_dmem_n421), .A2(MEM_stage_inst_dmem_n420), .ZN(MEM_stage_inst_dmem_n422) );
NAND2_X1 MEM_stage_inst_dmem_U581 ( .A1(MEM_stage_inst_dmem_ram_2400), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n420) );
NAND2_X1 MEM_stage_inst_dmem_U580 ( .A1(MEM_stage_inst_dmem_ram_2336), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n421) );
NAND2_X1 MEM_stage_inst_dmem_U579 ( .A1(MEM_stage_inst_dmem_n419), .A2(MEM_stage_inst_dmem_n418), .ZN(MEM_stage_inst_dmem_n423) );
NAND2_X1 MEM_stage_inst_dmem_U578 ( .A1(MEM_stage_inst_dmem_ram_2528), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n418) );
NAND2_X1 MEM_stage_inst_dmem_U577 ( .A1(MEM_stage_inst_dmem_ram_2320), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n419) );
NAND2_X1 MEM_stage_inst_dmem_U576 ( .A1(MEM_stage_inst_dmem_n417), .A2(MEM_stage_inst_dmem_n416), .ZN(MEM_stage_inst_dmem_n433) );
NOR2_X1 MEM_stage_inst_dmem_U575 ( .A1(MEM_stage_inst_dmem_n415), .A2(MEM_stage_inst_dmem_n414), .ZN(MEM_stage_inst_dmem_n416) );
NAND2_X1 MEM_stage_inst_dmem_U574 ( .A1(MEM_stage_inst_dmem_n413), .A2(MEM_stage_inst_dmem_n412), .ZN(MEM_stage_inst_dmem_n414) );
NAND2_X1 MEM_stage_inst_dmem_U573 ( .A1(MEM_stage_inst_dmem_ram_2688), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n412) );
NAND2_X1 MEM_stage_inst_dmem_U572 ( .A1(MEM_stage_inst_dmem_ram_2864), .A2(MEM_stage_inst_dmem_n8005), .ZN(MEM_stage_inst_dmem_n413) );
BUF_X1 MEM_stage_inst_dmem_U571 ( .A(MEM_stage_inst_dmem_n4740), .Z(MEM_stage_inst_dmem_n8005) );
NAND2_X1 MEM_stage_inst_dmem_U570 ( .A1(MEM_stage_inst_dmem_n411), .A2(MEM_stage_inst_dmem_n410), .ZN(MEM_stage_inst_dmem_n415) );
NAND2_X1 MEM_stage_inst_dmem_U569 ( .A1(MEM_stage_inst_dmem_ram_2096), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n410) );
NAND2_X1 MEM_stage_inst_dmem_U568 ( .A1(MEM_stage_inst_dmem_ram_2128), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n411) );
NOR2_X1 MEM_stage_inst_dmem_U567 ( .A1(MEM_stage_inst_dmem_n409), .A2(MEM_stage_inst_dmem_n408), .ZN(MEM_stage_inst_dmem_n417) );
NAND2_X1 MEM_stage_inst_dmem_U566 ( .A1(MEM_stage_inst_dmem_n407), .A2(MEM_stage_inst_dmem_n406), .ZN(MEM_stage_inst_dmem_n408) );
NAND2_X1 MEM_stage_inst_dmem_U565 ( .A1(MEM_stage_inst_dmem_ram_2720), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n406) );
NAND2_X1 MEM_stage_inst_dmem_U564 ( .A1(MEM_stage_inst_dmem_ram_2064), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n407) );
NAND2_X1 MEM_stage_inst_dmem_U563 ( .A1(MEM_stage_inst_dmem_n405), .A2(MEM_stage_inst_dmem_n404), .ZN(MEM_stage_inst_dmem_n409) );
NAND2_X1 MEM_stage_inst_dmem_U562 ( .A1(MEM_stage_inst_dmem_ram_2656), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n404) );
NAND2_X1 MEM_stage_inst_dmem_U561 ( .A1(MEM_stage_inst_dmem_ram_2624), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n405) );
NOR2_X1 MEM_stage_inst_dmem_U560 ( .A1(MEM_stage_inst_dmem_n403), .A2(MEM_stage_inst_dmem_n402), .ZN(MEM_stage_inst_dmem_n435) );
NAND2_X1 MEM_stage_inst_dmem_U559 ( .A1(MEM_stage_inst_dmem_n401), .A2(MEM_stage_inst_dmem_n400), .ZN(MEM_stage_inst_dmem_n402) );
NOR2_X1 MEM_stage_inst_dmem_U558 ( .A1(MEM_stage_inst_dmem_n399), .A2(MEM_stage_inst_dmem_n398), .ZN(MEM_stage_inst_dmem_n400) );
NAND2_X1 MEM_stage_inst_dmem_U557 ( .A1(MEM_stage_inst_dmem_n397), .A2(MEM_stage_inst_dmem_n396), .ZN(MEM_stage_inst_dmem_n398) );
NAND2_X1 MEM_stage_inst_dmem_U556 ( .A1(MEM_stage_inst_dmem_ram_3040), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n396) );
NAND2_X1 MEM_stage_inst_dmem_U555 ( .A1(MEM_stage_inst_dmem_ram_2784), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n397) );
NAND2_X1 MEM_stage_inst_dmem_U554 ( .A1(MEM_stage_inst_dmem_n395), .A2(MEM_stage_inst_dmem_n394), .ZN(MEM_stage_inst_dmem_n399) );
NAND2_X1 MEM_stage_inst_dmem_U553 ( .A1(MEM_stage_inst_dmem_ram_2928), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n394) );
NAND2_X1 MEM_stage_inst_dmem_U552 ( .A1(MEM_stage_inst_dmem_ram_2672), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n395) );
NOR2_X1 MEM_stage_inst_dmem_U551 ( .A1(MEM_stage_inst_dmem_n393), .A2(MEM_stage_inst_dmem_n392), .ZN(MEM_stage_inst_dmem_n401) );
NAND2_X1 MEM_stage_inst_dmem_U550 ( .A1(MEM_stage_inst_dmem_n391), .A2(MEM_stage_inst_dmem_n390), .ZN(MEM_stage_inst_dmem_n392) );
NAND2_X1 MEM_stage_inst_dmem_U549 ( .A1(MEM_stage_inst_dmem_ram_2944), .A2(MEM_stage_inst_dmem_n72), .ZN(MEM_stage_inst_dmem_n390) );
NAND2_X1 MEM_stage_inst_dmem_U548 ( .A1(MEM_stage_inst_dmem_ram_2560), .A2(MEM_stage_inst_dmem_n71), .ZN(MEM_stage_inst_dmem_n391) );
NAND2_X1 MEM_stage_inst_dmem_U547 ( .A1(MEM_stage_inst_dmem_n389), .A2(MEM_stage_inst_dmem_n388), .ZN(MEM_stage_inst_dmem_n393) );
NAND2_X1 MEM_stage_inst_dmem_U546 ( .A1(MEM_stage_inst_dmem_ram_3008), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n388) );
NAND2_X1 MEM_stage_inst_dmem_U545 ( .A1(MEM_stage_inst_dmem_ram_2288), .A2(MEM_stage_inst_dmem_n7914), .ZN(MEM_stage_inst_dmem_n389) );
BUF_X1 MEM_stage_inst_dmem_U544 ( .A(MEM_stage_inst_dmem_n4649), .Z(MEM_stage_inst_dmem_n7914) );
NAND2_X1 MEM_stage_inst_dmem_U543 ( .A1(MEM_stage_inst_dmem_n387), .A2(MEM_stage_inst_dmem_n386), .ZN(MEM_stage_inst_dmem_n403) );
NOR2_X1 MEM_stage_inst_dmem_U542 ( .A1(MEM_stage_inst_dmem_n385), .A2(MEM_stage_inst_dmem_n384), .ZN(MEM_stage_inst_dmem_n386) );
NAND2_X1 MEM_stage_inst_dmem_U541 ( .A1(MEM_stage_inst_dmem_n383), .A2(MEM_stage_inst_dmem_n382), .ZN(MEM_stage_inst_dmem_n384) );
NAND2_X1 MEM_stage_inst_dmem_U540 ( .A1(MEM_stage_inst_dmem_ram_2240), .A2(MEM_stage_inst_dmem_n36), .ZN(MEM_stage_inst_dmem_n382) );
NAND2_X1 MEM_stage_inst_dmem_U539 ( .A1(MEM_stage_inst_dmem_ram_2352), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n383) );
NAND2_X1 MEM_stage_inst_dmem_U538 ( .A1(MEM_stage_inst_dmem_n381), .A2(MEM_stage_inst_dmem_n380), .ZN(MEM_stage_inst_dmem_n385) );
NAND2_X1 MEM_stage_inst_dmem_U537 ( .A1(MEM_stage_inst_dmem_ram_3024), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n380) );
NAND2_X1 MEM_stage_inst_dmem_U536 ( .A1(MEM_stage_inst_dmem_ram_2848), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n381) );
NOR2_X1 MEM_stage_inst_dmem_U535 ( .A1(MEM_stage_inst_dmem_n379), .A2(MEM_stage_inst_dmem_n378), .ZN(MEM_stage_inst_dmem_n387) );
NAND2_X1 MEM_stage_inst_dmem_U534 ( .A1(MEM_stage_inst_dmem_n377), .A2(MEM_stage_inst_dmem_n376), .ZN(MEM_stage_inst_dmem_n378) );
NAND2_X1 MEM_stage_inst_dmem_U533 ( .A1(MEM_stage_inst_dmem_ram_2896), .A2(MEM_stage_inst_dmem_n8372), .ZN(MEM_stage_inst_dmem_n376) );
NAND2_X1 MEM_stage_inst_dmem_U532 ( .A1(MEM_stage_inst_dmem_ram_2160), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n377) );
NAND2_X1 MEM_stage_inst_dmem_U531 ( .A1(MEM_stage_inst_dmem_n375), .A2(MEM_stage_inst_dmem_n374), .ZN(MEM_stage_inst_dmem_n379) );
NAND2_X1 MEM_stage_inst_dmem_U530 ( .A1(MEM_stage_inst_dmem_ram_2816), .A2(MEM_stage_inst_dmem_n37), .ZN(MEM_stage_inst_dmem_n374) );
NAND2_X1 MEM_stage_inst_dmem_U529 ( .A1(MEM_stage_inst_dmem_ram_2432), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n375) );
NOR2_X1 MEM_stage_inst_dmem_U528 ( .A1(MEM_stage_inst_dmem_n373), .A2(MEM_stage_inst_dmem_n8551), .ZN(MEM_stage_inst_dmem_n502) );
NAND2_X1 MEM_stage_inst_dmem_U527 ( .A1(EX_pipeline_reg_out_28), .A2(EX_pipeline_reg_out_29), .ZN(MEM_stage_inst_dmem_n8551) );
NOR2_X1 MEM_stage_inst_dmem_U526 ( .A1(MEM_stage_inst_dmem_n372), .A2(MEM_stage_inst_dmem_n371), .ZN(MEM_stage_inst_dmem_n373) );
NAND2_X1 MEM_stage_inst_dmem_U525 ( .A1(MEM_stage_inst_dmem_n370), .A2(MEM_stage_inst_dmem_n369), .ZN(MEM_stage_inst_dmem_n371) );
NOR2_X1 MEM_stage_inst_dmem_U524 ( .A1(MEM_stage_inst_dmem_n368), .A2(MEM_stage_inst_dmem_n367), .ZN(MEM_stage_inst_dmem_n369) );
NAND2_X1 MEM_stage_inst_dmem_U523 ( .A1(MEM_stage_inst_dmem_n366), .A2(MEM_stage_inst_dmem_n365), .ZN(MEM_stage_inst_dmem_n367) );
NOR2_X1 MEM_stage_inst_dmem_U522 ( .A1(MEM_stage_inst_dmem_n364), .A2(MEM_stage_inst_dmem_n363), .ZN(MEM_stage_inst_dmem_n365) );
NAND2_X1 MEM_stage_inst_dmem_U521 ( .A1(MEM_stage_inst_dmem_n362), .A2(MEM_stage_inst_dmem_n361), .ZN(MEM_stage_inst_dmem_n363) );
NAND2_X1 MEM_stage_inst_dmem_U520 ( .A1(MEM_stage_inst_dmem_ram_640), .A2(MEM_stage_inst_dmem_n49), .ZN(MEM_stage_inst_dmem_n361) );
NOR2_X1 MEM_stage_inst_dmem_U519 ( .A1(MEM_stage_inst_dmem_n360), .A2(MEM_stage_inst_dmem_n359), .ZN(MEM_stage_inst_dmem_n7960) );
NAND2_X1 MEM_stage_inst_dmem_U518 ( .A1(MEM_stage_inst_dmem_ram_16), .A2(MEM_stage_inst_dmem_n70), .ZN(MEM_stage_inst_dmem_n362) );
NOR2_X1 MEM_stage_inst_dmem_U517 ( .A1(MEM_stage_inst_dmem_n358), .A2(MEM_stage_inst_dmem_n357), .ZN(MEM_stage_inst_dmem_n7887) );
NAND2_X1 MEM_stage_inst_dmem_U516 ( .A1(MEM_stage_inst_dmem_n356), .A2(MEM_stage_inst_dmem_n355), .ZN(MEM_stage_inst_dmem_n364) );
NAND2_X1 MEM_stage_inst_dmem_U515 ( .A1(MEM_stage_inst_dmem_ram_704), .A2(MEM_stage_inst_dmem_n59), .ZN(MEM_stage_inst_dmem_n355) );
NOR2_X1 MEM_stage_inst_dmem_U514 ( .A1(MEM_stage_inst_dmem_n354), .A2(MEM_stage_inst_dmem_n359), .ZN(MEM_stage_inst_dmem_n3192) );
NAND2_X1 MEM_stage_inst_dmem_U513 ( .A1(MEM_stage_inst_dmem_ram_128), .A2(MEM_stage_inst_dmem_n61), .ZN(MEM_stage_inst_dmem_n356) );
NOR2_X1 MEM_stage_inst_dmem_U512 ( .A1(MEM_stage_inst_dmem_n353), .A2(MEM_stage_inst_dmem_n360), .ZN(MEM_stage_inst_dmem_n3130) );
NOR2_X1 MEM_stage_inst_dmem_U511 ( .A1(MEM_stage_inst_dmem_n352), .A2(MEM_stage_inst_dmem_n351), .ZN(MEM_stage_inst_dmem_n366) );
NAND2_X1 MEM_stage_inst_dmem_U510 ( .A1(MEM_stage_inst_dmem_n350), .A2(MEM_stage_inst_dmem_n349), .ZN(MEM_stage_inst_dmem_n351) );
NAND2_X1 MEM_stage_inst_dmem_U509 ( .A1(MEM_stage_inst_dmem_ram_192), .A2(MEM_stage_inst_dmem_n36), .ZN(MEM_stage_inst_dmem_n349) );
NOR2_X1 MEM_stage_inst_dmem_U508 ( .A1(MEM_stage_inst_dmem_n353), .A2(MEM_stage_inst_dmem_n354), .ZN(MEM_stage_inst_dmem_n3082) );
NAND2_X1 MEM_stage_inst_dmem_U507 ( .A1(MEM_stage_inst_dmem_ram_336), .A2(MEM_stage_inst_dmem_n8451), .ZN(MEM_stage_inst_dmem_n350) );
BUF_X2 MEM_stage_inst_dmem_U506 ( .A(MEM_stage_inst_dmem_n3216), .Z(MEM_stage_inst_dmem_n8451) );
NAND2_X1 MEM_stage_inst_dmem_U505 ( .A1(MEM_stage_inst_dmem_n346), .A2(MEM_stage_inst_dmem_n345), .ZN(MEM_stage_inst_dmem_n352) );
NAND2_X1 MEM_stage_inst_dmem_U504 ( .A1(MEM_stage_inst_dmem_ram_320), .A2(MEM_stage_inst_dmem_n66), .ZN(MEM_stage_inst_dmem_n345) );
NOR2_X1 MEM_stage_inst_dmem_U503 ( .A1(MEM_stage_inst_dmem_n354), .A2(MEM_stage_inst_dmem_n348), .ZN(MEM_stage_inst_dmem_n4706) );
NAND2_X1 MEM_stage_inst_dmem_U502 ( .A1(MEM_stage_inst_dmem_ram_912), .A2(MEM_stage_inst_dmem_n24), .ZN(MEM_stage_inst_dmem_n346) );
NOR2_X1 MEM_stage_inst_dmem_U501 ( .A1(MEM_stage_inst_dmem_n357), .A2(MEM_stage_inst_dmem_n344), .ZN(MEM_stage_inst_dmem_n3073) );
NAND2_X1 MEM_stage_inst_dmem_U500 ( .A1(MEM_stage_inst_dmem_n343), .A2(MEM_stage_inst_dmem_n342), .ZN(MEM_stage_inst_dmem_n368) );
NOR2_X1 MEM_stage_inst_dmem_U499 ( .A1(MEM_stage_inst_dmem_n341), .A2(MEM_stage_inst_dmem_n340), .ZN(MEM_stage_inst_dmem_n342) );
NAND2_X1 MEM_stage_inst_dmem_U498 ( .A1(MEM_stage_inst_dmem_n339), .A2(MEM_stage_inst_dmem_n338), .ZN(MEM_stage_inst_dmem_n340) );
NAND2_X1 MEM_stage_inst_dmem_U497 ( .A1(MEM_stage_inst_dmem_ram_992), .A2(MEM_stage_inst_dmem_n47), .ZN(MEM_stage_inst_dmem_n338) );
NOR2_X1 MEM_stage_inst_dmem_U496 ( .A1(MEM_stage_inst_dmem_n337), .A2(MEM_stage_inst_dmem_n344), .ZN(MEM_stage_inst_dmem_n3113) );
NAND2_X1 MEM_stage_inst_dmem_U495 ( .A1(MEM_stage_inst_dmem_ram_112), .A2(MEM_stage_inst_dmem_n52), .ZN(MEM_stage_inst_dmem_n339) );
NOR2_X1 MEM_stage_inst_dmem_U494 ( .A1(MEM_stage_inst_dmem_n336), .A2(MEM_stage_inst_dmem_n358), .ZN(MEM_stage_inst_dmem_n4710) );
NAND2_X1 MEM_stage_inst_dmem_U493 ( .A1(MEM_stage_inst_dmem_n335), .A2(MEM_stage_inst_dmem_n334), .ZN(MEM_stage_inst_dmem_n341) );
NAND2_X1 MEM_stage_inst_dmem_U492 ( .A1(MEM_stage_inst_dmem_ram_352), .A2(MEM_stage_inst_dmem_n25), .ZN(MEM_stage_inst_dmem_n334) );
NOR2_X1 MEM_stage_inst_dmem_U491 ( .A1(MEM_stage_inst_dmem_n337), .A2(MEM_stage_inst_dmem_n348), .ZN(MEM_stage_inst_dmem_n3217) );
NAND2_X1 MEM_stage_inst_dmem_U490 ( .A1(MEM_stage_inst_dmem_ram_176), .A2(MEM_stage_inst_dmem_n8434), .ZN(MEM_stage_inst_dmem_n335) );
BUF_X1 MEM_stage_inst_dmem_U489 ( .A(MEM_stage_inst_dmem_n7937), .Z(MEM_stage_inst_dmem_n8434) );
NOR2_X1 MEM_stage_inst_dmem_U488 ( .A1(MEM_stage_inst_dmem_n353), .A2(MEM_stage_inst_dmem_n333), .ZN(MEM_stage_inst_dmem_n7937) );
NOR2_X1 MEM_stage_inst_dmem_U487 ( .A1(MEM_stage_inst_dmem_n332), .A2(MEM_stage_inst_dmem_n331), .ZN(MEM_stage_inst_dmem_n343) );
NAND2_X1 MEM_stage_inst_dmem_U486 ( .A1(MEM_stage_inst_dmem_n330), .A2(MEM_stage_inst_dmem_n329), .ZN(MEM_stage_inst_dmem_n331) );
NAND2_X1 MEM_stage_inst_dmem_U485 ( .A1(MEM_stage_inst_dmem_ram_864), .A2(MEM_stage_inst_dmem_n63), .ZN(MEM_stage_inst_dmem_n329) );
NOR2_X1 MEM_stage_inst_dmem_U484 ( .A1(MEM_stage_inst_dmem_n328), .A2(MEM_stage_inst_dmem_n337), .ZN(MEM_stage_inst_dmem_n7923) );
NAND2_X1 MEM_stage_inst_dmem_U483 ( .A1(MEM_stage_inst_dmem_ram_256), .A2(MEM_stage_inst_dmem_n7898), .ZN(MEM_stage_inst_dmem_n330) );
NAND2_X1 MEM_stage_inst_dmem_U482 ( .A1(MEM_stage_inst_dmem_n327), .A2(MEM_stage_inst_dmem_n326), .ZN(MEM_stage_inst_dmem_n332) );
NAND2_X1 MEM_stage_inst_dmem_U481 ( .A1(MEM_stage_inst_dmem_ram_800), .A2(MEM_stage_inst_dmem_n26), .ZN(MEM_stage_inst_dmem_n326) );
NOR2_X1 MEM_stage_inst_dmem_U480 ( .A1(MEM_stage_inst_dmem_n328), .A2(MEM_stage_inst_dmem_n325), .ZN(MEM_stage_inst_dmem_n3137) );
NAND2_X1 MEM_stage_inst_dmem_U479 ( .A1(MEM_stage_inst_dmem_ram_288), .A2(MEM_stage_inst_dmem_n67), .ZN(MEM_stage_inst_dmem_n327) );
NOR2_X1 MEM_stage_inst_dmem_U478 ( .A1(MEM_stage_inst_dmem_n348), .A2(MEM_stage_inst_dmem_n325), .ZN(MEM_stage_inst_dmem_n3209) );
NOR2_X1 MEM_stage_inst_dmem_U477 ( .A1(MEM_stage_inst_dmem_n324), .A2(MEM_stage_inst_dmem_n323), .ZN(MEM_stage_inst_dmem_n370) );
NAND2_X1 MEM_stage_inst_dmem_U476 ( .A1(MEM_stage_inst_dmem_n322), .A2(MEM_stage_inst_dmem_n321), .ZN(MEM_stage_inst_dmem_n323) );
NOR2_X1 MEM_stage_inst_dmem_U475 ( .A1(MEM_stage_inst_dmem_n320), .A2(MEM_stage_inst_dmem_n319), .ZN(MEM_stage_inst_dmem_n321) );
NAND2_X1 MEM_stage_inst_dmem_U474 ( .A1(MEM_stage_inst_dmem_n318), .A2(MEM_stage_inst_dmem_n317), .ZN(MEM_stage_inst_dmem_n319) );
NAND2_X1 MEM_stage_inst_dmem_U473 ( .A1(MEM_stage_inst_dmem_ram_496), .A2(MEM_stage_inst_dmem_n8535), .ZN(MEM_stage_inst_dmem_n317) );
BUF_X1 MEM_stage_inst_dmem_U472 ( .A(MEM_stage_inst_dmem_n3170), .Z(MEM_stage_inst_dmem_n8535) );
NOR2_X1 MEM_stage_inst_dmem_U471 ( .A1(MEM_stage_inst_dmem_n336), .A2(MEM_stage_inst_dmem_n316), .ZN(MEM_stage_inst_dmem_n3170) );
NAND2_X1 MEM_stage_inst_dmem_U470 ( .A1(MEM_stage_inst_dmem_ram_480), .A2(MEM_stage_inst_dmem_n19), .ZN(MEM_stage_inst_dmem_n318) );
NOR2_X1 MEM_stage_inst_dmem_U469 ( .A1(MEM_stage_inst_dmem_n337), .A2(MEM_stage_inst_dmem_n316), .ZN(MEM_stage_inst_dmem_n4667) );
NAND2_X1 MEM_stage_inst_dmem_U468 ( .A1(MEM_stage_inst_dmem_n315), .A2(MEM_stage_inst_dmem_n314), .ZN(MEM_stage_inst_dmem_n320) );
NAND2_X1 MEM_stage_inst_dmem_U467 ( .A1(MEM_stage_inst_dmem_ram_400), .A2(MEM_stage_inst_dmem_n23), .ZN(MEM_stage_inst_dmem_n314) );
NOR2_X1 MEM_stage_inst_dmem_U466 ( .A1(MEM_stage_inst_dmem_n316), .A2(MEM_stage_inst_dmem_n357), .ZN(MEM_stage_inst_dmem_n3160) );
NAND2_X1 MEM_stage_inst_dmem_U465 ( .A1(MEM_stage_inst_dmem_ram_816), .A2(MEM_stage_inst_dmem_n46), .ZN(MEM_stage_inst_dmem_n315) );
NOR2_X1 MEM_stage_inst_dmem_U464 ( .A1(MEM_stage_inst_dmem_n328), .A2(MEM_stage_inst_dmem_n333), .ZN(MEM_stage_inst_dmem_n4740) );
NOR2_X1 MEM_stage_inst_dmem_U463 ( .A1(MEM_stage_inst_dmem_n313), .A2(MEM_stage_inst_dmem_n312), .ZN(MEM_stage_inst_dmem_n322) );
NAND2_X1 MEM_stage_inst_dmem_U462 ( .A1(MEM_stage_inst_dmem_n311), .A2(MEM_stage_inst_dmem_n310), .ZN(MEM_stage_inst_dmem_n312) );
NAND2_X1 MEM_stage_inst_dmem_U461 ( .A1(MEM_stage_inst_dmem_ram_560), .A2(MEM_stage_inst_dmem_n41), .ZN(MEM_stage_inst_dmem_n310) );
NOR2_X1 MEM_stage_inst_dmem_U460 ( .A1(MEM_stage_inst_dmem_n333), .A2(MEM_stage_inst_dmem_n309), .ZN(MEM_stage_inst_dmem_n3085) );
NAND2_X1 MEM_stage_inst_dmem_U459 ( .A1(MEM_stage_inst_dmem_ram_672), .A2(MEM_stage_inst_dmem_n58), .ZN(MEM_stage_inst_dmem_n311) );
NOR2_X1 MEM_stage_inst_dmem_U458 ( .A1(MEM_stage_inst_dmem_n359), .A2(MEM_stage_inst_dmem_n325), .ZN(MEM_stage_inst_dmem_n3155) );
NAND2_X1 MEM_stage_inst_dmem_U457 ( .A1(MEM_stage_inst_dmem_n308), .A2(MEM_stage_inst_dmem_n307), .ZN(MEM_stage_inst_dmem_n313) );
NAND2_X1 MEM_stage_inst_dmem_U456 ( .A1(MEM_stage_inst_dmem_ram_32), .A2(MEM_stage_inst_dmem_n73), .ZN(MEM_stage_inst_dmem_n307) );
NOR2_X1 MEM_stage_inst_dmem_U455 ( .A1(MEM_stage_inst_dmem_n358), .A2(MEM_stage_inst_dmem_n325), .ZN(MEM_stage_inst_dmem_n3092) );
NAND2_X1 MEM_stage_inst_dmem_U454 ( .A1(MEM_stage_inst_dmem_ram_96), .A2(MEM_stage_inst_dmem_n56), .ZN(MEM_stage_inst_dmem_n308) );
NOR2_X1 MEM_stage_inst_dmem_U453 ( .A1(MEM_stage_inst_dmem_n337), .A2(MEM_stage_inst_dmem_n358), .ZN(MEM_stage_inst_dmem_n3179) );
NAND2_X1 MEM_stage_inst_dmem_U452 ( .A1(MEM_stage_inst_dmem_n306), .A2(MEM_stage_inst_dmem_n305), .ZN(MEM_stage_inst_dmem_n324) );
NOR2_X1 MEM_stage_inst_dmem_U451 ( .A1(MEM_stage_inst_dmem_n304), .A2(MEM_stage_inst_dmem_n303), .ZN(MEM_stage_inst_dmem_n305) );
NAND2_X1 MEM_stage_inst_dmem_U450 ( .A1(MEM_stage_inst_dmem_n302), .A2(MEM_stage_inst_dmem_n301), .ZN(MEM_stage_inst_dmem_n303) );
NAND2_X1 MEM_stage_inst_dmem_U449 ( .A1(MEM_stage_inst_dmem_ram_768), .A2(MEM_stage_inst_dmem_n8472), .ZN(MEM_stage_inst_dmem_n301) );
BUF_X1 MEM_stage_inst_dmem_U448 ( .A(MEM_stage_inst_dmem_n7992), .Z(MEM_stage_inst_dmem_n8472) );
NOR2_X1 MEM_stage_inst_dmem_U447 ( .A1(MEM_stage_inst_dmem_n328), .A2(MEM_stage_inst_dmem_n360), .ZN(MEM_stage_inst_dmem_n7992) );
NAND2_X1 MEM_stage_inst_dmem_U446 ( .A1(MEM_stage_inst_dmem_ram_304), .A2(MEM_stage_inst_dmem_n54), .ZN(MEM_stage_inst_dmem_n302) );
NOR2_X1 MEM_stage_inst_dmem_U445 ( .A1(MEM_stage_inst_dmem_n348), .A2(MEM_stage_inst_dmem_n333), .ZN(MEM_stage_inst_dmem_n4731) );
NAND2_X1 MEM_stage_inst_dmem_U444 ( .A1(MEM_stage_inst_dmem_n300), .A2(MEM_stage_inst_dmem_n299), .ZN(MEM_stage_inst_dmem_n304) );
NAND2_X1 MEM_stage_inst_dmem_U443 ( .A1(MEM_stage_inst_dmem_ram_976), .A2(MEM_stage_inst_dmem_n35), .ZN(MEM_stage_inst_dmem_n299) );
NOR2_X1 MEM_stage_inst_dmem_U442 ( .A1(MEM_stage_inst_dmem_n347), .A2(MEM_stage_inst_dmem_n344), .ZN(MEM_stage_inst_dmem_n7895) );
NAND2_X1 MEM_stage_inst_dmem_U441 ( .A1(MEM_stage_inst_dmem_ram_272), .A2(MEM_stage_inst_dmem_n62), .ZN(MEM_stage_inst_dmem_n300) );
NOR2_X1 MEM_stage_inst_dmem_U440 ( .A1(MEM_stage_inst_dmem_n348), .A2(MEM_stage_inst_dmem_n357), .ZN(MEM_stage_inst_dmem_n4672) );
NOR2_X1 MEM_stage_inst_dmem_U439 ( .A1(MEM_stage_inst_dmem_n298), .A2(MEM_stage_inst_dmem_n297), .ZN(MEM_stage_inst_dmem_n306) );
NAND2_X1 MEM_stage_inst_dmem_U438 ( .A1(MEM_stage_inst_dmem_n296), .A2(MEM_stage_inst_dmem_n295), .ZN(MEM_stage_inst_dmem_n297) );
NAND2_X1 MEM_stage_inst_dmem_U437 ( .A1(MEM_stage_inst_dmem_ram_928), .A2(MEM_stage_inst_dmem_n76), .ZN(MEM_stage_inst_dmem_n295) );
NOR2_X1 MEM_stage_inst_dmem_U436 ( .A1(MEM_stage_inst_dmem_n344), .A2(MEM_stage_inst_dmem_n325), .ZN(MEM_stage_inst_dmem_n4675) );
NAND2_X1 MEM_stage_inst_dmem_U435 ( .A1(MEM_stage_inst_dmem_ram_592), .A2(MEM_stage_inst_dmem_n53), .ZN(MEM_stage_inst_dmem_n296) );
NOR2_X1 MEM_stage_inst_dmem_U434 ( .A1(MEM_stage_inst_dmem_n347), .A2(MEM_stage_inst_dmem_n309), .ZN(MEM_stage_inst_dmem_n3140) );
NAND2_X1 MEM_stage_inst_dmem_U433 ( .A1(MEM_stage_inst_dmem_n294), .A2(MEM_stage_inst_dmem_n293), .ZN(MEM_stage_inst_dmem_n298) );
NAND2_X1 MEM_stage_inst_dmem_U432 ( .A1(MEM_stage_inst_dmem_ram_848), .A2(MEM_stage_inst_dmem_n3141), .ZN(MEM_stage_inst_dmem_n293) );
NAND2_X1 MEM_stage_inst_dmem_U431 ( .A1(MEM_stage_inst_dmem_ram_416), .A2(MEM_stage_inst_dmem_n8421), .ZN(MEM_stage_inst_dmem_n294) );
NAND2_X1 MEM_stage_inst_dmem_U430 ( .A1(MEM_stage_inst_dmem_n292), .A2(MEM_stage_inst_dmem_n291), .ZN(MEM_stage_inst_dmem_n372) );
NOR2_X1 MEM_stage_inst_dmem_U429 ( .A1(MEM_stage_inst_dmem_n290), .A2(MEM_stage_inst_dmem_n289), .ZN(MEM_stage_inst_dmem_n291) );
NAND2_X1 MEM_stage_inst_dmem_U428 ( .A1(MEM_stage_inst_dmem_n288), .A2(MEM_stage_inst_dmem_n287), .ZN(MEM_stage_inst_dmem_n289) );
NOR2_X1 MEM_stage_inst_dmem_U427 ( .A1(MEM_stage_inst_dmem_n286), .A2(MEM_stage_inst_dmem_n285), .ZN(MEM_stage_inst_dmem_n287) );
NAND2_X1 MEM_stage_inst_dmem_U426 ( .A1(MEM_stage_inst_dmem_n284), .A2(MEM_stage_inst_dmem_n283), .ZN(MEM_stage_inst_dmem_n285) );
NAND2_X1 MEM_stage_inst_dmem_U425 ( .A1(MEM_stage_inst_dmem_ram_64), .A2(MEM_stage_inst_dmem_n29), .ZN(MEM_stage_inst_dmem_n283) );
NOR2_X1 MEM_stage_inst_dmem_U424 ( .A1(MEM_stage_inst_dmem_n354), .A2(MEM_stage_inst_dmem_n358), .ZN(MEM_stage_inst_dmem_n3102) );
NAND2_X1 MEM_stage_inst_dmem_U423 ( .A1(MEM_stage_inst_dmem_ram_144), .A2(MEM_stage_inst_dmem_n44), .ZN(MEM_stage_inst_dmem_n284) );
NOR2_X1 MEM_stage_inst_dmem_U422 ( .A1(MEM_stage_inst_dmem_n353), .A2(MEM_stage_inst_dmem_n357), .ZN(MEM_stage_inst_dmem_n7903) );
NAND2_X1 MEM_stage_inst_dmem_U421 ( .A1(MEM_stage_inst_dmem_n282), .A2(MEM_stage_inst_dmem_n281), .ZN(MEM_stage_inst_dmem_n286) );
NAND2_X1 MEM_stage_inst_dmem_U420 ( .A1(MEM_stage_inst_dmem_ram_208), .A2(MEM_stage_inst_dmem_n51), .ZN(MEM_stage_inst_dmem_n281) );
NOR2_X1 MEM_stage_inst_dmem_U419 ( .A1(MEM_stage_inst_dmem_n353), .A2(MEM_stage_inst_dmem_n347), .ZN(MEM_stage_inst_dmem_n3220) );
NAND2_X1 MEM_stage_inst_dmem_U418 ( .A1(MEM_stage_inst_dmem_ram_736), .A2(MEM_stage_inst_dmem_n22), .ZN(MEM_stage_inst_dmem_n282) );
NOR2_X1 MEM_stage_inst_dmem_U417 ( .A1(MEM_stage_inst_dmem_n337), .A2(MEM_stage_inst_dmem_n359), .ZN(MEM_stage_inst_dmem_n4769) );
NOR2_X1 MEM_stage_inst_dmem_U416 ( .A1(MEM_stage_inst_dmem_n280), .A2(MEM_stage_inst_dmem_n279), .ZN(MEM_stage_inst_dmem_n288) );
NAND2_X1 MEM_stage_inst_dmem_U415 ( .A1(MEM_stage_inst_dmem_n278), .A2(MEM_stage_inst_dmem_n277), .ZN(MEM_stage_inst_dmem_n279) );
NAND2_X1 MEM_stage_inst_dmem_U414 ( .A1(MEM_stage_inst_dmem_ram_960), .A2(MEM_stage_inst_dmem_n42), .ZN(MEM_stage_inst_dmem_n277) );
NOR2_X1 MEM_stage_inst_dmem_U413 ( .A1(MEM_stage_inst_dmem_n354), .A2(MEM_stage_inst_dmem_n344), .ZN(MEM_stage_inst_dmem_n4728) );
NAND2_X1 MEM_stage_inst_dmem_U412 ( .A1(MEM_stage_inst_dmem_ram_448), .A2(MEM_stage_inst_dmem_n48), .ZN(MEM_stage_inst_dmem_n278) );
NOR2_X1 MEM_stage_inst_dmem_U411 ( .A1(MEM_stage_inst_dmem_n354), .A2(MEM_stage_inst_dmem_n316), .ZN(MEM_stage_inst_dmem_n3173) );
NAND2_X1 MEM_stage_inst_dmem_U410 ( .A1(MEM_stage_inst_dmem_n276), .A2(MEM_stage_inst_dmem_n275), .ZN(MEM_stage_inst_dmem_n280) );
NAND2_X1 MEM_stage_inst_dmem_U409 ( .A1(MEM_stage_inst_dmem_ram_944), .A2(MEM_stage_inst_dmem_n34), .ZN(MEM_stage_inst_dmem_n275) );
NOR2_X1 MEM_stage_inst_dmem_U408 ( .A1(MEM_stage_inst_dmem_n333), .A2(MEM_stage_inst_dmem_n344), .ZN(MEM_stage_inst_dmem_n3163) );
NAND2_X1 MEM_stage_inst_dmem_U407 ( .A1(MEM_stage_inst_dmem_ram_624), .A2(MEM_stage_inst_dmem_n32), .ZN(MEM_stage_inst_dmem_n276) );
NOR2_X1 MEM_stage_inst_dmem_U406 ( .A1(MEM_stage_inst_dmem_n336), .A2(MEM_stage_inst_dmem_n309), .ZN(MEM_stage_inst_dmem_n4652) );
NAND2_X1 MEM_stage_inst_dmem_U405 ( .A1(MEM_stage_inst_dmem_n274), .A2(MEM_stage_inst_dmem_n273), .ZN(MEM_stage_inst_dmem_n290) );
NOR2_X1 MEM_stage_inst_dmem_U404 ( .A1(MEM_stage_inst_dmem_n272), .A2(MEM_stage_inst_dmem_n271), .ZN(MEM_stage_inst_dmem_n273) );
NAND2_X1 MEM_stage_inst_dmem_U403 ( .A1(MEM_stage_inst_dmem_n270), .A2(MEM_stage_inst_dmem_n269), .ZN(MEM_stage_inst_dmem_n271) );
NAND2_X1 MEM_stage_inst_dmem_U402 ( .A1(MEM_stage_inst_dmem_ram_896), .A2(MEM_stage_inst_dmem_n72), .ZN(MEM_stage_inst_dmem_n269) );
NOR2_X1 MEM_stage_inst_dmem_U401 ( .A1(MEM_stage_inst_dmem_n360), .A2(MEM_stage_inst_dmem_n344), .ZN(MEM_stage_inst_dmem_n3123) );
NAND2_X1 MEM_stage_inst_dmem_U400 ( .A1(MEM_stage_inst_dmem_ram_0), .A2(MEM_stage_inst_dmem_n77), .ZN(MEM_stage_inst_dmem_n270) );
NOR2_X1 MEM_stage_inst_dmem_U399 ( .A1(MEM_stage_inst_dmem_n360), .A2(MEM_stage_inst_dmem_n358), .ZN(MEM_stage_inst_dmem_n7953) );
NAND2_X1 MEM_stage_inst_dmem_U398 ( .A1(MEM_stage_inst_dmem_n268), .A2(MEM_stage_inst_dmem_n267), .ZN(MEM_stage_inst_dmem_n272) );
NAND2_X1 MEM_stage_inst_dmem_U397 ( .A1(MEM_stage_inst_dmem_ram_880), .A2(MEM_stage_inst_dmem_n21), .ZN(MEM_stage_inst_dmem_n267) );
NOR2_X1 MEM_stage_inst_dmem_U396 ( .A1(MEM_stage_inst_dmem_n336), .A2(MEM_stage_inst_dmem_n328), .ZN(MEM_stage_inst_dmem_n3099) );
NAND2_X1 MEM_stage_inst_dmem_U395 ( .A1(MEM_stage_inst_dmem_ram_464), .A2(MEM_stage_inst_dmem_n65), .ZN(MEM_stage_inst_dmem_n268) );
NOR2_X1 MEM_stage_inst_dmem_U394 ( .A1(MEM_stage_inst_dmem_n316), .A2(MEM_stage_inst_dmem_n347), .ZN(MEM_stage_inst_dmem_n3174) );
NOR2_X1 MEM_stage_inst_dmem_U393 ( .A1(MEM_stage_inst_dmem_n266), .A2(MEM_stage_inst_dmem_n265), .ZN(MEM_stage_inst_dmem_n274) );
NAND2_X1 MEM_stage_inst_dmem_U392 ( .A1(MEM_stage_inst_dmem_n264), .A2(MEM_stage_inst_dmem_n263), .ZN(MEM_stage_inst_dmem_n265) );
NAND2_X1 MEM_stage_inst_dmem_U391 ( .A1(MEM_stage_inst_dmem_ram_432), .A2(MEM_stage_inst_dmem_n43), .ZN(MEM_stage_inst_dmem_n263) );
NOR2_X1 MEM_stage_inst_dmem_U390 ( .A1(MEM_stage_inst_dmem_n316), .A2(MEM_stage_inst_dmem_n333), .ZN(MEM_stage_inst_dmem_n7888) );
NAND2_X1 MEM_stage_inst_dmem_U389 ( .A1(MEM_stage_inst_dmem_ram_240), .A2(MEM_stage_inst_dmem_n39), .ZN(MEM_stage_inst_dmem_n264) );
NOR2_X1 MEM_stage_inst_dmem_U388 ( .A1(MEM_stage_inst_dmem_n336), .A2(MEM_stage_inst_dmem_n353), .ZN(MEM_stage_inst_dmem_n4649) );
NAND2_X1 MEM_stage_inst_dmem_U387 ( .A1(MEM_stage_inst_dmem_n262), .A2(MEM_stage_inst_dmem_n261), .ZN(MEM_stage_inst_dmem_n266) );
NAND2_X1 MEM_stage_inst_dmem_U386 ( .A1(MEM_stage_inst_dmem_ram_832), .A2(MEM_stage_inst_dmem_n57), .ZN(MEM_stage_inst_dmem_n261) );
NOR2_X1 MEM_stage_inst_dmem_U385 ( .A1(MEM_stage_inst_dmem_n328), .A2(MEM_stage_inst_dmem_n354), .ZN(MEM_stage_inst_dmem_n3120) );
NAND2_X1 MEM_stage_inst_dmem_U384 ( .A1(MEM_stage_inst_dmem_ram_1008), .A2(MEM_stage_inst_dmem_n60), .ZN(MEM_stage_inst_dmem_n262) );
NOR2_X1 MEM_stage_inst_dmem_U383 ( .A1(MEM_stage_inst_dmem_n336), .A2(MEM_stage_inst_dmem_n344), .ZN(MEM_stage_inst_dmem_n3199) );
NAND2_X1 MEM_stage_inst_dmem_U382 ( .A1(MEM_stage_inst_dmem_n260), .A2(MEM_stage_inst_dmem_n15966), .ZN(MEM_stage_inst_dmem_n344) );
NOR2_X1 MEM_stage_inst_dmem_U381 ( .A1(MEM_stage_inst_dmem_n259), .A2(MEM_stage_inst_dmem_n258), .ZN(MEM_stage_inst_dmem_n292) );
NAND2_X1 MEM_stage_inst_dmem_U380 ( .A1(MEM_stage_inst_dmem_n257), .A2(MEM_stage_inst_dmem_n256), .ZN(MEM_stage_inst_dmem_n258) );
NOR2_X1 MEM_stage_inst_dmem_U379 ( .A1(MEM_stage_inst_dmem_n255), .A2(MEM_stage_inst_dmem_n254), .ZN(MEM_stage_inst_dmem_n256) );
NAND2_X1 MEM_stage_inst_dmem_U378 ( .A1(MEM_stage_inst_dmem_n253), .A2(MEM_stage_inst_dmem_n252), .ZN(MEM_stage_inst_dmem_n254) );
NAND2_X1 MEM_stage_inst_dmem_U377 ( .A1(MEM_stage_inst_dmem_ram_48), .A2(MEM_stage_inst_dmem_n68), .ZN(MEM_stage_inst_dmem_n252) );
NOR2_X1 MEM_stage_inst_dmem_U376 ( .A1(MEM_stage_inst_dmem_n333), .A2(MEM_stage_inst_dmem_n358), .ZN(MEM_stage_inst_dmem_n3103) );
NAND2_X1 MEM_stage_inst_dmem_U375 ( .A1(MEM_stage_inst_dmem_ram_512), .A2(MEM_stage_inst_dmem_n71), .ZN(MEM_stage_inst_dmem_n253) );
NOR2_X1 MEM_stage_inst_dmem_U374 ( .A1(MEM_stage_inst_dmem_n360), .A2(MEM_stage_inst_dmem_n309), .ZN(MEM_stage_inst_dmem_n3182) );
NAND2_X1 MEM_stage_inst_dmem_U373 ( .A1(MEM_stage_inst_dmem_n251), .A2(MEM_stage_inst_dmem_n250), .ZN(MEM_stage_inst_dmem_n255) );
NAND2_X1 MEM_stage_inst_dmem_U372 ( .A1(MEM_stage_inst_dmem_ram_224), .A2(MEM_stage_inst_dmem_n28), .ZN(MEM_stage_inst_dmem_n250) );
NOR2_X1 MEM_stage_inst_dmem_U371 ( .A1(MEM_stage_inst_dmem_n353), .A2(MEM_stage_inst_dmem_n337), .ZN(MEM_stage_inst_dmem_n3152) );
NAND2_X1 MEM_stage_inst_dmem_U370 ( .A1(MEM_stage_inst_dmem_ram_528), .A2(MEM_stage_inst_dmem_n45), .ZN(MEM_stage_inst_dmem_n251) );
NOR2_X1 MEM_stage_inst_dmem_U369 ( .A1(MEM_stage_inst_dmem_n309), .A2(MEM_stage_inst_dmem_n357), .ZN(MEM_stage_inst_dmem_n7884) );
NOR2_X1 MEM_stage_inst_dmem_U368 ( .A1(MEM_stage_inst_dmem_n249), .A2(MEM_stage_inst_dmem_n248), .ZN(MEM_stage_inst_dmem_n257) );
NAND2_X1 MEM_stage_inst_dmem_U367 ( .A1(MEM_stage_inst_dmem_n247), .A2(MEM_stage_inst_dmem_n246), .ZN(MEM_stage_inst_dmem_n248) );
NAND2_X1 MEM_stage_inst_dmem_U366 ( .A1(MEM_stage_inst_dmem_ram_752), .A2(MEM_stage_inst_dmem_n20), .ZN(MEM_stage_inst_dmem_n246) );
NOR2_X1 MEM_stage_inst_dmem_U365 ( .A1(MEM_stage_inst_dmem_n336), .A2(MEM_stage_inst_dmem_n359), .ZN(MEM_stage_inst_dmem_n3202) );
NAND2_X1 MEM_stage_inst_dmem_U364 ( .A1(MEM_stage_inst_dmem_ram_656), .A2(MEM_stage_inst_dmem_n8325), .ZN(MEM_stage_inst_dmem_n247) );
NAND2_X1 MEM_stage_inst_dmem_U363 ( .A1(MEM_stage_inst_dmem_n245), .A2(MEM_stage_inst_dmem_n244), .ZN(MEM_stage_inst_dmem_n249) );
NAND2_X1 MEM_stage_inst_dmem_U362 ( .A1(MEM_stage_inst_dmem_ram_384), .A2(MEM_stage_inst_dmem_n75), .ZN(MEM_stage_inst_dmem_n244) );
NOR2_X1 MEM_stage_inst_dmem_U361 ( .A1(MEM_stage_inst_dmem_n360), .A2(MEM_stage_inst_dmem_n316), .ZN(MEM_stage_inst_dmem_n7930) );
NAND2_X1 MEM_stage_inst_dmem_U360 ( .A1(EX_pipeline_reg_out_27), .A2(MEM_stage_inst_dmem_n260), .ZN(MEM_stage_inst_dmem_n316) );
AND2_X1 MEM_stage_inst_dmem_U359 ( .A1(EX_pipeline_reg_out_26), .A2(EX_pipeline_reg_out_25), .ZN(MEM_stage_inst_dmem_n260) );
NAND2_X1 MEM_stage_inst_dmem_U358 ( .A1(MEM_stage_inst_dmem_n243), .A2(MEM_stage_inst_dmem_n8761), .ZN(MEM_stage_inst_dmem_n360) );
NAND2_X1 MEM_stage_inst_dmem_U357 ( .A1(MEM_stage_inst_dmem_ram_160), .A2(MEM_stage_inst_dmem_n69), .ZN(MEM_stage_inst_dmem_n245) );
NOR2_X1 MEM_stage_inst_dmem_U356 ( .A1(MEM_stage_inst_dmem_n353), .A2(MEM_stage_inst_dmem_n325), .ZN(MEM_stage_inst_dmem_n3081) );
NAND2_X1 MEM_stage_inst_dmem_U355 ( .A1(EX_pipeline_reg_out_27), .A2(MEM_stage_inst_dmem_n242), .ZN(MEM_stage_inst_dmem_n353) );
NAND2_X1 MEM_stage_inst_dmem_U354 ( .A1(MEM_stage_inst_dmem_n241), .A2(MEM_stage_inst_dmem_n240), .ZN(MEM_stage_inst_dmem_n259) );
NOR2_X1 MEM_stage_inst_dmem_U353 ( .A1(MEM_stage_inst_dmem_n239), .A2(MEM_stage_inst_dmem_n238), .ZN(MEM_stage_inst_dmem_n240) );
NAND2_X1 MEM_stage_inst_dmem_U352 ( .A1(MEM_stage_inst_dmem_n237), .A2(MEM_stage_inst_dmem_n236), .ZN(MEM_stage_inst_dmem_n238) );
NAND2_X1 MEM_stage_inst_dmem_U351 ( .A1(MEM_stage_inst_dmem_ram_688), .A2(MEM_stage_inst_dmem_n50), .ZN(MEM_stage_inst_dmem_n236) );
NOR2_X1 MEM_stage_inst_dmem_U350 ( .A1(MEM_stage_inst_dmem_n333), .A2(MEM_stage_inst_dmem_n359), .ZN(MEM_stage_inst_dmem_n4709) );
NAND2_X1 MEM_stage_inst_dmem_U349 ( .A1(EX_pipeline_reg_out_23), .A2(MEM_stage_inst_dmem_n235), .ZN(MEM_stage_inst_dmem_n333) );
NAND2_X1 MEM_stage_inst_dmem_U348 ( .A1(MEM_stage_inst_dmem_ram_80), .A2(MEM_stage_inst_dmem_n40), .ZN(MEM_stage_inst_dmem_n237) );
NOR2_X1 MEM_stage_inst_dmem_U347 ( .A1(MEM_stage_inst_dmem_n347), .A2(MEM_stage_inst_dmem_n358), .ZN(MEM_stage_inst_dmem_n7938) );
NAND2_X1 MEM_stage_inst_dmem_U346 ( .A1(EX_pipeline_reg_out_27), .A2(MEM_stage_inst_dmem_n234), .ZN(MEM_stage_inst_dmem_n358) );
NAND2_X1 MEM_stage_inst_dmem_U345 ( .A1(MEM_stage_inst_dmem_n233), .A2(MEM_stage_inst_dmem_n232), .ZN(MEM_stage_inst_dmem_n239) );
NAND2_X1 MEM_stage_inst_dmem_U344 ( .A1(MEM_stage_inst_dmem_ram_608), .A2(MEM_stage_inst_dmem_n30), .ZN(MEM_stage_inst_dmem_n232) );
NOR2_X1 MEM_stage_inst_dmem_U343 ( .A1(MEM_stage_inst_dmem_n337), .A2(MEM_stage_inst_dmem_n309), .ZN(MEM_stage_inst_dmem_n4701) );
NAND2_X1 MEM_stage_inst_dmem_U342 ( .A1(EX_pipeline_reg_out_23), .A2(MEM_stage_inst_dmem_n231), .ZN(MEM_stage_inst_dmem_n337) );
NAND2_X1 MEM_stage_inst_dmem_U341 ( .A1(MEM_stage_inst_dmem_ram_784), .A2(MEM_stage_inst_dmem_n38), .ZN(MEM_stage_inst_dmem_n233) );
NOR2_X1 MEM_stage_inst_dmem_U340 ( .A1(MEM_stage_inst_dmem_n328), .A2(MEM_stage_inst_dmem_n357), .ZN(MEM_stage_inst_dmem_n3191) );
NAND2_X1 MEM_stage_inst_dmem_U339 ( .A1(MEM_stage_inst_dmem_n235), .A2(MEM_stage_inst_dmem_n8761), .ZN(MEM_stage_inst_dmem_n357) );
NOR2_X1 MEM_stage_inst_dmem_U338 ( .A1(EX_pipeline_reg_out_24), .A2(MEM_stage_inst_dmem_n12963), .ZN(MEM_stage_inst_dmem_n235) );
NAND2_X1 MEM_stage_inst_dmem_U337 ( .A1(MEM_stage_inst_dmem_n230), .A2(MEM_stage_inst_dmem_n15966), .ZN(MEM_stage_inst_dmem_n328) );
NOR2_X1 MEM_stage_inst_dmem_U336 ( .A1(MEM_stage_inst_dmem_n229), .A2(MEM_stage_inst_dmem_n228), .ZN(MEM_stage_inst_dmem_n241) );
NAND2_X1 MEM_stage_inst_dmem_U335 ( .A1(MEM_stage_inst_dmem_n227), .A2(MEM_stage_inst_dmem_n226), .ZN(MEM_stage_inst_dmem_n228) );
NAND2_X1 MEM_stage_inst_dmem_U334 ( .A1(MEM_stage_inst_dmem_ram_544), .A2(MEM_stage_inst_dmem_n74), .ZN(MEM_stage_inst_dmem_n226) );
NOR2_X1 MEM_stage_inst_dmem_U333 ( .A1(MEM_stage_inst_dmem_n309), .A2(MEM_stage_inst_dmem_n325), .ZN(MEM_stage_inst_dmem_n4692) );
NAND2_X1 MEM_stage_inst_dmem_U332 ( .A1(EX_pipeline_reg_out_23), .A2(MEM_stage_inst_dmem_n243), .ZN(MEM_stage_inst_dmem_n325) );
NOR2_X1 MEM_stage_inst_dmem_U331 ( .A1(EX_pipeline_reg_out_22), .A2(EX_pipeline_reg_out_24), .ZN(MEM_stage_inst_dmem_n243) );
NAND2_X1 MEM_stage_inst_dmem_U330 ( .A1(MEM_stage_inst_dmem_ram_576), .A2(MEM_stage_inst_dmem_n27), .ZN(MEM_stage_inst_dmem_n227) );
NOR2_X1 MEM_stage_inst_dmem_U329 ( .A1(MEM_stage_inst_dmem_n354), .A2(MEM_stage_inst_dmem_n309), .ZN(MEM_stage_inst_dmem_n7973) );
NAND2_X1 MEM_stage_inst_dmem_U328 ( .A1(MEM_stage_inst_dmem_n234), .A2(MEM_stage_inst_dmem_n15966), .ZN(MEM_stage_inst_dmem_n309) );
NOR2_X1 MEM_stage_inst_dmem_U327 ( .A1(EX_pipeline_reg_out_26), .A2(EX_pipeline_reg_out_25), .ZN(MEM_stage_inst_dmem_n234) );
NAND2_X1 MEM_stage_inst_dmem_U326 ( .A1(MEM_stage_inst_dmem_n231), .A2(MEM_stage_inst_dmem_n8761), .ZN(MEM_stage_inst_dmem_n354) );
NOR2_X1 MEM_stage_inst_dmem_U325 ( .A1(EX_pipeline_reg_out_22), .A2(MEM_stage_inst_dmem_n8762), .ZN(MEM_stage_inst_dmem_n231) );
NAND2_X1 MEM_stage_inst_dmem_U324 ( .A1(MEM_stage_inst_dmem_n225), .A2(MEM_stage_inst_dmem_n224), .ZN(MEM_stage_inst_dmem_n229) );
NAND2_X1 MEM_stage_inst_dmem_U323 ( .A1(MEM_stage_inst_dmem_ram_720), .A2(MEM_stage_inst_dmem_n31), .ZN(MEM_stage_inst_dmem_n224) );
NOR2_X1 MEM_stage_inst_dmem_U322 ( .A1(MEM_stage_inst_dmem_n347), .A2(MEM_stage_inst_dmem_n359), .ZN(MEM_stage_inst_dmem_n3112) );
NAND2_X1 MEM_stage_inst_dmem_U321 ( .A1(MEM_stage_inst_dmem_n242), .A2(MEM_stage_inst_dmem_n15966), .ZN(MEM_stage_inst_dmem_n359) );
INV_X1 MEM_stage_inst_dmem_U320 ( .A(EX_pipeline_reg_out_27), .ZN(MEM_stage_inst_dmem_n15966) );
NOR2_X1 MEM_stage_inst_dmem_U319 ( .A1(EX_pipeline_reg_out_26), .A2(MEM_stage_inst_dmem_n12964), .ZN(MEM_stage_inst_dmem_n242) );
NAND2_X1 MEM_stage_inst_dmem_U318 ( .A1(MEM_stage_inst_dmem_n223), .A2(MEM_stage_inst_dmem_n8761), .ZN(MEM_stage_inst_dmem_n347) );
INV_X1 MEM_stage_inst_dmem_U317 ( .A(EX_pipeline_reg_out_23), .ZN(MEM_stage_inst_dmem_n8761) );
NAND2_X1 MEM_stage_inst_dmem_U316 ( .A1(MEM_stage_inst_dmem_ram_368), .A2(MEM_stage_inst_dmem_n33), .ZN(MEM_stage_inst_dmem_n225) );
NOR2_X1 MEM_stage_inst_dmem_U315 ( .A1(MEM_stage_inst_dmem_n336), .A2(MEM_stage_inst_dmem_n348), .ZN(MEM_stage_inst_dmem_n4721) );
AND2_X1 MEM_stage_inst_dmem_U314 ( .A1(MEM_stage_inst_dmem_n12964), .A2(EX_pipeline_reg_out_26), .ZN(MEM_stage_inst_dmem_n230) );
INV_X1 MEM_stage_inst_dmem_U313 ( .A(EX_pipeline_reg_out_25), .ZN(MEM_stage_inst_dmem_n12964) );
NAND2_X1 MEM_stage_inst_dmem_U312 ( .A1(MEM_stage_inst_dmem_n223), .A2(EX_pipeline_reg_out_23), .ZN(MEM_stage_inst_dmem_n336) );
NOR2_X1 MEM_stage_inst_dmem_U311 ( .A1(MEM_stage_inst_dmem_n12963), .A2(MEM_stage_inst_dmem_n8762), .ZN(MEM_stage_inst_dmem_n223) );
INV_X1 MEM_stage_inst_dmem_U310 ( .A(EX_pipeline_reg_out_24), .ZN(MEM_stage_inst_dmem_n8762) );
INV_X1 MEM_stage_inst_dmem_U309 ( .A(EX_pipeline_reg_out_22), .ZN(MEM_stage_inst_dmem_n12963) );
INV_X1 MEM_stage_inst_dmem_U308 ( .A(MEM_stage_inst_dmem_n8655), .ZN(MEM_stage_inst_dmem_n8656) );
INV_X1 MEM_stage_inst_dmem_U307 ( .A(MEM_stage_inst_dmem_n12996), .ZN(MEM_stage_inst_dmem_n12997) );
INV_X1 MEM_stage_inst_dmem_U306 ( .A(MEM_stage_inst_dmem_n13106), .ZN(MEM_stage_inst_dmem_n13107) );
INV_X1 MEM_stage_inst_dmem_U305 ( .A(MEM_stage_inst_dmem_n13176), .ZN(MEM_stage_inst_dmem_n13177) );
INV_X1 MEM_stage_inst_dmem_U304 ( .A(MEM_stage_inst_dmem_n13418), .ZN(MEM_stage_inst_dmem_n13419) );
INV_X1 MEM_stage_inst_dmem_U303 ( .A(MEM_stage_inst_dmem_n13690), .ZN(MEM_stage_inst_dmem_n13691) );
INV_X1 MEM_stage_inst_dmem_U302 ( .A(MEM_stage_inst_dmem_n13940), .ZN(MEM_stage_inst_dmem_n13941) );
INV_X1 MEM_stage_inst_dmem_U301 ( .A(MEM_stage_inst_dmem_n14212), .ZN(MEM_stage_inst_dmem_n14213) );
INV_X1 MEM_stage_inst_dmem_U300 ( .A(MEM_stage_inst_dmem_n14451), .ZN(MEM_stage_inst_dmem_n14452) );
INV_X1 MEM_stage_inst_dmem_U299 ( .A(MEM_stage_inst_dmem_n14689), .ZN(MEM_stage_inst_dmem_n14690) );
INV_X1 MEM_stage_inst_dmem_U298 ( .A(MEM_stage_inst_dmem_n14936), .ZN(MEM_stage_inst_dmem_n14937) );
INV_X1 MEM_stage_inst_dmem_U297 ( .A(MEM_stage_inst_dmem_n15451), .ZN(MEM_stage_inst_dmem_n15452) );
INV_X1 MEM_stage_inst_dmem_U296 ( .A(MEM_stage_inst_dmem_n15587), .ZN(MEM_stage_inst_dmem_n15588) );
INV_X1 MEM_stage_inst_dmem_U295 ( .A(MEM_stage_inst_dmem_n15893), .ZN(MEM_stage_inst_dmem_n15894) );
BUF_X1 MEM_stage_inst_dmem_U294 ( .A(MEM_stage_inst_dmem_n20530), .Z(MEM_stage_inst_dmem_n16361) );
INV_X1 MEM_stage_inst_dmem_U293 ( .A(MEM_stage_inst_dmem_n16339), .ZN(MEM_stage_inst_dmem_n16340) );
INV_X1 MEM_stage_inst_dmem_U292 ( .A(MEM_stage_inst_dmem_n16618), .ZN(MEM_stage_inst_dmem_n16619) );
INV_X1 MEM_stage_inst_dmem_U291 ( .A(MEM_stage_inst_dmem_n16829), .ZN(MEM_stage_inst_dmem_n16830) );
INV_X1 MEM_stage_inst_dmem_U290 ( .A(MEM_stage_inst_dmem_n16863), .ZN(MEM_stage_inst_dmem_n16864) );
INV_X1 MEM_stage_inst_dmem_U289 ( .A(MEM_stage_inst_dmem_n17102), .ZN(MEM_stage_inst_dmem_n17103) );
INV_X1 MEM_stage_inst_dmem_U288 ( .A(MEM_stage_inst_dmem_n17374), .ZN(MEM_stage_inst_dmem_n17375) );
INV_X1 MEM_stage_inst_dmem_U287 ( .A(MEM_stage_inst_dmem_n17613), .ZN(MEM_stage_inst_dmem_n17614) );
INV_X1 MEM_stage_inst_dmem_U286 ( .A(MEM_stage_inst_dmem_n17888), .ZN(MEM_stage_inst_dmem_n17889) );
INV_X1 MEM_stage_inst_dmem_U285 ( .A(MEM_stage_inst_dmem_n18373), .ZN(MEM_stage_inst_dmem_n18374) );
INV_X1 MEM_stage_inst_dmem_U284 ( .A(MEM_stage_inst_dmem_n18611), .ZN(MEM_stage_inst_dmem_n18612) );
INV_X1 MEM_stage_inst_dmem_U283 ( .A(MEM_stage_inst_dmem_n18851), .ZN(MEM_stage_inst_dmem_n18852) );
INV_X1 MEM_stage_inst_dmem_U282 ( .A(MEM_stage_inst_dmem_n19130), .ZN(MEM_stage_inst_dmem_n19131) );
BUF_X1 MEM_stage_inst_dmem_U281 ( .A(MEM_stage_inst_dmem_n20515), .Z(MEM_stage_inst_dmem_n21474) );
INV_X1 MEM_stage_inst_dmem_U280 ( .A(MEM_stage_inst_dmem_n19580), .ZN(MEM_stage_inst_dmem_n19581) );
INV_X1 MEM_stage_inst_dmem_U279 ( .A(MEM_stage_inst_dmem_n19854), .ZN(MEM_stage_inst_dmem_n19855) );
INV_X1 MEM_stage_inst_dmem_U278 ( .A(MEM_stage_inst_dmem_n20092), .ZN(MEM_stage_inst_dmem_n20093) );
INV_X1 MEM_stage_inst_dmem_U277 ( .A(MEM_stage_inst_dmem_n20365), .ZN(MEM_stage_inst_dmem_n20366) );
BUF_X1 MEM_stage_inst_dmem_U276 ( .A(MEM_stage_inst_dmem_n20518), .Z(MEM_stage_inst_dmem_n20904) );
INV_X1 MEM_stage_inst_dmem_U275 ( .A(MEM_stage_inst_dmem_n20619), .ZN(MEM_stage_inst_dmem_n20620) );
INV_X1 MEM_stage_inst_dmem_U274 ( .A(MEM_stage_inst_dmem_n20857), .ZN(MEM_stage_inst_dmem_n20858) );
INV_X1 MEM_stage_inst_dmem_U273 ( .A(MEM_stage_inst_dmem_n21140), .ZN(MEM_stage_inst_dmem_n21141) );
INV_X1 MEM_stage_inst_dmem_U272 ( .A(MEM_stage_inst_dmem_n21390), .ZN(MEM_stage_inst_dmem_n21391) );
INV_X1 MEM_stage_inst_dmem_U271 ( .A(MEM_stage_inst_dmem_n21499), .ZN(MEM_stage_inst_dmem_n21500) );
BUF_X1 MEM_stage_inst_dmem_U270 ( .A(MEM_stage_inst_dmem_n15110), .Z(MEM_stage_inst_dmem_n16758) );
BUF_X1 MEM_stage_inst_dmem_U269 ( .A(MEM_stage_inst_dmem_n14693), .Z(MEM_stage_inst_dmem_n21320) );
BUF_X1 MEM_stage_inst_dmem_U268 ( .A(MEM_stage_inst_dmem_n14705), .Z(MEM_stage_inst_dmem_n18864) );
BUF_X1 MEM_stage_inst_dmem_U267 ( .A(MEM_stage_inst_dmem_n20512), .Z(MEM_stage_inst_dmem_n19242) );
BUF_X1 MEM_stage_inst_dmem_U266 ( .A(MEM_stage_inst_dmem_n20512), .Z(MEM_stage_inst_dmem_n15116) );
BUF_X1 MEM_stage_inst_dmem_U264 ( .A(MEM_stage_inst_dmem_n14702), .Z(MEM_stage_inst_dmem_n18861) );
BUF_X1 MEM_stage_inst_dmem_U262 ( .A(MEM_stage_inst_dmem_n20509), .Z(MEM_stage_inst_dmem_n15113) );
BUF_X1 MEM_stage_inst_dmem_U261 ( .A(MEM_stage_inst_dmem_n20509), .Z(MEM_stage_inst_dmem_n14696) );
BUF_X1 MEM_stage_inst_dmem_U260 ( .A(MEM_stage_inst_dmem_n20533), .Z(MEM_stage_inst_dmem_n14717) );
BUF_X1 MEM_stage_inst_dmem_U259 ( .A(MEM_stage_inst_dmem_n20551), .Z(MEM_stage_inst_dmem_n19275) );
BUF_X1 MEM_stage_inst_dmem_U258 ( .A(MEM_stage_inst_dmem_n20551), .Z(MEM_stage_inst_dmem_n15145) );
BUF_X1 MEM_stage_inst_dmem_U257 ( .A(MEM_stage_inst_dmem_n20551), .Z(MEM_stage_inst_dmem_n14732) );
BUF_X1 MEM_stage_inst_dmem_U256 ( .A(MEM_stage_inst_dmem_n6), .Z(MEM_stage_inst_dmem_n16784) );
BUF_X1 MEM_stage_inst_dmem_U255 ( .A(MEM_stage_inst_dmem_n6), .Z(MEM_stage_inst_dmem_n16368) );
BUF_X2 MEM_stage_inst_dmem_U254 ( .A(MEM_stage_inst_dmem_n4772), .Z(MEM_stage_inst_dmem_n8421) );
BUF_X2 MEM_stage_inst_dmem_U253 ( .A(MEM_stage_inst_dmem_n7898), .Z(MEM_stage_inst_dmem_n5857) );
BUF_X2 MEM_stage_inst_dmem_U252 ( .A(MEM_stage_inst_dmem_n3076), .Z(MEM_stage_inst_dmem_n8325) );
NOR2_X2 MEM_stage_inst_dmem_U251 ( .A1(MEM_stage_inst_dmem_n348), .A2(MEM_stage_inst_dmem_n347), .ZN(MEM_stage_inst_dmem_n3216) );
BUF_X2 MEM_stage_inst_dmem_U250 ( .A(MEM_stage_inst_dmem_n3141), .Z(MEM_stage_inst_dmem_n8372) );
NOR2_X2 MEM_stage_inst_dmem_U249 ( .A1(MEM_stage_inst_dmem_n316), .A2(MEM_stage_inst_dmem_n325), .ZN(MEM_stage_inst_dmem_n4772) );
NOR2_X2 MEM_stage_inst_dmem_U248 ( .A1(MEM_stage_inst_dmem_n328), .A2(MEM_stage_inst_dmem_n347), .ZN(MEM_stage_inst_dmem_n3141) );
NOR2_X2 MEM_stage_inst_dmem_U247 ( .A1(MEM_stage_inst_dmem_n357), .A2(MEM_stage_inst_dmem_n359), .ZN(MEM_stage_inst_dmem_n3076) );
NOR2_X2 MEM_stage_inst_dmem_U246 ( .A1(MEM_stage_inst_dmem_n360), .A2(MEM_stage_inst_dmem_n348), .ZN(MEM_stage_inst_dmem_n7898) );
NAND2_X1 MEM_stage_inst_dmem_U245 ( .A1(EX_pipeline_reg_out_27), .A2(MEM_stage_inst_dmem_n230), .ZN(MEM_stage_inst_dmem_n348) );
BUF_X2 MEM_stage_inst_dmem_U139 ( .A(EX_pipeline_reg_out_14), .Z(MEM_stage_inst_dmem_n13880) );
BUF_X2 MEM_stage_inst_dmem_U138 ( .A(EX_pipeline_reg_out_15), .Z(MEM_stage_inst_dmem_n13877) );
BUF_X2 MEM_stage_inst_dmem_U137 ( .A(MEM_stage_inst_dmem_n20506), .Z(MEM_stage_inst_dmem_n114) );
BUF_X2 MEM_stage_inst_dmem_U135 ( .A(EX_pipeline_reg_out_7), .Z(MEM_stage_inst_dmem_n13900) );
BUF_X2 MEM_stage_inst_dmem_U134 ( .A(EX_pipeline_reg_out_8), .Z(MEM_stage_inst_dmem_n13897) );
BUF_X2 MEM_stage_inst_dmem_U133 ( .A(MEM_stage_inst_dmem_n20544), .Z(MEM_stage_inst_dmem_n113) );
BUF_X2 MEM_stage_inst_dmem_U132 ( .A(EX_pipeline_reg_out_10), .Z(MEM_stage_inst_dmem_n13892) );
BUF_X2 MEM_stage_inst_dmem_U131 ( .A(EX_pipeline_reg_out_11), .Z(MEM_stage_inst_dmem_n13889) );
BUF_X2 MEM_stage_inst_dmem_U130 ( .A(EX_pipeline_reg_out_20), .Z(MEM_stage_inst_dmem_n17994) );
BUF_X2 MEM_stage_inst_dmem_U129 ( .A(EX_pipeline_reg_out_16), .Z(MEM_stage_inst_dmem_n13874) );
BUF_X2 MEM_stage_inst_dmem_U128 ( .A(EX_pipeline_reg_out_17), .Z(MEM_stage_inst_dmem_n13871) );
BUF_X2 MEM_stage_inst_dmem_U127 ( .A(MEM_stage_inst_dmem_n20515), .Z(MEM_stage_inst_dmem_n105) );
BUF_X2 MEM_stage_inst_dmem_U126 ( .A(MEM_stage_inst_dmem_n20527), .Z(MEM_stage_inst_dmem_n104) );
BUF_X2 MEM_stage_inst_dmem_U125 ( .A(MEM_stage_inst_dmem_n20518), .Z(MEM_stage_inst_dmem_n103) );
BUF_X2 MEM_stage_inst_dmem_U124 ( .A(MEM_stage_inst_dmem_n20521), .Z(MEM_stage_inst_dmem_n102) );
BUF_X2 MEM_stage_inst_dmem_U123 ( .A(MEM_stage_inst_dmem_n20530), .Z(MEM_stage_inst_dmem_n101) );
BUF_X2 MEM_stage_inst_dmem_U122 ( .A(MEM_stage_inst_dmem_n20524), .Z(MEM_stage_inst_dmem_n100) );
BUF_X2 MEM_stage_inst_dmem_U118 ( .A(MEM_stage_inst_dmem_n20521), .Z(MEM_stage_inst_dmem_n16354) );
BUF_X2 MEM_stage_inst_dmem_U116 ( .A(MEM_stage_inst_dmem_n20544), .Z(MEM_stage_inst_dmem_n16373) );
BUF_X4 MEM_stage_inst_dmem_U96 ( .A(MEM_stage_inst_dmem_n7953), .Z(MEM_stage_inst_dmem_n77) );
BUF_X4 MEM_stage_inst_dmem_U95 ( .A(MEM_stage_inst_dmem_n4675), .Z(MEM_stage_inst_dmem_n76) );
BUF_X4 MEM_stage_inst_dmem_U94 ( .A(MEM_stage_inst_dmem_n7930), .Z(MEM_stage_inst_dmem_n75) );
BUF_X4 MEM_stage_inst_dmem_U93 ( .A(MEM_stage_inst_dmem_n4692), .Z(MEM_stage_inst_dmem_n74) );
BUF_X4 MEM_stage_inst_dmem_U92 ( .A(MEM_stage_inst_dmem_n3092), .Z(MEM_stage_inst_dmem_n73) );
BUF_X2 MEM_stage_inst_dmem_U91 ( .A(MEM_stage_inst_dmem_n3123), .Z(MEM_stage_inst_dmem_n72) );
BUF_X2 MEM_stage_inst_dmem_U90 ( .A(MEM_stage_inst_dmem_n3182), .Z(MEM_stage_inst_dmem_n71) );
BUF_X4 MEM_stage_inst_dmem_U89 ( .A(MEM_stage_inst_dmem_n7887), .Z(MEM_stage_inst_dmem_n70) );
BUF_X4 MEM_stage_inst_dmem_U88 ( .A(MEM_stage_inst_dmem_n3081), .Z(MEM_stage_inst_dmem_n69) );
BUF_X4 MEM_stage_inst_dmem_U87 ( .A(MEM_stage_inst_dmem_n3103), .Z(MEM_stage_inst_dmem_n68) );
BUF_X4 MEM_stage_inst_dmem_U86 ( .A(MEM_stage_inst_dmem_n3209), .Z(MEM_stage_inst_dmem_n67) );
BUF_X4 MEM_stage_inst_dmem_U85 ( .A(MEM_stage_inst_dmem_n4706), .Z(MEM_stage_inst_dmem_n66) );
BUF_X4 MEM_stage_inst_dmem_U84 ( .A(MEM_stage_inst_dmem_n3174), .Z(MEM_stage_inst_dmem_n65) );
BUF_X2 MEM_stage_inst_dmem_U83 ( .A(MEM_stage_inst_dmem_n3170), .Z(MEM_stage_inst_dmem_n64) );
BUF_X4 MEM_stage_inst_dmem_U82 ( .A(MEM_stage_inst_dmem_n7923), .Z(MEM_stage_inst_dmem_n63) );
BUF_X4 MEM_stage_inst_dmem_U81 ( .A(MEM_stage_inst_dmem_n4672), .Z(MEM_stage_inst_dmem_n62) );
BUF_X2 MEM_stage_inst_dmem_U80 ( .A(MEM_stage_inst_dmem_n3130), .Z(MEM_stage_inst_dmem_n61) );
BUF_X4 MEM_stage_inst_dmem_U79 ( .A(MEM_stage_inst_dmem_n3199), .Z(MEM_stage_inst_dmem_n60) );
BUF_X4 MEM_stage_inst_dmem_U78 ( .A(MEM_stage_inst_dmem_n3192), .Z(MEM_stage_inst_dmem_n59) );
BUF_X4 MEM_stage_inst_dmem_U77 ( .A(MEM_stage_inst_dmem_n3155), .Z(MEM_stage_inst_dmem_n58) );
BUF_X4 MEM_stage_inst_dmem_U76 ( .A(MEM_stage_inst_dmem_n3120), .Z(MEM_stage_inst_dmem_n57) );
BUF_X4 MEM_stage_inst_dmem_U75 ( .A(MEM_stage_inst_dmem_n3179), .Z(MEM_stage_inst_dmem_n56) );
BUF_X2 MEM_stage_inst_dmem_U74 ( .A(MEM_stage_inst_dmem_n7937), .Z(MEM_stage_inst_dmem_n55) );
BUF_X4 MEM_stage_inst_dmem_U73 ( .A(MEM_stage_inst_dmem_n4731), .Z(MEM_stage_inst_dmem_n54) );
BUF_X4 MEM_stage_inst_dmem_U72 ( .A(MEM_stage_inst_dmem_n3140), .Z(MEM_stage_inst_dmem_n53) );
BUF_X4 MEM_stage_inst_dmem_U71 ( .A(MEM_stage_inst_dmem_n4710), .Z(MEM_stage_inst_dmem_n52) );
BUF_X2 MEM_stage_inst_dmem_U70 ( .A(MEM_stage_inst_dmem_n3220), .Z(MEM_stage_inst_dmem_n51) );
BUF_X4 MEM_stage_inst_dmem_U69 ( .A(MEM_stage_inst_dmem_n4709), .Z(MEM_stage_inst_dmem_n50) );
BUF_X4 MEM_stage_inst_dmem_U68 ( .A(MEM_stage_inst_dmem_n7960), .Z(MEM_stage_inst_dmem_n49) );
BUF_X4 MEM_stage_inst_dmem_U67 ( .A(MEM_stage_inst_dmem_n3173), .Z(MEM_stage_inst_dmem_n48) );
BUF_X4 MEM_stage_inst_dmem_U66 ( .A(MEM_stage_inst_dmem_n3113), .Z(MEM_stage_inst_dmem_n47) );
BUF_X2 MEM_stage_inst_dmem_U65 ( .A(MEM_stage_inst_dmem_n4740), .Z(MEM_stage_inst_dmem_n46) );
BUF_X4 MEM_stage_inst_dmem_U64 ( .A(MEM_stage_inst_dmem_n7884), .Z(MEM_stage_inst_dmem_n45) );
BUF_X2 MEM_stage_inst_dmem_U63 ( .A(MEM_stage_inst_dmem_n7903), .Z(MEM_stage_inst_dmem_n44) );
BUF_X4 MEM_stage_inst_dmem_U62 ( .A(MEM_stage_inst_dmem_n7888), .Z(MEM_stage_inst_dmem_n43) );
BUF_X4 MEM_stage_inst_dmem_U61 ( .A(MEM_stage_inst_dmem_n4728), .Z(MEM_stage_inst_dmem_n42) );
BUF_X2 MEM_stage_inst_dmem_U60 ( .A(MEM_stage_inst_dmem_n3085), .Z(MEM_stage_inst_dmem_n41) );
BUF_X4 MEM_stage_inst_dmem_U59 ( .A(MEM_stage_inst_dmem_n7938), .Z(MEM_stage_inst_dmem_n40) );
BUF_X2 MEM_stage_inst_dmem_U58 ( .A(MEM_stage_inst_dmem_n4649), .Z(MEM_stage_inst_dmem_n39) );
BUF_X4 MEM_stage_inst_dmem_U57 ( .A(MEM_stage_inst_dmem_n3191), .Z(MEM_stage_inst_dmem_n38) );
BUF_X2 MEM_stage_inst_dmem_U56 ( .A(MEM_stage_inst_dmem_n7992), .Z(MEM_stage_inst_dmem_n37) );
BUF_X2 MEM_stage_inst_dmem_U55 ( .A(MEM_stage_inst_dmem_n3082), .Z(MEM_stage_inst_dmem_n36) );
BUF_X4 MEM_stage_inst_dmem_U54 ( .A(MEM_stage_inst_dmem_n7895), .Z(MEM_stage_inst_dmem_n35) );
BUF_X4 MEM_stage_inst_dmem_U53 ( .A(MEM_stage_inst_dmem_n3163), .Z(MEM_stage_inst_dmem_n34) );
BUF_X4 MEM_stage_inst_dmem_U52 ( .A(MEM_stage_inst_dmem_n4721), .Z(MEM_stage_inst_dmem_n33) );
BUF_X4 MEM_stage_inst_dmem_U51 ( .A(MEM_stage_inst_dmem_n4652), .Z(MEM_stage_inst_dmem_n32) );
BUF_X4 MEM_stage_inst_dmem_U50 ( .A(MEM_stage_inst_dmem_n3112), .Z(MEM_stage_inst_dmem_n31) );
BUF_X4 MEM_stage_inst_dmem_U49 ( .A(MEM_stage_inst_dmem_n4701), .Z(MEM_stage_inst_dmem_n30) );
BUF_X4 MEM_stage_inst_dmem_U48 ( .A(MEM_stage_inst_dmem_n3102), .Z(MEM_stage_inst_dmem_n29) );
BUF_X4 MEM_stage_inst_dmem_U47 ( .A(MEM_stage_inst_dmem_n3152), .Z(MEM_stage_inst_dmem_n28) );
BUF_X4 MEM_stage_inst_dmem_U46 ( .A(MEM_stage_inst_dmem_n7973), .Z(MEM_stage_inst_dmem_n27) );
BUF_X4 MEM_stage_inst_dmem_U45 ( .A(MEM_stage_inst_dmem_n3137), .Z(MEM_stage_inst_dmem_n26) );
BUF_X4 MEM_stage_inst_dmem_U44 ( .A(MEM_stage_inst_dmem_n3217), .Z(MEM_stage_inst_dmem_n25) );
BUF_X4 MEM_stage_inst_dmem_U43 ( .A(MEM_stage_inst_dmem_n3073), .Z(MEM_stage_inst_dmem_n24) );
BUF_X4 MEM_stage_inst_dmem_U42 ( .A(MEM_stage_inst_dmem_n3160), .Z(MEM_stage_inst_dmem_n23) );
BUF_X4 MEM_stage_inst_dmem_U41 ( .A(MEM_stage_inst_dmem_n4769), .Z(MEM_stage_inst_dmem_n22) );
BUF_X4 MEM_stage_inst_dmem_U40 ( .A(MEM_stage_inst_dmem_n3099), .Z(MEM_stage_inst_dmem_n21) );
BUF_X4 MEM_stage_inst_dmem_U39 ( .A(MEM_stage_inst_dmem_n3202), .Z(MEM_stage_inst_dmem_n20) );
BUF_X4 MEM_stage_inst_dmem_U38 ( .A(MEM_stage_inst_dmem_n4667), .Z(MEM_stage_inst_dmem_n19) );
INV_X1 MEM_stage_inst_dmem_U37 ( .A(MEM_stage_inst_dmem_n16), .ZN(MEM_stage_inst_dmem_n18) );
INV_X1 MEM_stage_inst_dmem_U36 ( .A(MEM_stage_inst_dmem_n16), .ZN(MEM_stage_inst_dmem_n17) );
INV_X1 MEM_stage_inst_dmem_U35 ( .A(MEM_stage_inst_dmem_n112), .ZN(MEM_stage_inst_dmem_n16) );
INV_X1 MEM_stage_inst_dmem_U34 ( .A(MEM_stage_inst_dmem_n109), .ZN(MEM_stage_inst_dmem_n13) );
BUF_X1 MEM_stage_inst_dmem_U33 ( .A(MEM_stage_inst_dmem_n20512), .Z(MEM_stage_inst_dmem_n116) );
INV_X4 MEM_stage_inst_dmem_U32 ( .A(MEM_stage_inst_dmem_n11), .ZN(MEM_stage_inst_dmem_n12) );
INV_X1 MEM_stage_inst_dmem_U31 ( .A(MEM_stage_inst_dmem_n116), .ZN(MEM_stage_inst_dmem_n11) );
BUF_X1 MEM_stage_inst_dmem_U30 ( .A(MEM_stage_inst_dmem_n20509), .Z(MEM_stage_inst_dmem_n115) );
INV_X4 MEM_stage_inst_dmem_U29 ( .A(MEM_stage_inst_dmem_n9), .ZN(MEM_stage_inst_dmem_n10) );
INV_X1 MEM_stage_inst_dmem_U28 ( .A(MEM_stage_inst_dmem_n115), .ZN(MEM_stage_inst_dmem_n9) );
INV_X4 MEM_stage_inst_dmem_U26 ( .A(MEM_stage_inst_dmem_n7), .ZN(MEM_stage_inst_dmem_n8) );
INV_X1 MEM_stage_inst_dmem_U25 ( .A(MEM_stage_inst_dmem_n20551), .ZN(MEM_stage_inst_dmem_n7) );
BUF_X1 MEM_stage_inst_dmem_U24 ( .A(EX_pipeline_reg_out_9), .Z(MEM_stage_inst_dmem_n18022) );
INV_X1 MEM_stage_inst_dmem_U23 ( .A(MEM_stage_inst_dmem_n18022), .ZN(MEM_stage_inst_dmem_n5) );
BUF_X1 MEM_stage_inst_dmem_U22 ( .A(MEM_stage_inst_dmem_n13883), .Z(MEM_stage_inst_dmem_n111) );
INV_X2 MEM_stage_inst_dmem_U21 ( .A(MEM_stage_inst_dmem_n3), .ZN(MEM_stage_inst_dmem_n4) );
INV_X1 MEM_stage_inst_dmem_U20 ( .A(MEM_stage_inst_dmem_n111), .ZN(MEM_stage_inst_dmem_n3) );
BUF_X1 MEM_stage_inst_dmem_U18 ( .A(MEM_stage_inst_dmem_n100), .Z(MEM_stage_inst_dmem_n96) );
INV_X2 MEM_stage_inst_dmem_U17 ( .A(MEM_stage_inst_dmem_n1), .ZN(MEM_stage_inst_dmem_n2) );
INV_X1 MEM_stage_inst_dmem_U16 ( .A(MEM_stage_inst_dmem_n96), .ZN(MEM_stage_inst_dmem_n1) );
BUF_X1 MEM_stage_inst_dmem_U14 ( .A(MEM_stage_inst_dmem_n13886), .Z(MEM_stage_inst_dmem_n112) );
BUF_X1 MEM_stage_inst_dmem_U13 ( .A(MEM_stage_inst_dmem_n20547), .Z(MEM_stage_inst_dmem_n109) );
BUF_X4 MEM_stage_inst_dmem_U12 ( .A(EX_pipeline_reg_out_11), .Z(MEM_stage_inst_dmem_n20533) );
BUF_X1 MEM_stage_inst_dmem_U10 ( .A(MEM_stage_inst_dmem_n20506), .Z(MEM_stage_inst_dmem_n14693) );
BUF_X1 MEM_stage_inst_dmem_U9 ( .A(MEM_stage_inst_dmem_n20506), .Z(MEM_stage_inst_dmem_n15110) );
BUF_X1 MEM_stage_inst_dmem_U8 ( .A(MEM_stage_inst_dmem_n20515), .Z(MEM_stage_inst_dmem_n14702) );
BUF_X1 MEM_stage_inst_dmem_U7 ( .A(MEM_stage_inst_dmem_n20518), .Z(MEM_stage_inst_dmem_n14705) );
BUF_X4 MEM_stage_inst_dmem_U6 ( .A(EX_pipeline_reg_out_8), .Z(MEM_stage_inst_dmem_n20541) );
BUF_X4 MEM_stage_inst_dmem_U5 ( .A(EX_pipeline_reg_out_10), .Z(MEM_stage_inst_dmem_n20536) );
INV_X4 MEM_stage_inst_dmem_U4 ( .A(MEM_stage_inst_dmem_n13), .ZN(MEM_stage_inst_dmem_n14) );
INV_X4 MEM_stage_inst_dmem_U3 ( .A(MEM_stage_inst_dmem_n13), .ZN(MEM_stage_inst_dmem_n15) );
endmodule