module s13207 ( g1, g10, g1000, g1006, g1008, g1015, g1016, g1017, g1080, g11, g1193, g1194, g1195, g1196, g1197, g1198, g1201, g1202, g1203, g1205, g1206, g1234, g1246, g1553, g1554, g1724, g1783, g1798, g1804, g1810, g1817, g1824, g1829, g1870, g1871, g1894, g1911, g1944, g206, g21, g22, g23, g24, g25, g26, g2662, g27, g28, g2844, g2888, g29, g291, g30, g3077, g3096, g31, g3130, g3159, g3191, g32, g37, g372, g3829, g3854, g3856, g3857, g3859, g3860, g41, g42, g4267, g43, g4316, g4370, g4371, g4372, g4373, g44, g45, g453, g4655, g4657, g4660, g4661, g4663, g4664, g49, g5143, g5164, g534, g5571, g5669, g5678, g5682, g5684, g5687, g5729, g594, g6207, g6212, g6223, g6236, g6269, g6288, g6289, g6290, g6291, g6292, g6293, g6294, g6295, g6296, g6297, g6298, g6299, g6300, g6301, g6302, g6303, g6304, g6305, g6306, g6307, g6308, g633, g634, g635, g6376, g6425, g645, g647, g648, g6648, g6653, g6675, g6849, g6850, g6895, g690, g6909, g694, g698, g702, g7048, g7063, g7103, g722, g723, g7298, g7423, g7424, g7425, g7474, g7504, g7505, g7506, g7507, g7508, g751, g7514, g752, g753, g754, g755, g756, g757, g7729, g7730, g7731, g7732, g7763, g781, g785, g786, g795, g8216, g8217, g8218, g8219, g8234, g8663, g8872, g8958, g9, g9128, g9132, g9204, g9280, g929, g9297, g9299, g9305, g9308, g9310, g9312, g9314, g9378, g941, g955, g962 , g9116, g6373, g6858, g7116, g6328, g7745, g8871, n1517, g9031, g6855, g9098, g6874, g5745, n1418, g7749, g9086, g7753, g8227, g6385, g6386, g5180, g7735, g6392, g6869, n1522, g5186, g7106, g5737, n1498, g9102, n1509, g7762, g7112, g6365, g6383, g6880, g9085, g7742, g7524, g9029, g9088, g6360, n1518, g9360, n1515, n1485, n1519, g7518, g6349, g5183, g7109, n1416, g7771, g6879, g4654, n1523, g7101, g6352, g7517, g7759, g7772, g7111, g5166, g9097, g9030, g8675, g7113, g8226, g6332, g7302, n1514, g6882, g6316, g8662, g5742, g6317, n1499, g5181, g6353, g9386, g6343, g6851, n1483, g7741, g6330, g8875, g4598, g5736, g6878, g6342, g6891, g6351, g6358, g5173, g5178, g6868, g9114, n1516, n1479, g5185, g8222, g4656, g7512, g7308, g6311, g9107, g5741, g6870, g9034, g8959, g6372, g9090, g6866, g6856, g4665, n1487, g7775, g5739, g8667, g9389, g6345, g7309, g7530, g8224, g7740, g6871, g7299, g5730, g4658, g7304, g9036, g6862, g5163, g7107, g7523, g6388, g6333, g9374, g7733, n1500, g6356, g7743, g6863, g8869, g6380, g9095, g7303, g6873, n1401, n1512, g6354, g5179, g7119, g7305, g5182, g8865, g7110, g6883, g7516, g6357, g6340, g6326, g7525, g7099, g7306, g8665, g9117, g6366, g6889, g8678, g6315, g6852, g7773, g7766, g6337, g6329, g7511, g4668, g7307, g6391, g5170, g9027, g5176, g6344, g3849, g7513, g6312, g5174, g5172, g9115, g7108, g6363, g6374, g9111, g6310, g5177, g6390, g8220, g5738, g6336, g6887, g5732, g6364, g7746, g8956, g6334, g7115, g5175, g6320, g1235, g6379, g6382, g9093, n1521, g7510, g7117, g8957, g8867, g3836, g7118, n1495, g6387, g7768, g7756, g7104, g6362, g7754, g9145, g9091, g9028, g7747, g5168, g5740, g9362, g7100, g7526, g3861, g6369, g7755, g9087, g8674, g5165, g6860, g6319, g7102, n1478, g7737, g8223, g7515, g6861, g7527, g6350, g7105, n1501, g7744, g6377, g6876, g5735, n1407, g9104, g8672, g5731, g6339, g9103, g6359, g7522, g9032, g9100, g6314, g6890, g3863, g7114, g9101, g5184, g9133, g7769, g6865, g6322, g8664, n1520, g6885, g6888, g6886, g7774, n1507, g6325, g7300, g6318, g6355, g6321, g6378, g7529, g6367, g6854, g9109, g7750, g6348, g8676, g6864, g8673, g8666, g7758, g6324, n1489, g7748, g7739, n1493, g5169, g8669, g7520, g6346, g9106, g6884, g3842, g9094, g6313, g9112, g5167, g6338, g9033, g9108, g5743, g9373, g7757, n1491, g6853, g6371, g9372, g8870, g2652, g6881, g9089, g6393, n1497, g6370, g6381, g7761, g5733, g8221, g9099, g7738, g6331, n1481, g7770, g8874, g6384, g9361, g9375, g9092, g7765, g6872, g9376, g7751, g8873, g5187, g9134, g8670, g7767, g6347, g7519, g7764, n1503, g9113, g6335, g7296, g6875, g6323, g6375, g8671, g8225, g9096, g6309, g6857, g7528, g6327, g5746, g6859, g6877, g9110, g6368, g9105, g4669, g3838, g6389, g7752, g9026, g8960, g7521, g8668, g6361, g6867, g5744, g7736, g6341, g8864, g9035, g7301, g71, g12, DFF_635net860, g1179, g5158, g1450, g1360, g462, g1494, g603, g1313, n1404, g995, g1134, DFF_622net847, g435, g154, DFF_619net844, g597, g1351, g381, n1436, g459, g339, g384, g3848, g1204, g866, g411, g162, DFF_605net830, g306, g607, g673, DFF_601net826, g3852, g94, DFF_597net822, g414, g1311, g321, g1158, g432, g324, g539, g584, g1519, g1253, n1439, g1393, g973, g1057, g376, g677, DFF_578net803, g1318, g1118, g765, g300, g521, g258, n1387, g2661, g1155, g1348, g1148, g348, DFF_564net789, g524, DFF_562net787, g5150, g5153, g1330, g1130, n1427, g2673, g3846, n1425, g999, g540, g205, g236, g216, g4659, g764, g395, g1416, g446, g4646, g1159, g1307, g185, g1391, g1191, n1406, g1403, g1514, g1200, g378, g1461, g762, DFF_527net752, g1061, g1106, g3844, g1325, g201, DFF_521net746, g875, DFF_518net743, g4650, g863, g1319, g595, g181, g125, g303, g275, g570, g86, g394, g210, g1398, g1149, g184, g476, g440, g5160, g146, g759, g871, g408, g1329, g950, g1401, g182, g605, g1312, g2663, g616, g591, g121, g874, g489, g1354, g1154, g543, g1097, g1481, g769, g1342, g1142, g734, g714, g1266, g274, g373, g1395, g267, g1033, g4639, g1322, g495, g4641, g1122, g1065, g5155, g601, g1336, n1467, g849, n1437, g429, g5157, g1114, g945, g604, g478, n1426, g2646, n1443, g249, g4651, g630, g610, g108, g547, g507, g1245, g399, g573, g888, g83, g1399, g1199, g233, g213, g602, g618, g377, DFF_422net647, g443, g1069, n1438, g4644, g1270, g2649, g1405, g1005, DFF_412net637, g1176, g953, g356, g4667, g1431, g195, g944, g5146, g492, DFF_402net627, g828, g1192, g599, g837, g129, g1462, n1435, g706, g228, DFF_391net616, g237, g4640, g626, g1409, g556, g1254, g103, g609, DFF_381net606, g47, g2644, g1489, DFF_377net602, g566, g613, g2650, g1402, DFF_371net596, g296, g1310, g1110, g4649, g855, g3855, g477, g1435, g620, g1244, g949, g255, g550, g173, g887, g6841, g628, g345, g456, g933, g336, g316, g617, g1320, g4645, g560, n1385, g93, g1404, g1004, g890, g3845, g770, g1439, g290, g3850, g199, g778, g2653, g536, g516, g261, g852, g68, g375, g1357, g1157, g264, g330, g252, g1053, g1432, DFF_314net539, g4662, g342, g458, g318, g1156, g74, g1390, g501, g623, g553, g1460, g815, g468, g62, g371, g544, g665, g504, g1317, g55, g6843, g1013, g235, g215, g510, g563, g98, g374, g1147, g4599, g405, g436, n1389, g1472, g518, g2660, g859, g773, g150, g5145, g1146, g293, g1327, g831, g77, g661, g627, g158, g4647, DFF_260net485, g557, g231, g834, g211, g309, g92, g1326, DFF_252net477, g1126, g652, g234, g214, g2654, g333, g313, g567, g812, g799, g951, g33, g475, g990, g232, DFF_236net461, g212, g145, g5147, g954, g297, g1041, g998, g402, g1257, g615, g580, g1263, g952, n1448, g1021, g533, DFF_218net443, g513, DFF_215net440, g471, g486, g457, g317, g1467, g588, g1018, g766, g1509, g141, g1396, g474, g1333, g825, DFF_200net425, g104, g4648, g631, g611, g1308, g819, g281, g225, g5149, g5148, g669, g1247, g1430, g614, n1442, g579, g1428, g846, g806, DFF_180net405, g426, g219, g5152, g284, g2664, g5151, g5154, g517, g246, g4642, n1466, g632, g38, g612, g396, g480, g758, n1392, DFF_160net385, DFF_159net384, g959, g760, g186, DFF_155net380, g1045, g99, g4643, g2647, g355, g1087, g685, g174, g768, DFF_144net369, g1025, g822, g583, DFF_140net365, g1185, g1504, g365, g840, g387, DFF_133net358, n1384, g420, g222, g1268, g596, g5156, g479, g240, g200, g1098, g1049, g109, g351, g437, g681, g417, g625, g390, g889, g1309, g1138, g180, g133, g113, g619, g354, g985, g398, g1429, DFF_101net326, g1029, g1389, DFF_98net323, g327, g1412, g646, g52, g1012, g606, g13, n1434, g587, n1386, g3847, g1454, DFF_84net309, g621, g775, g483, g1102, g1037, g295, g730, g710, g763, g270, g362, n1381, g624, g179, DFF_68net293, g3851, g598, g718, DFF_63net288, g278, g1513, g527, g137, g117, g984, g1014, g2651, g622, g2648, g455, g315, g843, g803, g771, g423, g600, g1269, g1444, g80, g1499, g243, g1304, g2645, g774, g465, g608, n1447, g1477, g294, g2659, g1077, g393, g767, g2672, g20, g1339, DFF_24net249, g359, g183, I8024, g772, g292, g535, g5159, g454, g1092, g314, g498, g976, g940, g1153, g5161, g629, g948, g452, g273, g312, g1271, g397, DFF_20net245 );
input g1, g10, g1000, g1008, g1016, g1080, g11, g1194, g1196, g1198, g1202, g1203, g1206, g1234, g1553, g1554, g21, g22, g23, g24, g25, g26, g27, g28, g29, g30, g31, g32, g37, g41, g42, g43, g44, g45, g49, g633, g634, g635, g645, g647, g648, g690, g694, g698, g702, g722, g723, g751, g752, g753, g754, g755, g756, g757, g781, g786, g795, g9, g929, g941, g955, g962, g4370, g1193, g7423, g2844, g7424, g4373, g1871, g1911, g1944, g1195, g4267, g1870, g5571, g3130, g3096, g2888, g4371, g3191, g1197, g3159, g7425, g6223, g1201, g4316, g4372, g1205, g71, g12, DFF_635net860, g1179, g5158, g1450, g1360, g462, g1494, g603, g1313, n1404, g995, g1134, DFF_622net847, g435, g154, DFF_619net844, g597, g1351, g381, n1436, g459, g339, g384, g3848, g1204, g866, g411, g162, DFF_605net830, g306, g607, g673, DFF_601net826, g3852, g94, DFF_597net822, g414, g1311, g321, g1158, g432, g324, g539, g584, g1519, g1253, n1439, g1393, g973, g1057, g376, g677, DFF_578net803, g1318, g1118, g765, g300, g521, g258, n1387, g2661, g1155, g1348, g1148, g348, DFF_564net789, g524, DFF_562net787, g5150, g5153, g1330, g1130, n1427, g2673, g3846, n1425, g999, g540, g205, g236, g216, g4659, g764, g395, g1416, g446, g4646, g1159, g1307, g185, g1391, g1191, n1406, g1403, g1514, g1200, g378, g1461, g762, DFF_527net752, g1061, g1106, g3844, g1325, g201, DFF_521net746, g875, DFF_518net743, g4650, g863, g1319, g595, g181, g125, g303, g275, g570, g86, g394, g210, g1398, g1149, g184, g476, g440, g5160, g146, g759, g871, g408, g1329, g950, g1401, g182, g605, g1312, g2663, g616, g591, g121, g874, g489, g1354, g1154, g543, g1097, g1481, g769, g1342, g1142, g734, g714, g1266, g274, g373, g1395, g267, g1033, g4639, g1322, g495, g4641, g1122, g1065, g5155, g601, g1336, n1467, g849, n1437, g429, g5157, g1114, g945, g604, g478, n1426, g2646, n1443, g249, g4651, g630, g610, g108, g547, g507, g1245, g399, g573, g888, g83, g1399, g1199, g233, g213, g602, g618, g377, DFF_422net647, g443, g1069, n1438, g4644, g1270, g2649, g1405, g1005, DFF_412net637, g1176, g953, g356, g4667, g1431, g195, g944, g5146, g492, DFF_402net627, g828, g1192, g599, g837, g129, g1462, n1435, g706, g228, DFF_391net616, g237, g4640, g626, g1409, g556, g1254, g103, g609, DFF_381net606, g47, g2644, g1489, DFF_377net602, g566, g613, g2650, g1402, DFF_371net596, g296, g1310, g1110, g4649, g855, g3855, g477, g1435, g620, g1244, g949, g255, g550, g173, g887, g6841, g628, g345, g456, g933, g336, g316, g617, g1320, g4645, g560, n1385, g93, g1404, g1004, g890, g3845, g770, g1439, g290, g3850, g199, g778, g2653, g536, g516, g261, g852, g68, g375, g1357, g1157, g264, g330, g252, g1053, g1432, DFF_314net539, g4662, g342, g458, g318, g1156, g74, g1390, g501, g623, g553, g1460, g815, g468, g62, g371, g544, g665, g504, g1317, g55, g6843, g1013, g235, g215, g510, g563, g98, g374, g1147, g4599, g405, g436, n1389, g1472, g518, g2660, g859, g773, g150, g5145, g1146, g293, g1327, g831, g77, g661, g627, g158, g4647, DFF_260net485, g557, g231, g834, g211, g309, g92, g1326, DFF_252net477, g1126, g652, g234, g214, g2654, g333, g313, g567, g812, g799, g951, g33, g475, g990, g232, DFF_236net461, g212, g145, g5147, g954, g297, g1041, g998, g402, g1257, g615, g580, g1263, g952, n1448, g1021, g533, DFF_218net443, g513, DFF_215net440, g471, g486, g457, g317, g1467, g588, g1018, g766, g1509, g141, g1396, g474, g1333, g825, DFF_200net425, g104, g4648, g631, g611, g1308, g819, g281, g225, g5149, g5148, g669, g1247, g1430, g614, n1442, g579, g1428, g846, g806, DFF_180net405, g426, g219, g5152, g284, g2664, g5151, g5154, g517, g246, g4642, n1466, g632, g38, g612, g396, g480, g758, n1392, DFF_160net385, DFF_159net384, g959, g760, g186, DFF_155net380, g1045, g99, g4643, g2647, g355, g1087, g685, g174, g768, DFF_144net369, g1025, g822, g583, DFF_140net365, g1185, g1504, g365, g840, g387, DFF_133net358, n1384, g420, g222, g1268, g596, g5156, g479, g240, g200, g1098, g1049, g109, g351, g437, g681, g417, g625, g390, g889, g1309, g1138, g180, g133, g113, g619, g354, g985, g398, g1429, DFF_101net326, g1029, g1389, DFF_98net323, g327, g1412, g646, g52, g1012, g606, g13, n1434, g587, n1386, g3847, g1454, DFF_84net309, g621, g775, g483, g1102, g1037, g295, g730, g710, g763, g270, g362, n1381, g624, g179, DFF_68net293, g3851, g598, g718, DFF_63net288, g278, g1513, g527, g137, g117, g984, g1014, g2651, g622, g2648, g455, g315, g843, g803, g771, g423, g600, g1269, g1444, g80, g1499, g243, g1304, g2645, g774, g465, g608, n1447, g1477, g294, g2659, g1077, g393, g767, g2672, g20, g1339, DFF_24net249, g359, g183, I8024, g772, g292, g535, g5159, g454, g1092, g314, g498, g976, g940, g1153, g5161, g629, g948, g452, g273, g312, g1271, g397, DFF_20net245;
output g1006, g1015, g1017, g1246, g1724, g1783, g1798, g1804, g1810, g1817, g1824, g1829, g1894, g206, g2662, g291, g3077, g372, g3829, g3854, g3856, g3857, g3859, g3860, g453, g4655, g4657, g4660, g4661, g4663, g4664, g5143, g5164, g534, g5669, g5678, g5682, g5684, g5687, g5729, g594, g6207, g6212, g6236, g6269, g6288, g6289, g6290, g6291, g6292, g6293, g6294, g6295, g6296, g6297, g6298, g6299, g6300, g6301, g6302, g6303, g6304, g6305, g6306, g6307, g6308, g6376, g6425, g6648, g6653, g6675, g6849, g6850, g6895, g6909, g7048, g7063, g7103, g7298, g7474, g7504, g7505, g7506, g7507, g7508, g7514, g7729, g7730, g7731, g7732, g7763, g785, g8216, g8217, g8218, g8219, g8234, g8663, g8872, g8958, g9128, g9132, g9204, g9280, g9297, g9299, g9305, g9308, g9310, g9312, g9314, g9378, g9116, g6373, g6858, g7116, g6328, g7745, g8871, n1517, g9031, g6855, g9098, g6874, g5745, n1418, g7749, g9086, g7753, g8227, g6385, g6386, g5180, g7735, g6392, g6869, n1522, g5186, g7106, g5737, n1498, g9102, n1509, g7762, g7112, g6365, g6383, g6880, g9085, g7742, g7524, g9029, g9088, g6360, n1518, g9360, n1515, n1485, n1519, g7518, g6349, g5183, g7109, n1416, g7771, g6879, g4654, n1523, g7101, g6352, g7517, g7759, g7772, g7111, g5166, g9097, g9030, g8675, g7113, g8226, g6332, g7302, n1514, g6882, g6316, g8662, g5742, g6317, n1499, g5181, g6353, g9386, g6343, g6851, n1483, g7741, g6330, g8875, g4598, g5736, g6878, g6342, g6891, g6351, g6358, g5173, g5178, g6868, g9114, n1516, n1479, g5185, g8222, g4656, g7512, g7308, g6311, g9107, g5741, g6870, g9034, g8959, g6372, g9090, g6866, g6856, g4665, n1487, g7775, g5739, g8667, g9389, g6345, g7309, g7530, g8224, g7740, g6871, g7299, g5730, g4658, g7304, g9036, g6862, g5163, g7107, g7523, g6388, g6333, g9374, g7733, n1500, g6356, g7743, g6863, g8869, g6380, g9095, g7303, g6873, n1401, n1512, g6354, g5179, g7119, g7305, g5182, g8865, g7110, g6883, g7516, g6357, g6340, g6326, g7525, g7099, g7306, g8665, g9117, g6366, g6889, g8678, g6315, g6852, g7773, g7766, g6337, g6329, g7511, g4668, g7307, g6391, g5170, g9027, g5176, g6344, g3849, g7513, g6312, g5174, g5172, g9115, g7108, g6363, g6374, g9111, g6310, g5177, g6390, g8220, g5738, g6336, g6887, g5732, g6364, g7746, g8956, g6334, g7115, g5175, g6320, g1235, g6379, g6382, g9093, n1521, g7510, g7117, g8957, g8867, g3836, g7118, n1495, g6387, g7768, g7756, g7104, g6362, g7754, g9145, g9091, g9028, g7747, g5168, g5740, g9362, g7100, g7526, g3861, g6369, g7755, g9087, g8674, g5165, g6860, g6319, g7102, n1478, g7737, g8223, g7515, g6861, g7527, g6350, g7105, n1501, g7744, g6377, g6876, g5735, n1407, g9104, g8672, g5731, g6339, g9103, g6359, g7522, g9032, g9100, g6314, g6890, g3863, g7114, g9101, g5184, g9133, g7769, g6865, g6322, g8664, n1520, g6885, g6888, g6886, g7774, n1507, g6325, g7300, g6318, g6355, g6321, g6378, g7529, g6367, g6854, g9109, g7750, g6348, g8676, g6864, g8673, g8666, g7758, g6324, n1489, g7748, g7739, n1493, g5169, g8669, g7520, g6346, g9106, g6884, g3842, g9094, g6313, g9112, g5167, g6338, g9033, g9108, g5743, g9373, g7757, n1491, g6853, g6371, g9372, g8870, g2652, g6881, g9089, g6393, n1497, g6370, g6381, g7761, g5733, g8221, g9099, g7738, g6331, n1481, g7770, g8874, g6384, g9361, g9375, g9092, g7765, g6872, g9376, g7751, g8873, g5187, g9134, g8670, g7767, g6347, g7519, g7764, n1503, g9113, g6335, g7296, g6875, g6323, g6375, g8671, g8225, g9096, g6309, g6857, g7528, g6327, g5746, g6859, g6877, g9110, g6368, g9105, g4669, g3838, g6389, g7752, g9026, g8960, g7521, g8668, g6361, g6867, g5744, g7736, g6341, g8864, g9035, g7301;
wire g1000, g1008, g11, g1554, g21, g25, g30, g31, g32, g41, g42, g44, g49, g9, g8955, g7509, g7071, g9291, g8625, g6745, g8627, g9261, g3528, g7252, I5528, g9285, g1683, g9264, g9288, g7322, g8633, g9267, g6056, g6952, g7248, g2801, g9363, g6565, g8630, g3084, g9282, g2474, g3516, g3555, g4302, g3505, g3504, g9294, n1379, n1380, n1382, n1383, n1388, n1390, n1391, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1402, n1403, n1405, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1417, n1419, n1420, n1421, n1422, n1423, n1424, n1428, n1429, n1430, n1431, n1432, n1433, n1440, n1441, n1444, n1445, n1446, n1449, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1477, n1480, n1482, n1484, n1486, n1488, n1490, n1492, n1494, n1496, n1502, n1504, n1505, n1506, n1508, n1510, n1511, n1513, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, DFF_630net855 , DFF_576net801 , DFF_550net775 , DFF_517net742 , DFF_404net629 , DFF_373net598 , DFF_365net590 , DFF_342net567 , DFF_313net538 , DFF_286net511 , DFF_270net495 , DFF_175net400 , DFF_171net396 , DFF_166net391 , DFF_66net291;
nb1s1 U3371 ( .Q(g6269), .DIN(g1000) );
nb1s1 U3372 ( .Q(g6909), .DIN(g1008) );
nb1s1 U3373 ( .Q(g6290), .DIN(g11) );
nb1s1 U3374 ( .Q(g5143), .DIN(g1554) );
nb1s1 U3375 ( .Q(g6299), .DIN(g21) );
nb1s1 U3376 ( .Q(g6376), .DIN(g25) );
nb1s1 U3377 ( .Q(g6295), .DIN(g25) );
nb1s1 U3378 ( .Q(g6301), .DIN(g30) );
nb1s1 U3379 ( .Q(g6302), .DIN(g31) );
nb1s1 U3380 ( .Q(g6303), .DIN(g32) );
nb1s1 U3381 ( .Q(g6305), .DIN(g41) );
nb1s1 U3382 ( .Q(g6306), .DIN(g42) );
nb1s1 U3383 ( .Q(g6307), .DIN(g44) );
nb1s1 U3384 ( .Q(g5729), .DIN(g49) );
nb1s1 U3385 ( .Q(g6288), .DIN(g9) );
nb1s1 U3386 ( .Q(g6291), .DIN(g6309) );
nb1s1 U3387 ( .Q(g6309), .DIN(g10) );
nb1s1 U3388 ( .Q(g7506), .DIN(g20) );
nb1s1 U3389 ( .Q(g5682), .DIN(g20) );
nb1s1 U3390 ( .Q(g1810), .DIN(g2647) );
nb1s1 U3391 ( .Q(g7504), .DIN(g13) );
nb1s1 U3392 ( .Q(g5669), .DIN(g13) );
nb1s1 U3393 ( .Q(g6851), .DIN(g43) );
nb1s1 U3394 ( .Q(g7730), .DIN(g1389) );
nb1s1 U3395 ( .Q(g6212), .DIN(g1389) );
nb1s1 U3396 ( .Q(g3077), .DIN(g1029) );
nb1s1 U3397 ( .Q(g1017), .DIN(g1029) );
nb1s1 U3398 ( .Q(g1817), .DIN(g2648) );
nb1s1 U3399 ( .Q(g7508), .DIN(g38) );
nb1s1 U3400 ( .Q(g5687), .DIN(g38) );
nb1s1 U3401 ( .Q(g1804), .DIN(g2646) );
nb1s1 U3402 ( .Q(g8217), .DIN(g4662) );
nb1s1 U3403 ( .Q(g6653), .DIN(g4662) );
nb1s1 U3404 ( .Q(g6298), .DIN(g6389) );
nb1s1 U3405 ( .Q(g6389), .DIN(g28) );
nb1s1 U3406 ( .Q(g6308), .DIN(g8955) );
nb1s1 U3407 ( .Q(g8955), .DIN(g45) );
nb1s1 U3408 ( .Q(g7507), .DIN(g33) );
nb1s1 U3409 ( .Q(g5684), .DIN(g33) );
nb1s1 U3410 ( .Q(g6300), .DIN(g6390) );
nb1s1 U3411 ( .Q(g6390), .DIN(g29) );
nb1s1 U3412 ( .Q(g1829), .DIN(g2650) );
nb1s1 U3413 ( .Q(g1783), .DIN(g2651) );
nb1s1 U3414 ( .Q(g1235), .DIN(g1234) );
nb1s1 U3415 ( .Q(g3842), .DIN(g1202) );
nb1s1 U3416 ( .Q(g594), .DIN(g1460) );
nb1s1 U3417 ( .Q(g534), .DIN(g1460) );
nb1s1 U3418 ( .Q(g453), .DIN(g1460) );
nb1s1 U3419 ( .Q(g372), .DIN(g1460) );
nb1s1 U3420 ( .Q(g291), .DIN(g1460) );
nb1s1 U3421 ( .Q(g206), .DIN(g1460) );
nb1s1 U3422 ( .Q(g8216), .DIN(g4659) );
nb1s1 U3423 ( .Q(g6648), .DIN(g4659) );
nb1s1 U3424 ( .Q(g3836), .DIN(g1194) );
nb1s1 U3425 ( .Q(g7729), .DIN(g173) );
nb1s1 U3426 ( .Q(g6207), .DIN(g173) );
nb1s1 U3427 ( .Q(g3838), .DIN(g1198) );
nb1s1 U3428 ( .Q(g6297), .DIN(g6388) );
nb1s1 U3429 ( .Q(g6388), .DIN(g27) );
nb1s1 U3430 ( .Q(g2662), .DIN(g1254) );
nb1s1 U3431 ( .Q(g1724), .DIN(g1409) );
nb1s1 U3432 ( .Q(g2652), .DIN(g941) );
nb1s1 U3433 ( .Q(g1824), .DIN(g2649) );
nb1s1 U3434 ( .Q(g6296), .DIN(g6387) );
nb1s1 U3435 ( .Q(g6387), .DIN(g26) );
nb1s1 U3436 ( .Q(g6294), .DIN(g6375) );
nb1s1 U3437 ( .Q(g6375), .DIN(g24) );
nb1s1 U3438 ( .Q(g7731), .DIN(g3861) );
nb1s1 U3439 ( .Q(g6236), .DIN(g3861) );
nb1s1 U3440 ( .Q(g785), .DIN(g888) );
nb1s1 U3441 ( .Q(g1246), .DIN(g1245) );
nb1s1 U3442 ( .Q(g1798), .DIN(g2645) );
nb1s1 U3443 ( .Q(g6293), .DIN(g6374) );
nb1s1 U3444 ( .Q(g6374), .DIN(g23) );
nb1s1 U3445 ( .Q(g6289), .DIN(g6310) );
nb1s1 U3446 ( .Q(g6310), .DIN(g1) );
nb1s1 U3447 ( .Q(g6304), .DIN(g6393) );
nb1s1 U3448 ( .Q(g6393), .DIN(g37) );
nb1s1 U3449 ( .Q(g3860), .DIN(g1461) );
nb1s1 U3450 ( .Q(g3859), .DIN(g1461) );
nb1s1 U3451 ( .Q(g3829), .DIN(g1461) );
nb1s1 U3452 ( .Q(g6292), .DIN(g6373) );
nb1s1 U3453 ( .Q(g6373), .DIN(g22) );
nb1s1 U3454 ( .Q(g8218), .DIN(g4599) );
nb1s1 U3455 ( .Q(g6425), .DIN(g4599) );
nb1s1 U3456 ( .Q(g3849), .DIN(g1206) );
nb1s1 U3457 ( .Q(g1894), .DIN(g2660) );
nb1s1 U3458 ( .Q(g7505), .DIN(g2664) );
nb1s1 U3459 ( .Q(g5678), .DIN(g2664) );
nb1s1 U3460 ( .Q(g7048), .DIN(g8662) );
nb1s1 U3461 ( .Q(g7298), .DIN(g7071) );
nb1s1 U3462 ( .Q(g9312), .DIN(g9291) );
nb1s1 U3463 ( .Q(g6895), .DIN(I8024) );
nb1s1 U3464 ( .Q(g1006), .DIN(g8625) );
nb1s1 U3465 ( .Q(g7103), .DIN(g6745) );
nb1s1 U3466 ( .Q(g8958), .DIN(g8627) );
nb1s1 U3467 ( .Q(g9280), .DIN(g9261) );
nb1s1 U3468 ( .Q(g4660), .DIN(g3528) );
nb1s1 U3469 ( .Q(g7514), .DIN(g7252) );
nb1s1 U3470 ( .Q(g6850), .DIN(I5528) );
nb1s1 U3471 ( .Q(g9308), .DIN(g9285) );
nb1s1 U3472 ( .Q(g3854), .DIN(g1683) );
nb1s1 U3473 ( .Q(g9297), .DIN(g9264) );
nb1s1 U3474 ( .Q(g9310), .DIN(g9288) );
nb1s1 U3475 ( .Q(g7763), .DIN(g7322) );
nb1s1 U3476 ( .Q(g8872), .DIN(g8633) );
nb1s1 U3477 ( .Q(g9299), .DIN(g9267) );
nb1s1 U3478 ( .Q(g6849), .DIN(g6056) );
nb1s1 U3479 ( .Q(g9204), .DIN(g6952) );
nb1s1 U3480 ( .Q(g9128), .DIN(g6952) );
nb1s1 U3481 ( .Q(g7474), .DIN(g7248) );
nb1s1 U3482 ( .Q(g4655), .DIN(g2801) );
nb1s1 U3483 ( .Q(g9378), .DIN(g9363) );
nb1s1 U3484 ( .Q(g9132), .DIN(g6565) );
nb1s1 U3485 ( .Q(g8234), .DIN(g6565) );
nb1s1 U3486 ( .Q(g1015), .DIN(g8630) );
nb1s1 U3487 ( .Q(g3857), .DIN(g3084) );
nb1s1 U3488 ( .Q(g9305), .DIN(g9282) );
nb1s1 U3489 ( .Q(g8663), .DIN(g2474) );
nb1s1 U3490 ( .Q(g7063), .DIN(g2474) );
nb1s1 U3491 ( .Q(g4664), .DIN(g3516) );
nb1s1 U3492 ( .Q(g4663), .DIN(g3555) );
nb1s1 U3493 ( .Q(g5164), .DIN(g4302) );
nb1s1 U3494 ( .Q(g4661), .DIN(g3505) );
nb1s1 U3495 ( .Q(g4657), .DIN(g3504) );
nb1s1 U3496 ( .Q(g9314), .DIN(g9294) );
nb1s1 U3497 ( .Q(g7732), .DIN(g6223) );
nb1s1 U3498 ( .Q(g8219), .DIN(g6675) );
and2s1 U1791 ( .Q(g7739), .DIN1(g154), .DIN2(DFF_133net358) );
hi1s1 U1792 ( .Q(g7741), .DIN(n2189) );
hi1s1 U1793 ( .Q(n2189), .DIN(g162) );
hi1s1 U1794 ( .Q(g7746), .DIN(n2184) );
hi1s1 U1795 ( .Q(n2184), .DIN(g673) );
hi1s1 U1796 ( .Q(g7747), .DIN(n2183) );
hi1s1 U1797 ( .Q(n2183), .DIN(g677) );
hi1s1 U1798 ( .Q(g8222), .DIN(n2118) );
hi1s1 U1799 ( .Q(n2118), .DIN(n2119) );
hi1s1 U1800 ( .Q(g7735), .DIN(n2194) );
hi1s1 U1801 ( .Q(n2194), .DIN(g146) );
hi1s1 U1802 ( .Q(g7755), .DIN(n2174) );
hi1s1 U1803 ( .Q(n2174), .DIN(g734) );
hi1s1 U1804 ( .Q(g7752), .DIN(n2177) );
hi1s1 U1805 ( .Q(n2177), .DIN(g714) );
hi1s1 U1806 ( .Q(g4598), .DIN(n1443) );
hi1s1 U1807 ( .Q(g8956), .DIN(n2038) );
hi1s1 U1808 ( .Q(n2038), .DIN(n2039) );
hi1s1 U1809 ( .Q(g7750), .DIN(n2180) );
hi1s1 U1810 ( .Q(n2180), .DIN(g706) );
hi1s1 U1811 ( .Q(g8220), .DIN(n2121) );
hi1s1 U1812 ( .Q(n2121), .DIN(g855) );
hi1s1 U1813 ( .Q(g7736), .DIN(n2193) );
hi1s1 U1814 ( .Q(n2193), .DIN(g173) );
hi1s1 U1815 ( .Q(g7744), .DIN(n2186) );
hi1s1 U1816 ( .Q(n2186), .DIN(g665) );
hi1s1 U1817 ( .Q(g8221), .DIN(n2120) );
hi1s1 U1818 ( .Q(n2120), .DIN(g859) );
hi1s1 U1819 ( .Q(g7738), .DIN(n2191) );
hi1s1 U1820 ( .Q(n2191), .DIN(g150) );
hi1s1 U1821 ( .Q(g7743), .DIN(n2187) );
hi1s1 U1822 ( .Q(n2187), .DIN(g661) );
hi1s1 U1823 ( .Q(g7740), .DIN(n2190) );
hi1s1 U1824 ( .Q(n2190), .DIN(g158) );
hi1s1 U1825 ( .Q(g7742), .DIN(n2188) );
hi1s1 U1826 ( .Q(n2188), .DIN(g2654) );
hi1s1 U1827 ( .Q(g7745), .DIN(n2185) );
hi1s1 U1828 ( .Q(n2185), .DIN(g669) );
hi1s1 U1829 ( .Q(g7749), .DIN(n2181) );
hi1s1 U1830 ( .Q(n2181), .DIN(g685) );
hi1s1 U1831 ( .Q(g7737), .DIN(n2192) );
hi1s1 U1832 ( .Q(n2192), .DIN(g174) );
hi1s1 U1833 ( .Q(g7748), .DIN(n2182) );
hi1s1 U1834 ( .Q(n2182), .DIN(g681) );
hi1s1 U1835 ( .Q(g9386), .DIN(n1524) );
hi1s1 U1836 ( .Q(n1524), .DIN(n1525) );
hi1s1 U1837 ( .Q(g7754), .DIN(n2175) );
hi1s1 U1838 ( .Q(n2175), .DIN(g730) );
hi1s1 U1839 ( .Q(g7751), .DIN(n2178) );
hi1s1 U1840 ( .Q(n2178), .DIN(g710) );
hi1s1 U1841 ( .Q(g7753), .DIN(n2176) );
hi1s1 U1842 ( .Q(n2176), .DIN(g718) );
hi1s1 U1843 ( .Q(n1478), .DIN(n1477) );
hi1s1 U1844 ( .Q(n1479), .DIN(n1543) );
hi1s1 U1845 ( .Q(n1481), .DIN(n1480) );
hi1s1 U1846 ( .Q(n1483), .DIN(n1482) );
hi1s1 U1847 ( .Q(n1485), .DIN(n1484) );
hi1s1 U1848 ( .Q(n1487), .DIN(n1486) );
hi1s1 U1849 ( .Q(n1489), .DIN(n1488) );
hi1s1 U1850 ( .Q(n1491), .DIN(n1490) );
hi1s1 U1851 ( .Q(n1493), .DIN(n1492) );
hi1s1 U1852 ( .Q(n1495), .DIN(n1494) );
hi1s1 U1853 ( .Q(n1497), .DIN(n1496) );
hi1s1 U1854 ( .Q(n1498), .DIN(n1447) );
hi1s1 U1855 ( .Q(n1499), .DIN(n1447) );
hi1s1 U1856 ( .Q(n1500), .DIN(n1428) );
hi1s1 U1857 ( .Q(n1501), .DIN(n1428) );
hi1s1 U1858 ( .Q(n1503), .DIN(n1502) );
hi1s1 U1859 ( .Q(n1505), .DIN(n1504) );
hi1s1 U1860 ( .Q(n1507), .DIN(n1506) );
hi1s1 U1861 ( .Q(n1509), .DIN(n1508) );
hi1s1 U1862 ( .Q(n1510), .DIN(n1944) );
hi1s1 U1863 ( .Q(n1512), .DIN(n1511) );
hi1s1 U1864 ( .Q(n1514), .DIN(n1513) );
hi1s1 U1865 ( .Q(n1515), .DIN(n1429) );
hi1s1 U1866 ( .Q(n1516), .DIN(n1412) );
hi1s1 U1867 ( .Q(n1517), .DIN(n1412) );
hi1s1 U1868 ( .Q(n1520), .DIN(n1414) );
hi1s1 U1869 ( .Q(n1518), .DIN(n1414) );
hi1s1 U1870 ( .Q(n1519), .DIN(n1414) );
hi1s1 U1871 ( .Q(n1521), .DIN(n1413) );
hi1s1 U1872 ( .Q(n1523), .DIN(n1413) );
hi1s1 U1873 ( .Q(n1522), .DIN(n1413) );
nnd2s1 U1886 ( .Q(n1525), .DIN1(n1434), .DIN2(n1526) );
nnd4s1 U1887 ( .Q(n1526), .DIN1(g9389), .DIN2(n1527), .DIN3(n1528), .DIN4(n1529) );
nor2s1 U1888 ( .Q(n1528), .DIN1(g8955), .DIN2(g44) );
or2s1 U1889 ( .Q(g9363), .DIN1(n1388), .DIN2(g9389) );
nnd2s1 U1890 ( .Q(g9389), .DIN1(n1530), .DIN2(n1531) );
nnd2s1 U1891 ( .Q(n1531), .DIN1(n1532), .DIN2(g44) );
xor2s1 U1892 ( .Q(n1532), .DIN1(n1533), .DIN2(n1534) );
xor2s1 U1893 ( .Q(n1534), .DIN1(n1535), .DIN2(n1536) );
xor2s1 U1894 ( .Q(n1536), .DIN1(g9375), .DIN2(n1537) );
xor2s1 U1895 ( .Q(n1535), .DIN1(g9376), .DIN2(g9374) );
xor2s1 U1896 ( .Q(n1533), .DIN1(n1538), .DIN2(n1539) );
xor2s1 U1897 ( .Q(n1539), .DIN1(g9373), .DIN2(g9372) );
xor2s1 U1898 ( .Q(n1538), .DIN1(g9360), .DIN2(g9362) );
or3s1 U1899 ( .Q(n1530), .DIN1(n1540), .DIN2(n1541), .DIN3(g44) );
hi1s1 U1900 ( .Q(g9361), .DIN(n1537) );
or2s1 U1901 ( .Q(g9294), .DIN1(n1388), .DIN2(g9376) );
or4s1 U1902 ( .Q(g9376), .DIN1(n1542), .DIN2(n1543), .DIN3(n1544), .DIN4(n1545) );
nnd4s1 U1903 ( .Q(n1545), .DIN1(n1546), .DIN2(n1547), .DIN3(n1548), .DIN4(n1549) );
and3s1 U1904 ( .Q(n1549), .DIN1(n1550), .DIN2(n1551), .DIN3(n1552) );
nnd2s1 U1905 ( .Q(n1552), .DIN1(g255), .DIN2(n1553) );
nnd2s1 U1906 ( .Q(n1551), .DIN1(g614), .DIN2(n1554) );
nnd2s1 U1907 ( .Q(n1550), .DIN1(g336), .DIN2(n1555) );
nnd2s1 U1908 ( .Q(n1548), .DIN1(g563), .DIN2(n1556) );
nnd2s1 U1909 ( .Q(n1547), .DIN1(n1557), .DIN2(n1558) );
nnd4s1 U1910 ( .Q(n1558), .DIN1(n1559), .DIN2(n1560), .DIN3(n1561), .DIN4(n1562) );
nor2s1 U1911 ( .Q(n1562), .DIN1(n1563), .DIN2(n1564) );
and2s1 U1912 ( .Q(n1564), .DIN1(n1565), .DIN2(g767) );
and2s1 U1913 ( .Q(n1563), .DIN1(n1566), .DIN2(g759) );
nnd2s1 U1914 ( .Q(n1561), .DIN1(g831), .DIN2(n1567) );
nnd2s1 U1915 ( .Q(n1560), .DIN1(n1568), .DIN2(n1569) );
nnd4s1 U1916 ( .Q(n1569), .DIN1(n1570), .DIN2(n1571), .DIN3(n1572), .DIN4(n1573) );
nor2s1 U1917 ( .Q(n1573), .DIN1(n1574), .DIN2(n1575) );
and2s1 U1918 ( .Q(n1575), .DIN1(n1576), .DIN2(g690) );
and2s1 U1919 ( .Q(n1574), .DIN1(n1577), .DIN2(g706) );
nnd2s1 U1920 ( .Q(n1572), .DIN1(g498), .DIN2(n1578) );
nnd2s1 U1921 ( .Q(n1570), .DIN1(g751), .DIN2(n1579) );
nnd2s1 U1922 ( .Q(n1559), .DIN1(n1580), .DIN2(n1512) );
nnd2s1 U1923 ( .Q(n1546), .DIN1(g417), .DIN2(n1581) );
nnd3s1 U1924 ( .Q(n1544), .DIN1(n1582), .DIN2(n1583), .DIN3(n1584) );
nnd2s1 U1925 ( .Q(n1584), .DIN1(g5153), .DIN2(n1585) );
nnd2s1 U1926 ( .Q(n1583), .DIN1(g601), .DIN2(n1586) );
nnd2s1 U1927 ( .Q(n1582), .DIN1(g625), .DIN2(n1587) );
hi1s1 U1928 ( .Q(n1543), .DIN(g7509) );
and2s1 U1929 ( .Q(n1542), .DIN1(n1588), .DIN2(g146) );
or2s1 U1930 ( .Q(g9291), .DIN1(n1388), .DIN2(g9375) );
or3s1 U1931 ( .Q(g9375), .DIN1(n1589), .DIN2(n1590), .DIN3(n1591) );
nnd4s1 U1932 ( .Q(n1591), .DIN1(n1592), .DIN2(n1593), .DIN3(n1594), .DIN4(n1595) );
and3s1 U1933 ( .Q(n1595), .DIN1(n1596), .DIN2(n1597), .DIN3(n1598) );
nnd2s1 U1934 ( .Q(n1598), .DIN1(g183), .DIN2(n1599) );
nnd2s1 U1935 ( .Q(n1597), .DIN1(g615), .DIN2(n1554) );
nnd2s1 U1936 ( .Q(n1596), .DIN1(g339), .DIN2(n1555) );
nnd2s1 U1937 ( .Q(n1594), .DIN1(g570), .DIN2(n1556) );
nnd2s1 U1938 ( .Q(n1593), .DIN1(n1557), .DIN2(n1600) );
nnd4s1 U1939 ( .Q(n1600), .DIN1(n1601), .DIN2(n1602), .DIN3(n1603), .DIN4(n1604) );
nor2s1 U1940 ( .Q(n1604), .DIN1(n1605), .DIN2(n1606) );
and2s1 U1941 ( .Q(n1606), .DIN1(n1565), .DIN2(g768) );
and2s1 U1942 ( .Q(n1605), .DIN1(n1566), .DIN2(g760) );
nnd2s1 U1943 ( .Q(n1603), .DIN1(g834), .DIN2(n1567) );
nnd2s1 U1944 ( .Q(n1602), .DIN1(n1568), .DIN2(n1607) );
nnd4s1 U1945 ( .Q(n1607), .DIN1(n1608), .DIN2(n1571), .DIN3(n1609), .DIN4(n1610) );
nor2s1 U1946 ( .Q(n1610), .DIN1(n1611), .DIN2(n1612) );
and2s1 U1947 ( .Q(n1612), .DIN1(n1576), .DIN2(g633) );
and2s1 U1948 ( .Q(n1611), .DIN1(n1577), .DIN2(g661) );
nnd2s1 U1949 ( .Q(n1609), .DIN1(g501), .DIN2(n1578) );
nnd2s1 U1950 ( .Q(n1608), .DIN1(g755), .DIN2(n1579) );
nnd2s1 U1951 ( .Q(n1601), .DIN1(n1580), .DIN2(n1515) );
nnd2s1 U1952 ( .Q(n1592), .DIN1(g420), .DIN2(n1581) );
nnd3s1 U1953 ( .Q(n1590), .DIN1(n1613), .DIN2(n1614), .DIN3(g7509) );
nnd2s1 U1954 ( .Q(n1614), .DIN1(g5154), .DIN2(n1585) );
nnd2s1 U1955 ( .Q(n1613), .DIN1(g173), .DIN2(n1588) );
nnd3s1 U1956 ( .Q(n1589), .DIN1(n1615), .DIN2(n1616), .DIN3(n1617) );
nnd2s1 U1957 ( .Q(n1617), .DIN1(g626), .DIN2(n1587) );
nnd2s1 U1958 ( .Q(n1616), .DIN1(g258), .DIN2(n1553) );
nnd2s1 U1959 ( .Q(n1615), .DIN1(g602), .DIN2(n1586) );
or2s1 U1960 ( .Q(g9288), .DIN1(n1388), .DIN2(g9374) );
or3s1 U1961 ( .Q(g9374), .DIN1(n1618), .DIN2(n1619), .DIN3(n1620) );
nnd4s1 U1962 ( .Q(n1620), .DIN1(n1621), .DIN2(n1622), .DIN3(n1623), .DIN4(n1624) );
and3s1 U1963 ( .Q(n1624), .DIN1(n1625), .DIN2(n1626), .DIN3(n1627) );
nnd2s1 U1964 ( .Q(n1627), .DIN1(g184), .DIN2(n1599) );
nnd2s1 U1965 ( .Q(n1626), .DIN1(g616), .DIN2(n1554) );
nnd2s1 U1966 ( .Q(n1625), .DIN1(g342), .DIN2(n1555) );
nnd2s1 U1967 ( .Q(n1623), .DIN1(g588), .DIN2(n1556) );
nnd2s1 U1968 ( .Q(n1622), .DIN1(n1557), .DIN2(n1628) );
nnd4s1 U1969 ( .Q(n1628), .DIN1(n1629), .DIN2(n1630), .DIN3(n1631), .DIN4(n1632) );
nor2s1 U1970 ( .Q(n1632), .DIN1(n1633), .DIN2(n1634) );
and2s1 U1971 ( .Q(n1634), .DIN1(n1565), .DIN2(g769) );
nor2s1 U1972 ( .Q(n1633), .DIN1(n1635), .DIN2(n1425) );
nnd2s1 U1973 ( .Q(n1631), .DIN1(g837), .DIN2(n1567) );
nnd2s1 U1974 ( .Q(n1630), .DIN1(n1568), .DIN2(n1636) );
nnd4s1 U1975 ( .Q(n1636), .DIN1(n1637), .DIN2(n1571), .DIN3(n1638), .DIN4(n1639) );
nor2s1 U1976 ( .Q(n1639), .DIN1(n1640), .DIN2(n1641) );
and2s1 U1977 ( .Q(n1641), .DIN1(n1576), .DIN2(g634) );
and2s1 U1978 ( .Q(n1640), .DIN1(n1577), .DIN2(g665) );
nnd2s1 U1979 ( .Q(n1638), .DIN1(g504), .DIN2(n1578) );
nnd2s1 U1980 ( .Q(n1637), .DIN1(g754), .DIN2(n1579) );
nnd2s1 U1981 ( .Q(n1629), .DIN1(n1580), .DIN2(n1497) );
nnd2s1 U1982 ( .Q(n1621), .DIN1(g423), .DIN2(n1581) );
nnd3s1 U1983 ( .Q(n1619), .DIN1(n1642), .DIN2(n1643), .DIN3(g7509) );
nnd2s1 U1984 ( .Q(n1643), .DIN1(g5155), .DIN2(n1585) );
nnd2s1 U1985 ( .Q(n1642), .DIN1(g150), .DIN2(n1588) );
nnd3s1 U1986 ( .Q(n1618), .DIN1(n1644), .DIN2(n1645), .DIN3(n1646) );
nnd2s1 U1987 ( .Q(n1646), .DIN1(g627), .DIN2(n1587) );
nnd2s1 U1988 ( .Q(n1645), .DIN1(g261), .DIN2(n1553) );
nnd2s1 U1989 ( .Q(n1644), .DIN1(g603), .DIN2(n1586) );
or2s1 U1990 ( .Q(g9285), .DIN1(n1388), .DIN2(g9373) );
or4s1 U1991 ( .Q(g9373), .DIN1(n1647), .DIN2(n1648), .DIN3(n1649), .DIN4(n1650) );
nnd4s1 U1992 ( .Q(n1650), .DIN1(n1651), .DIN2(n1652), .DIN3(n1653), .DIN4(n1654) );
nnd2s1 U1993 ( .Q(n1654), .DIN1(n1557), .DIN2(n1655) );
nnd4s1 U1994 ( .Q(n1655), .DIN1(n1656), .DIN2(n1657), .DIN3(n1658), .DIN4(n1659) );
nnd2s1 U1995 ( .Q(n1659), .DIN1(g840), .DIN2(n1567) );
nor2s1 U1996 ( .Q(n1658), .DIN1(n1660), .DIN2(n1661) );
and2s1 U1997 ( .Q(n1661), .DIN1(n1516), .DIN2(n1580) );
nor2s1 U1998 ( .Q(n1660), .DIN1(n1662), .DIN2(n1663) );
nor2s1 U1999 ( .Q(n1662), .DIN1(n1664), .DIN2(n1665) );
nnd4s1 U2000 ( .Q(n1665), .DIN1(n1666), .DIN2(n1667), .DIN3(n1668), .DIN4(n1669) );
nnd2s1 U2001 ( .Q(n1669), .DIN1(g730), .DIN2(n1670) );
nnd2s1 U2002 ( .Q(n1668), .DIN1(g669), .DIN2(n1577) );
nnd2s1 U2003 ( .Q(n1667), .DIN1(g723), .DIN2(n1671) );
nnd2s1 U2004 ( .Q(n1666), .DIN1(g635), .DIN2(n1576) );
nnd4s1 U2005 ( .Q(n1664), .DIN1(n1672), .DIN2(n1673), .DIN3(n1674), .DIN4(n1571) );
nnd2s1 U2006 ( .Q(n1674), .DIN1(g752), .DIN2(n1579) );
nnd2s1 U2007 ( .Q(n1673), .DIN1(g507), .DIN2(n1578) );
nnd2s1 U2008 ( .Q(n1672), .DIN1(g459), .DIN2(n1675) );
nnd2s1 U2009 ( .Q(n1657), .DIN1(g762), .DIN2(n1566) );
nnd2s1 U2010 ( .Q(n1656), .DIN1(g770), .DIN2(n1565) );
nnd2s1 U2011 ( .Q(n1653), .DIN1(g216), .DIN2(n1676) );
nnd2s1 U2012 ( .Q(n1652), .DIN1(g378), .DIN2(n1677) );
nnd2s1 U2013 ( .Q(n1651), .DIN1(g591), .DIN2(n1556) );
nnd4s1 U2014 ( .Q(n1649), .DIN1(n1678), .DIN2(n1679), .DIN3(n1680), .DIN4(n1681) );
nnd2s1 U2015 ( .Q(n1681), .DIN1(g5156), .DIN2(n1585) );
nor2s1 U2016 ( .Q(n1680), .DIN1(n1682), .DIN2(n1683) );
nor2s1 U2017 ( .Q(n1683), .DIN1(n1684), .DIN2(DFF_270net495) );
and2s1 U2018 ( .Q(n1682), .DIN1(n1587), .DIN2(g628) );
nnd2s1 U2019 ( .Q(n1679), .DIN1(g297), .DIN2(n1685) );
nnd2s1 U2020 ( .Q(n1678), .DIN1(g174), .DIN2(n1588) );
nnd4s1 U2021 ( .Q(n1648), .DIN1(g7509), .DIN2(n1686), .DIN3(n1687), .DIN4(n1688) );
nnd2s1 U2022 ( .Q(n1688), .DIN1(g345), .DIN2(n1555) );
nnd2s1 U2023 ( .Q(n1687), .DIN1(g179), .DIN2(n1599) );
nnd2s1 U2024 ( .Q(n1686), .DIN1(g264), .DIN2(n1553) );
nnd4s1 U2025 ( .Q(n1647), .DIN1(n1689), .DIN2(n1690), .DIN3(n1691), .DIN4(n1692) );
nor2s1 U2026 ( .Q(n1692), .DIN1(n1693), .DIN2(n1694) );
and2s1 U2027 ( .Q(n1694), .DIN1(n1581), .DIN2(g426) );
and2s1 U2028 ( .Q(n1693), .DIN1(n1695), .DIN2(g596) );
nnd2s1 U2029 ( .Q(n1691), .DIN1(g604), .DIN2(n1586) );
nnd2s1 U2030 ( .Q(n1690), .DIN1(g617), .DIN2(n1554) );
nnd2s1 U2031 ( .Q(n1689), .DIN1(g609), .DIN2(n1696) );
or2s1 U2032 ( .Q(g9282), .DIN1(n1388), .DIN2(g9372) );
or4s1 U2033 ( .Q(g9372), .DIN1(n1697), .DIN2(n1698), .DIN3(n1699), .DIN4(n1700) );
nnd4s1 U2034 ( .Q(n1700), .DIN1(n1701), .DIN2(n1702), .DIN3(n1703), .DIN4(n1704) );
nnd2s1 U2035 ( .Q(n1704), .DIN1(n1557), .DIN2(n1705) );
nnd4s1 U2036 ( .Q(n1705), .DIN1(n1706), .DIN2(n1707), .DIN3(n1708), .DIN4(n1709) );
nnd2s1 U2037 ( .Q(n1709), .DIN1(g843), .DIN2(n1567) );
nor2s1 U2038 ( .Q(n1708), .DIN1(n1710), .DIN2(n1711) );
and2s1 U2039 ( .Q(n1711), .DIN1(n1498), .DIN2(n1580) );
nor2s1 U2040 ( .Q(n1710), .DIN1(n1712), .DIN2(n1663) );
nor2s1 U2041 ( .Q(n1712), .DIN1(n1713), .DIN2(n1714) );
nnd4s1 U2042 ( .Q(n1714), .DIN1(n1715), .DIN2(n1716), .DIN3(n1717), .DIN4(n1718) );
nnd2s1 U2043 ( .Q(n1718), .DIN1(g734), .DIN2(n1670) );
nnd2s1 U2044 ( .Q(n1717), .DIN1(g673), .DIN2(n1577) );
nnd2s1 U2045 ( .Q(n1716), .DIN1(g722), .DIN2(n1671) );
nnd2s1 U2046 ( .Q(n1715), .DIN1(g645), .DIN2(n1576) );
nnd4s1 U2047 ( .Q(n1713), .DIN1(n1719), .DIN2(n1720), .DIN3(n1721), .DIN4(n1571) );
nnd2s1 U2048 ( .Q(n1721), .DIN1(g753), .DIN2(n1579) );
nnd2s1 U2049 ( .Q(n1720), .DIN1(g510), .DIN2(n1578) );
nnd2s1 U2050 ( .Q(n1719), .DIN1(g462), .DIN2(n1675) );
nnd2s1 U2051 ( .Q(n1707), .DIN1(g763), .DIN2(n1566) );
nnd2s1 U2052 ( .Q(n1706), .DIN1(g771), .DIN2(n1565) );
nnd2s1 U2053 ( .Q(n1703), .DIN1(g219), .DIN2(n1676) );
nnd2s1 U2054 ( .Q(n1702), .DIN1(g381), .DIN2(n1677) );
nnd2s1 U2055 ( .Q(n1701), .DIN1(g573), .DIN2(n1556) );
nnd4s1 U2056 ( .Q(n1699), .DIN1(n1722), .DIN2(n1723), .DIN3(n1724), .DIN4(n1725) );
nnd2s1 U2057 ( .Q(n1725), .DIN1(g5149), .DIN2(n1585) );
nor2s1 U2058 ( .Q(n1724), .DIN1(n1726), .DIN2(n1727) );
nor2s1 U2059 ( .Q(n1727), .DIN1(n1684), .DIN2(DFF_404net629) );
and2s1 U2060 ( .Q(n1726), .DIN1(n1587), .DIN2(g629) );
nnd2s1 U2061 ( .Q(n1723), .DIN1(g300), .DIN2(n1685) );
nnd2s1 U2062 ( .Q(n1722), .DIN1(g154), .DIN2(n1588) );
nnd4s1 U2063 ( .Q(n1698), .DIN1(g7509), .DIN2(n1728), .DIN3(n1729), .DIN4(n1730) );
nnd2s1 U2064 ( .Q(n1730), .DIN1(g348), .DIN2(n1555) );
nnd2s1 U2065 ( .Q(n1729), .DIN1(g180), .DIN2(n1599) );
nnd2s1 U2066 ( .Q(n1728), .DIN1(g267), .DIN2(n1553) );
nnd4s1 U2067 ( .Q(n1697), .DIN1(n1731), .DIN2(n1732), .DIN3(n1733), .DIN4(n1734) );
nor2s1 U2068 ( .Q(n1734), .DIN1(n1735), .DIN2(n1736) );
and2s1 U2069 ( .Q(n1736), .DIN1(n1581), .DIN2(g429) );
and2s1 U2070 ( .Q(n1735), .DIN1(n1695), .DIN2(g597) );
nnd2s1 U2071 ( .Q(n1733), .DIN1(g605), .DIN2(n1586) );
nnd2s1 U2072 ( .Q(n1732), .DIN1(g618), .DIN2(n1554) );
nnd2s1 U2073 ( .Q(n1731), .DIN1(g610), .DIN2(n1696) );
nnd2s1 U2074 ( .Q(g9267), .DIN1(g62), .DIN2(n1537) );
nor4s1 U2075 ( .Q(n1537), .DIN1(n1737), .DIN2(n1738), .DIN3(n1739), .DIN4(n1740) );
nnd4s1 U2076 ( .Q(n1740), .DIN1(n1741), .DIN2(n1742), .DIN3(n1743), .DIN4(n1744) );
nnd2s1 U2077 ( .Q(n1744), .DIN1(g181), .DIN2(n1599) );
nor2s1 U2078 ( .Q(n1743), .DIN1(n1745), .DIN2(n1746) );
and2s1 U2079 ( .Q(n1746), .DIN1(n1555), .DIN2(g351) );
and2s1 U2080 ( .Q(n1745), .DIN1(n1696), .DIN2(g611) );
nnd2s1 U2081 ( .Q(n1742), .DIN1(g270), .DIN2(n1553) );
nnd2s1 U2082 ( .Q(n1741), .DIN1(g606), .DIN2(n1586) );
nnd4s1 U2083 ( .Q(n1739), .DIN1(n1747), .DIN2(n1748), .DIN3(n1749), .DIN4(n1750) );
nor2s1 U2084 ( .Q(n1750), .DIN1(n1751), .DIN2(n1752) );
and2s1 U2085 ( .Q(n1752), .DIN1(n1554), .DIN2(g619) );
and2s1 U2086 ( .Q(n1751), .DIN1(n1556), .DIN2(g547) );
nnd2s1 U2087 ( .Q(n1749), .DIN1(g432), .DIN2(n1581) );
nnd2s1 U2088 ( .Q(n1748), .DIN1(g622), .DIN2(n1753) );
nnd2s1 U2089 ( .Q(n1747), .DIN1(n1557), .DIN2(n1754) );
nnd4s1 U2090 ( .Q(n1754), .DIN1(n1755), .DIN2(n1756), .DIN3(n1757), .DIN4(n1758) );
and3s1 U2091 ( .Q(n1758), .DIN1(n1759), .DIN2(n1760), .DIN3(n1761) );
nnd2s1 U2092 ( .Q(n1761), .DIN1(g772), .DIN2(n1565) );
nnd2s1 U2093 ( .Q(n1760), .DIN1(g846), .DIN2(n1567) );
nnd2s1 U2094 ( .Q(n1759), .DIN1(g764), .DIN2(n1566) );
nnd2s1 U2095 ( .Q(n1757), .DIN1(n1580), .DIN2(n1519) );
nnd2s1 U2096 ( .Q(n1756), .DIN1(g863), .DIN2(n1762) );
or2s1 U2097 ( .Q(n1755), .DIN1(n1763), .DIN2(n1663) );
nor2s1 U2098 ( .Q(n1763), .DIN1(n1764), .DIN2(n1765) );
nnd4s1 U2099 ( .Q(n1765), .DIN1(n1766), .DIN2(n1767), .DIN3(n1768), .DIN4(n1769) );
nnd2s1 U2100 ( .Q(n1769), .DIN1(g718), .DIN2(n1670) );
nnd2s1 U2101 ( .Q(n1768), .DIN1(g677), .DIN2(n1577) );
nnd2s1 U2102 ( .Q(n1767), .DIN1(g702), .DIN2(n1671) );
nnd2s1 U2103 ( .Q(n1766), .DIN1(g652), .DIN2(n1576) );
nnd4s1 U2104 ( .Q(n1764), .DIN1(n1770), .DIN2(n1771), .DIN3(n1772), .DIN4(n1571) );
nnd2s1 U2105 ( .Q(n1772), .DIN1(g756), .DIN2(n1579) );
nnd2s1 U2106 ( .Q(n1771), .DIN1(g513), .DIN2(n1578) );
nnd2s1 U2107 ( .Q(n1770), .DIN1(g465), .DIN2(n1675) );
nnd4s1 U2108 ( .Q(n1738), .DIN1(g7509), .DIN2(n1773), .DIN3(n1774), .DIN4(n1775) );
nnd2s1 U2109 ( .Q(n1775), .DIN1(g222), .DIN2(n1676) );
nnd2s1 U2110 ( .Q(n1774), .DIN1(g384), .DIN2(n1510) );
nnd2s1 U2111 ( .Q(n1773), .DIN1(n1588), .DIN2(g158) );
nnd4s1 U2112 ( .Q(n1737), .DIN1(n1776), .DIN2(n1777), .DIN3(n1778), .DIN4(n1779) );
nnd2s1 U2113 ( .Q(n1779), .DIN1(g5157), .DIN2(n1780) );
nor2s1 U2114 ( .Q(n1778), .DIN1(n1781), .DIN2(n1782) );
and2s1 U2115 ( .Q(n1782), .DIN1(n1587), .DIN2(g630) );
and2s1 U2116 ( .Q(n1781), .DIN1(n1695), .DIN2(g598) );
nnd2s1 U2117 ( .Q(n1777), .DIN1(g5150), .DIN2(n1585) );
nnd2s1 U2118 ( .Q(n1776), .DIN1(g303), .DIN2(n1685) );
or2s1 U2119 ( .Q(g9264), .DIN1(n1388), .DIN2(g9360) );
or4s1 U2120 ( .Q(g9360), .DIN1(n1783), .DIN2(n1784), .DIN3(n1785), .DIN4(n1786) );
nnd4s1 U2121 ( .Q(n1786), .DIN1(n1787), .DIN2(n1788), .DIN3(n1789), .DIN4(n1790) );
nor2s1 U2122 ( .Q(n1790), .DIN1(n1791), .DIN2(n1792) );
and2s1 U2123 ( .Q(n1792), .DIN1(n1554), .DIN2(g620) );
and2s1 U2124 ( .Q(n1791), .DIN1(n1556), .DIN2(g550) );
nnd2s1 U2125 ( .Q(n1789), .DIN1(g387), .DIN2(n1510) );
nnd2s1 U2126 ( .Q(n1788), .DIN1(n1557), .DIN2(n1793) );
nnd4s1 U2127 ( .Q(n1793), .DIN1(n1794), .DIN2(n1795), .DIN3(n1796), .DIN4(n1797) );
and3s1 U2128 ( .Q(n1797), .DIN1(n1798), .DIN2(n1799), .DIN3(n1800) );
nnd2s1 U2129 ( .Q(n1800), .DIN1(g773), .DIN2(n1565) );
nnd2s1 U2130 ( .Q(n1799), .DIN1(g849), .DIN2(n1567) );
nnd2s1 U2131 ( .Q(n1798), .DIN1(g765), .DIN2(n1566) );
nnd2s1 U2132 ( .Q(n1796), .DIN1(n1580), .DIN2(n1500) );
nnd2s1 U2133 ( .Q(n1795), .DIN1(g859), .DIN2(n1762) );
nnd2s1 U2134 ( .Q(n1794), .DIN1(n1568), .DIN2(n1801) );
or4s1 U2135 ( .Q(n1801), .DIN1(n1802), .DIN2(n1803), .DIN3(n1804), .DIN4(n1805) );
nnd4s1 U2136 ( .Q(n1805), .DIN1(n1806), .DIN2(n1807), .DIN3(n1808), .DIN4(n1809) );
nnd2s1 U2137 ( .Q(n1809), .DIN1(g714), .DIN2(n1670) );
nnd2s1 U2138 ( .Q(n1808), .DIN1(g681), .DIN2(n1577) );
nnd2s1 U2139 ( .Q(n1807), .DIN1(g698), .DIN2(n1671) );
nnd2s1 U2140 ( .Q(n1806), .DIN1(g647), .DIN2(n1576) );
nnd3s1 U2141 ( .Q(n1804), .DIN1(n1810), .DIN2(n1571), .DIN3(n1811) );
nnd2s1 U2142 ( .Q(n1811), .DIN1(g524), .DIN2(n1578) );
nnd2s1 U2143 ( .Q(n1810), .DIN1(g757), .DIN2(n1579) );
nor2s1 U2144 ( .Q(n1803), .DIN1(n1812), .DIN2(n1434) );
and2s1 U2145 ( .Q(n1802), .DIN1(n1675), .DIN2(g468) );
nnd2s1 U2146 ( .Q(n1787), .DIN1(g225), .DIN2(n1676) );
nnd4s1 U2147 ( .Q(n1785), .DIN1(n1813), .DIN2(n1814), .DIN3(n1815), .DIN4(n1816) );
nnd2s1 U2148 ( .Q(n1816), .DIN1(g5147), .DIN2(n1780) );
nor2s1 U2149 ( .Q(n1815), .DIN1(n1817), .DIN2(n1818) );
and2s1 U2150 ( .Q(n1818), .DIN1(n1587), .DIN2(g631) );
and2s1 U2151 ( .Q(n1817), .DIN1(n1753), .DIN2(g623) );
nnd2s1 U2152 ( .Q(n1814), .DIN1(g5151), .DIN2(n1585) );
nnd2s1 U2153 ( .Q(n1813), .DIN1(g306), .DIN2(n1685) );
nnd4s1 U2154 ( .Q(n1784), .DIN1(g7509), .DIN2(n1819), .DIN3(n1820), .DIN4(n1821) );
nnd2s1 U2155 ( .Q(n1821), .DIN1(g182), .DIN2(n1599) );
nnd2s1 U2156 ( .Q(n1820), .DIN1(g281), .DIN2(n1553) );
nnd2s1 U2157 ( .Q(n1819), .DIN1(g162), .DIN2(n1588) );
nnd4s1 U2158 ( .Q(n1783), .DIN1(n1822), .DIN2(n1823), .DIN3(n1824), .DIN4(n1825) );
nor2s1 U2159 ( .Q(n1825), .DIN1(n1826), .DIN2(n1827) );
and2s1 U2160 ( .Q(n1827), .DIN1(n1555), .DIN2(g362) );
and2s1 U2161 ( .Q(n1826), .DIN1(n1581), .DIN2(g443) );
nnd2s1 U2162 ( .Q(n1824), .DIN1(g599), .DIN2(n1695) );
nnd2s1 U2163 ( .Q(n1823), .DIN1(g612), .DIN2(n1696) );
nnd2s1 U2164 ( .Q(n1822), .DIN1(g607), .DIN2(n1586) );
or2s1 U2165 ( .Q(g9261), .DIN1(n1388), .DIN2(g9362) );
or4s1 U2166 ( .Q(g9362), .DIN1(n1828), .DIN2(n1829), .DIN3(n1830), .DIN4(n1831) );
nnd4s1 U2167 ( .Q(n1831), .DIN1(n1832), .DIN2(n1833), .DIN3(n1834), .DIN4(n1835) );
nor2s1 U2168 ( .Q(n1835), .DIN1(n1836), .DIN2(n1837) );
and2s1 U2169 ( .Q(n1837), .DIN1(n1554), .DIN2(g621) );
and2s1 U2170 ( .Q(n1836), .DIN1(n1556), .DIN2(g553) );
and2s1 U2171 ( .Q(n1556), .DIN1(n1838), .DIN2(n1839) );
nnd2s1 U2172 ( .Q(n1834), .DIN1(g390), .DIN2(n1677) );
nnd2s1 U2173 ( .Q(n1833), .DIN1(n1557), .DIN2(n1840) );
nnd4s1 U2174 ( .Q(n1840), .DIN1(n1841), .DIN2(n1842), .DIN3(n1843), .DIN4(n1844) );
and4s1 U2175 ( .Q(n1844), .DIN1(n1845), .DIN2(n1846), .DIN3(n1847), .DIN4(n1848) );
nnd3s1 U2176 ( .Q(n1848), .DIN1(n1849), .DIN2(n1850), .DIN3(g758) );
nnd2s1 U2177 ( .Q(n1847), .DIN1(g855), .DIN2(n1762) );
nnd2s1 U2178 ( .Q(n1846), .DIN1(n1580), .DIN2(n1521) );
nor2s1 U2179 ( .Q(n1580), .DIN1(n1851), .DIN2(g74) );
nnd2s1 U2180 ( .Q(n1845), .DIN1(g852), .DIN2(n1567) );
and2s1 U2181 ( .Q(n1567), .DIN1(n1852), .DIN2(n1839) );
nnd2s1 U2182 ( .Q(n1843), .DIN1(g774), .DIN2(n1565) );
and2s1 U2183 ( .Q(n1565), .DIN1(n1853), .DIN2(n1854) );
nnd2s1 U2184 ( .Q(n1842), .DIN1(n1568), .DIN2(n1855) );
or4s1 U2185 ( .Q(n1855), .DIN1(n1856), .DIN2(n1857), .DIN3(n1858), .DIN4(n1859) );
nnd4s1 U2186 ( .Q(n1859), .DIN1(n1860), .DIN2(n1861), .DIN3(n1862), .DIN4(n1863) );
nnd2s1 U2187 ( .Q(n1863), .DIN1(g710), .DIN2(n1670) );
hi1s1 U2188 ( .Q(n1670), .DIN(n1864) );
nnd2s1 U2189 ( .Q(n1862), .DIN1(g685), .DIN2(n1577) );
hi1s1 U2190 ( .Q(n1577), .DIN(n1865) );
nnd2s1 U2191 ( .Q(n1861), .DIN1(g694), .DIN2(n1671) );
nnd2s1 U2192 ( .Q(n1860), .DIN1(g648), .DIN2(n1576) );
hi1s1 U2193 ( .Q(n1576), .DIN(n1866) );
nnd3s1 U2194 ( .Q(n1858), .DIN1(n1867), .DIN2(n1571), .DIN3(n1868) );
nnd2s1 U2195 ( .Q(n1868), .DIN1(g527), .DIN2(n1578) );
hi1s1 U2196 ( .Q(n1578), .DIN(n1851) );
or2s1 U2197 ( .Q(n1571), .DIN1(n1869), .DIN2(n1870) );
nnd4s1 U2198 ( .Q(n1870), .DIN1(n1871), .DIN2(n1812), .DIN3(n1864), .DIN4(n1872) );
nnd2s1 U2199 ( .Q(n1871), .DIN1(n1873), .DIN2(n1874) );
nnd4s1 U2200 ( .Q(n1869), .DIN1(n1875), .DIN2(n1865), .DIN3(n1866), .DIN4(n1851) );
nnd2s1 U2201 ( .Q(n1851), .DIN1(n1852), .DIN2(n1854) );
nnd2s1 U2202 ( .Q(n1867), .DIN1(g49), .DIN2(n1579) );
hi1s1 U2203 ( .Q(n1579), .DIN(n1875) );
nnd4s1 U2204 ( .Q(n1875), .DIN1(n1876), .DIN2(n1849), .DIN3(g52), .DIN4(n1877) );
and2s1 U2205 ( .Q(n1877), .DIN1(g83), .DIN2(g86) );
nor2s1 U2206 ( .Q(n1857), .DIN1(n1812), .DIN2(n1435) );
and2s1 U2207 ( .Q(n1856), .DIN1(n1675), .DIN2(g471) );
hi1s1 U2208 ( .Q(n1568), .DIN(n1663) );
nnd3s1 U2209 ( .Q(n1663), .DIN1(n1878), .DIN2(n1879), .DIN3(n1880) );
nnd2s1 U2210 ( .Q(n1880), .DIN1(n1852), .DIN2(n1391) );
nnd2s1 U2211 ( .Q(n1841), .DIN1(g766), .DIN2(n1566) );
hi1s1 U2212 ( .Q(n1566), .DIN(n1635) );
nnd2s1 U2213 ( .Q(n1635), .DIN1(n1839), .DIN2(n1850) );
nor4s1 U2214 ( .Q(n1557), .DIN1(n1599), .DIN2(n1554), .DIN3(n1881), .DIN4(n1882) );
nnd4s1 U2215 ( .Q(n1882), .DIN1(n1684), .DIN2(n1883), .DIN3(n1884), .DIN4(n1885) );
nor2s1 U2216 ( .Q(n1885), .DIN1(n1886), .DIN2(n1696) );
nnd3s1 U2217 ( .Q(n1881), .DIN1(n1887), .DIN2(n1888), .DIN3(n1889) );
and2s1 U2218 ( .Q(n1554), .DIN1(n1890), .DIN2(n1839) );
nnd2s1 U2219 ( .Q(n1832), .DIN1(g228), .DIN2(n1676) );
nnd4s1 U2220 ( .Q(n1830), .DIN1(n1891), .DIN2(n1892), .DIN3(n1893), .DIN4(n1894) );
nnd2s1 U2221 ( .Q(n1894), .DIN1(g5148), .DIN2(n1780) );
hi1s1 U2222 ( .Q(n1780), .DIN(n1684) );
nnd2s1 U2223 ( .Q(n1684), .DIN1(n1895), .DIN2(n1849) );
nor2s1 U2224 ( .Q(n1893), .DIN1(n1896), .DIN2(n1897) );
and2s1 U2225 ( .Q(n1897), .DIN1(n1587), .DIN2(g632) );
and2s1 U2226 ( .Q(n1587), .DIN1(n1854), .DIN2(n1850) );
and2s1 U2227 ( .Q(n1896), .DIN1(n1753), .DIN2(g624) );
and2s1 U2228 ( .Q(n1753), .DIN1(n1874), .DIN2(n1850) );
hi1s1 U2229 ( .Q(n1850), .DIN(n1879) );
nnd4s1 U2230 ( .Q(n1879), .DIN1(g80), .DIN2(n1898), .DIN3(n1391), .DIN4(n1409) );
nnd2s1 U2231 ( .Q(n1892), .DIN1(g5152), .DIN2(n1585) );
hi1s1 U2232 ( .Q(n1585), .DIN(n1887) );
nnd2s1 U2233 ( .Q(n1887), .DIN1(n1839), .DIN2(n1895) );
nnd2s1 U2234 ( .Q(n1891), .DIN1(g309), .DIN2(n1685) );
nnd4s1 U2235 ( .Q(n1829), .DIN1(g7509), .DIN2(n1899), .DIN3(n1900), .DIN4(n1901) );
nnd2s1 U2236 ( .Q(n1901), .DIN1(g185), .DIN2(n1599) );
and2s1 U2237 ( .Q(n1599), .DIN1(n1895), .DIN2(n1854) );
nnd2s1 U2238 ( .Q(n1900), .DIN1(g284), .DIN2(n1553) );
and2s1 U2239 ( .Q(n1553), .DIN1(n1886), .DIN2(n1854) );
nnd2s1 U2240 ( .Q(n1899), .DIN1(g2654), .DIN2(n1588) );
hi1s1 U2241 ( .Q(n1588), .DIN(n1888) );
nnd4s1 U2242 ( .Q(n1828), .DIN1(n1902), .DIN2(n1903), .DIN3(n1904), .DIN4(n1905) );
nor2s1 U2243 ( .Q(n1905), .DIN1(n1906), .DIN2(n1907) );
and2s1 U2244 ( .Q(n1907), .DIN1(n1555), .DIN2(g365) );
and2s1 U2245 ( .Q(n1555), .DIN1(n1886), .DIN2(n1839) );
and2s1 U2246 ( .Q(n1906), .DIN1(n1581), .DIN2(g446) );
and2s1 U2247 ( .Q(n1581), .DIN1(n1838), .DIN2(n1854) );
nnd2s1 U2248 ( .Q(n1904), .DIN1(g600), .DIN2(n1695) );
hi1s1 U2249 ( .Q(n1695), .DIN(n1884) );
nnd2s1 U2250 ( .Q(n1884), .DIN1(n1890), .DIN2(n1874) );
nnd2s1 U2251 ( .Q(n1903), .DIN1(g613), .DIN2(n1696) );
and2s1 U2252 ( .Q(n1696), .DIN1(n1890), .DIN2(n1849) );
nnd2s1 U2253 ( .Q(n1902), .DIN1(g608), .DIN2(n1586) );
hi1s1 U2254 ( .Q(n1586), .DIN(n1889) );
nnd2s1 U2255 ( .Q(n1889), .DIN1(n1890), .DIN2(n1854) );
and3s1 U2256 ( .Q(n1890), .DIN1(g74), .DIN2(n1908), .DIN3(g77) );
nnd2s1 U2257 ( .Q(g9145), .DIN1(n1909), .DIN2(n1910) );
nnd2s1 U2258 ( .Q(n1910), .DIN1(g1069), .DIN2(n1911) );
nnd2s1 U2259 ( .Q(n1909), .DIN1(n1912), .DIN2(g4267) );
nnd2s1 U2260 ( .Q(g9134), .DIN1(n1913), .DIN2(n1914) );
nnd2s1 U2261 ( .Q(n1914), .DIN1(n1911), .DIN2(n1470) );
and3s1 U2262 ( .Q(n1911), .DIN1(n1915), .DIN2(n1916), .DIN3(g1065) );
nnd2s1 U2263 ( .Q(n1913), .DIN1(g1069), .DIN2(n1917) );
nnd2s1 U2264 ( .Q(n1917), .DIN1(n1918), .DIN2(n1919) );
nnd2s1 U2265 ( .Q(n1919), .DIN1(n1920), .DIN2(n1440) );
hi1s1 U2266 ( .Q(n1918), .DIN(n1921) );
nor2s1 U2267 ( .Q(g9133), .DIN1(g2653), .DIN2(n1922) );
nnd2s1 U2268 ( .Q(g9117), .DIN1(n1923), .DIN2(n1924) );
nnd2s1 U2269 ( .Q(n1924), .DIN1(g1065), .DIN2(n1921) );
nnd3s1 U2270 ( .Q(n1923), .DIN1(n1915), .DIN2(n1916), .DIN3(n1440) );
hi1s1 U2271 ( .Q(n1916), .DIN(n1925) );
nnd2s1 U2272 ( .Q(g9116), .DIN1(n1926), .DIN2(n1927) );
nnd2s1 U2273 ( .Q(n1927), .DIN1(g513), .DIN2(n1872) );
nnd2s1 U2274 ( .Q(n1926), .DIN1(g495), .DIN2(n1675) );
nnd2s1 U2275 ( .Q(g9115), .DIN1(n1928), .DIN2(n1929) );
nnd2s1 U2276 ( .Q(n1929), .DIN1(g510), .DIN2(n1872) );
nnd2s1 U2277 ( .Q(n1928), .DIN1(g492), .DIN2(n1675) );
nnd2s1 U2278 ( .Q(g9114), .DIN1(n1930), .DIN2(n1931) );
nnd2s1 U2279 ( .Q(n1931), .DIN1(g507), .DIN2(n1872) );
nnd2s1 U2280 ( .Q(n1930), .DIN1(g489), .DIN2(n1675) );
nnd2s1 U2281 ( .Q(g9113), .DIN1(n1932), .DIN2(n1933) );
nnd2s1 U2282 ( .Q(n1933), .DIN1(g504), .DIN2(n1872) );
nnd2s1 U2283 ( .Q(n1932), .DIN1(g486), .DIN2(n1675) );
nnd2s1 U2284 ( .Q(g9112), .DIN1(n1934), .DIN2(n1935) );
nnd2s1 U2285 ( .Q(n1935), .DIN1(g501), .DIN2(n1872) );
nnd2s1 U2286 ( .Q(n1934), .DIN1(g483), .DIN2(n1675) );
nnd2s1 U2287 ( .Q(g9111), .DIN1(n1936), .DIN2(n1937) );
nnd2s1 U2288 ( .Q(n1937), .DIN1(g498), .DIN2(n1872) );
nnd2s1 U2289 ( .Q(n1936), .DIN1(g480), .DIN2(n1675) );
nnd2s1 U2290 ( .Q(g9110), .DIN1(n1938), .DIN2(n1939) );
nnd2s1 U2291 ( .Q(n1939), .DIN1(g527), .DIN2(n1872) );
nnd2s1 U2292 ( .Q(n1938), .DIN1(g521), .DIN2(n1675) );
nnd2s1 U2293 ( .Q(g9109), .DIN1(n1940), .DIN2(n1941) );
nnd2s1 U2294 ( .Q(n1941), .DIN1(g524), .DIN2(n1872) );
nnd2s1 U2295 ( .Q(n1940), .DIN1(g518), .DIN2(n1675) );
hi1s1 U2296 ( .Q(n1675), .DIN(n1872) );
nnd4s1 U2297 ( .Q(n1872), .DIN1(n1852), .DIN2(g7509), .DIN3(g74), .DIN4(n1874) );
and3s1 U2298 ( .Q(n1852), .DIN1(g80), .DIN2(n1898), .DIN3(g77) );
nnd2s1 U2299 ( .Q(g9108), .DIN1(n1942), .DIN2(n1943) );
nnd2s1 U2300 ( .Q(n1943), .DIN1(g432), .DIN2(n1944) );
nnd2s1 U2301 ( .Q(n1942), .DIN1(g414), .DIN2(n1677) );
nnd2s1 U2302 ( .Q(g9107), .DIN1(n1945), .DIN2(n1946) );
nnd2s1 U2303 ( .Q(n1946), .DIN1(g429), .DIN2(n1944) );
nnd2s1 U2304 ( .Q(n1945), .DIN1(g411), .DIN2(n1677) );
nnd2s1 U2305 ( .Q(g9106), .DIN1(n1947), .DIN2(n1948) );
nnd2s1 U2306 ( .Q(n1948), .DIN1(g426), .DIN2(n1944) );
nnd2s1 U2307 ( .Q(n1947), .DIN1(g408), .DIN2(n1677) );
nnd2s1 U2308 ( .Q(g9105), .DIN1(n1949), .DIN2(n1950) );
nnd2s1 U2309 ( .Q(n1950), .DIN1(g423), .DIN2(n1944) );
nnd2s1 U2310 ( .Q(n1949), .DIN1(g405), .DIN2(n1677) );
nnd2s1 U2311 ( .Q(g9104), .DIN1(n1951), .DIN2(n1952) );
nnd2s1 U2312 ( .Q(n1952), .DIN1(g420), .DIN2(n1944) );
nnd2s1 U2313 ( .Q(n1951), .DIN1(g402), .DIN2(n1677) );
nnd2s1 U2314 ( .Q(g9103), .DIN1(n1953), .DIN2(n1954) );
nnd2s1 U2315 ( .Q(n1954), .DIN1(g417), .DIN2(n1944) );
nnd2s1 U2316 ( .Q(n1953), .DIN1(g399), .DIN2(n1677) );
nnd2s1 U2317 ( .Q(g9102), .DIN1(n1955), .DIN2(n1956) );
nnd2s1 U2318 ( .Q(n1956), .DIN1(g446), .DIN2(n1944) );
nnd2s1 U2319 ( .Q(n1955), .DIN1(g440), .DIN2(n1677) );
nnd2s1 U2320 ( .Q(g9101), .DIN1(n1957), .DIN2(n1958) );
nnd2s1 U2321 ( .Q(n1958), .DIN1(g443), .DIN2(n1944) );
nnd2s1 U2322 ( .Q(n1957), .DIN1(g437), .DIN2(n1677) );
nnd2s1 U2323 ( .Q(g9100), .DIN1(n1959), .DIN2(n1960) );
nnd2s1 U2324 ( .Q(n1960), .DIN1(g351), .DIN2(n1961) );
nnd2s1 U2325 ( .Q(n1959), .DIN1(g333), .DIN2(n1685) );
nnd2s1 U2326 ( .Q(g9099), .DIN1(n1962), .DIN2(n1963) );
nnd2s1 U2327 ( .Q(n1963), .DIN1(g348), .DIN2(n1961) );
nnd2s1 U2328 ( .Q(n1962), .DIN1(g330), .DIN2(n1685) );
nnd2s1 U2329 ( .Q(g9098), .DIN1(n1964), .DIN2(n1965) );
nnd2s1 U2330 ( .Q(n1965), .DIN1(g345), .DIN2(n1961) );
nnd2s1 U2331 ( .Q(n1964), .DIN1(g327), .DIN2(n1685) );
nnd2s1 U2332 ( .Q(g9097), .DIN1(n1966), .DIN2(n1967) );
nnd2s1 U2333 ( .Q(n1967), .DIN1(g342), .DIN2(n1961) );
nnd2s1 U2334 ( .Q(n1966), .DIN1(g324), .DIN2(n1685) );
nnd2s1 U2335 ( .Q(g9096), .DIN1(n1968), .DIN2(n1969) );
nnd2s1 U2336 ( .Q(n1969), .DIN1(g339), .DIN2(n1961) );
nnd2s1 U2337 ( .Q(n1968), .DIN1(g321), .DIN2(n1685) );
nnd2s1 U2338 ( .Q(g9095), .DIN1(n1970), .DIN2(n1971) );
nnd2s1 U2339 ( .Q(n1971), .DIN1(g336), .DIN2(n1961) );
nnd2s1 U2340 ( .Q(n1970), .DIN1(g318), .DIN2(n1685) );
nnd2s1 U2341 ( .Q(g9094), .DIN1(n1972), .DIN2(n1973) );
nnd2s1 U2342 ( .Q(n1973), .DIN1(g365), .DIN2(n1961) );
nnd2s1 U2343 ( .Q(n1972), .DIN1(g359), .DIN2(n1685) );
nnd2s1 U2344 ( .Q(g9093), .DIN1(n1974), .DIN2(n1975) );
nnd2s1 U2345 ( .Q(n1975), .DIN1(g362), .DIN2(n1961) );
nnd2s1 U2346 ( .Q(n1974), .DIN1(g356), .DIN2(n1685) );
hi1s1 U2347 ( .Q(n1685), .DIN(n1961) );
nnd3s1 U2348 ( .Q(n1961), .DIN1(g7509), .DIN2(n1849), .DIN3(n1886) );
nnd2s1 U2349 ( .Q(g9092), .DIN1(n1976), .DIN2(n1977) );
nnd2s1 U2350 ( .Q(n1977), .DIN1(g270), .DIN2(n1978) );
nnd2s1 U2351 ( .Q(n1976), .DIN1(g252), .DIN2(n1676) );
nnd2s1 U2352 ( .Q(g9091), .DIN1(n1979), .DIN2(n1980) );
nnd2s1 U2353 ( .Q(n1980), .DIN1(g267), .DIN2(n1978) );
nnd2s1 U2354 ( .Q(n1979), .DIN1(g249), .DIN2(n1676) );
nnd2s1 U2355 ( .Q(g9090), .DIN1(n1981), .DIN2(n1982) );
nnd2s1 U2356 ( .Q(n1982), .DIN1(g264), .DIN2(n1978) );
nnd2s1 U2357 ( .Q(n1981), .DIN1(g246), .DIN2(n1676) );
nnd2s1 U2358 ( .Q(g9089), .DIN1(n1983), .DIN2(n1984) );
nnd2s1 U2359 ( .Q(n1984), .DIN1(g261), .DIN2(n1978) );
nnd2s1 U2360 ( .Q(n1983), .DIN1(g243), .DIN2(n1676) );
nnd2s1 U2361 ( .Q(g9088), .DIN1(n1985), .DIN2(n1986) );
nnd2s1 U2362 ( .Q(n1986), .DIN1(g258), .DIN2(n1978) );
nnd2s1 U2363 ( .Q(n1985), .DIN1(g240), .DIN2(n1676) );
nnd2s1 U2364 ( .Q(g9087), .DIN1(n1987), .DIN2(n1988) );
nnd2s1 U2365 ( .Q(n1988), .DIN1(g255), .DIN2(n1978) );
nnd2s1 U2366 ( .Q(n1987), .DIN1(g237), .DIN2(n1676) );
nnd2s1 U2367 ( .Q(g9086), .DIN1(n1989), .DIN2(n1990) );
nnd2s1 U2368 ( .Q(n1990), .DIN1(g284), .DIN2(n1978) );
nnd2s1 U2369 ( .Q(n1989), .DIN1(g278), .DIN2(n1676) );
nnd2s1 U2370 ( .Q(g9085), .DIN1(n1991), .DIN2(n1992) );
nnd2s1 U2371 ( .Q(n1992), .DIN1(g281), .DIN2(n1978) );
nnd2s1 U2372 ( .Q(n1991), .DIN1(g275), .DIN2(n1676) );
hi1s1 U2373 ( .Q(n1676), .DIN(n1978) );
nnd3s1 U2374 ( .Q(n1978), .DIN1(g7509), .DIN2(n1874), .DIN3(n1886) );
and3s1 U2375 ( .Q(n1886), .DIN1(n1908), .DIN2(n1409), .DIN3(g74) );
nor2s1 U2376 ( .Q(g9036), .DIN1(n1993), .DIN2(n1994) );
xor2s1 U2377 ( .Q(n1993), .DIN1(g1477), .DIN2(n1995) );
nnd2s1 U2378 ( .Q(n1995), .DIN1(n1996), .DIN2(g1472) );
nnd2s1 U2379 ( .Q(g9035), .DIN1(n1997), .DIN2(n1998) );
nnd4s1 U2380 ( .Q(n1998), .DIN1(n1915), .DIN2(g1057), .DIN3(n1999), .DIN4(n1925) );
nnd2s1 U2381 ( .Q(n1997), .DIN1(g1061), .DIN2(n1921) );
nnd2s1 U2382 ( .Q(n1921), .DIN1(n2000), .DIN2(n2001) );
nnd2s1 U2383 ( .Q(n2001), .DIN1(n1925), .DIN2(n1920) );
nnd3s1 U2384 ( .Q(n1925), .DIN1(g1057), .DIN2(n1999), .DIN3(g1061) );
and2s1 U2385 ( .Q(g9034), .DIN1(n2002), .DIN2(n2003) );
nnd3s1 U2386 ( .Q(n2002), .DIN1(n2004), .DIN2(g6565), .DIN3(n2005) );
hi1s1 U2387 ( .Q(n2005), .DIN(n2006) );
or3s1 U2388 ( .Q(n2004), .DIN1(g1021), .DIN2(g1025), .DIN3(n1433) );
nnd2s1 U2389 ( .Q(g9033), .DIN1(n2007), .DIN2(n2008) );
nnd2s1 U2390 ( .Q(n2008), .DIN1(g573), .DIN2(n1944) );
nnd2s1 U2391 ( .Q(n2007), .DIN1(g560), .DIN2(n1677) );
nnd2s1 U2392 ( .Q(g9032), .DIN1(n2009), .DIN2(n2010) );
nnd2s1 U2393 ( .Q(n2010), .DIN1(g591), .DIN2(n1944) );
nnd2s1 U2394 ( .Q(n2009), .DIN1(g584), .DIN2(n1677) );
nnd2s1 U2395 ( .Q(g9031), .DIN1(n2011), .DIN2(n2012) );
nnd2s1 U2396 ( .Q(n2012), .DIN1(g588), .DIN2(n1944) );
nnd2s1 U2397 ( .Q(n2011), .DIN1(g580), .DIN2(n1677) );
nnd2s1 U2398 ( .Q(g9030), .DIN1(n2013), .DIN2(n2014) );
nnd2s1 U2399 ( .Q(n2014), .DIN1(g570), .DIN2(n1944) );
nnd2s1 U2400 ( .Q(n2013), .DIN1(g567), .DIN2(n1677) );
nnd2s1 U2401 ( .Q(g9029), .DIN1(n2015), .DIN2(n2016) );
nnd2s1 U2402 ( .Q(n2016), .DIN1(g563), .DIN2(n1944) );
nnd2s1 U2403 ( .Q(n2015), .DIN1(g557), .DIN2(n1677) );
nnd2s1 U2404 ( .Q(g9028), .DIN1(n2017), .DIN2(n2018) );
nnd2s1 U2405 ( .Q(n2018), .DIN1(g553), .DIN2(n1944) );
nnd2s1 U2406 ( .Q(n2017), .DIN1(g544), .DIN2(n1677) );
nnd2s1 U2407 ( .Q(g9027), .DIN1(n2019), .DIN2(n2020) );
nnd2s1 U2408 ( .Q(n2020), .DIN1(g550), .DIN2(n1944) );
nnd2s1 U2409 ( .Q(n2019), .DIN1(g540), .DIN2(n1677) );
nnd2s1 U2410 ( .Q(g9026), .DIN1(n2021), .DIN2(n2022) );
nnd2s1 U2411 ( .Q(n2022), .DIN1(g547), .DIN2(n1944) );
nnd2s1 U2412 ( .Q(n2021), .DIN1(g536), .DIN2(n1677) );
hi1s1 U2413 ( .Q(n1677), .DIN(n1944) );
nnd3s1 U2414 ( .Q(n1944), .DIN1(g7509), .DIN2(n1874), .DIN3(n1838) );
hi1s1 U2415 ( .Q(n1838), .DIN(n1883) );
nnd3s1 U2416 ( .Q(n1883), .DIN1(n1908), .DIN2(n1391), .DIN3(g77) );
nor2s1 U2417 ( .Q(g8960), .DIN1(n2023), .DIN2(n1994) );
xor2s1 U2418 ( .Q(n2023), .DIN1(n2024), .DIN2(g1472) );
nnd2s1 U2419 ( .Q(g8959), .DIN1(n2025), .DIN2(n2026) );
nnd2s1 U2420 ( .Q(n2026), .DIN1(g1057), .DIN2(n2027) );
nnd3s1 U2421 ( .Q(n2025), .DIN1(n1915), .DIN2(n1999), .DIN3(n1459) );
hi1s1 U2422 ( .Q(n1999), .DIN(n2028) );
nor2s1 U2423 ( .Q(g8957), .DIN1(n2029), .DIN2(n2030) );
nor2s1 U2424 ( .Q(n2030), .DIN1(g4599), .DIN2(n2006) );
nnd3s1 U2425 ( .Q(n2006), .DIN1(n2031), .DIN2(n2032), .DIN3(n1922) );
nnd4s1 U2426 ( .Q(n2032), .DIN1(g998), .DIN2(n2033), .DIN3(g999), .DIN4(n2034) );
or4s1 U2427 ( .Q(n2031), .DIN1(DFF_160net385), .DIN2(n2035), .DIN3(n2036), .DIN4(n2034) );
or3s1 U2428 ( .Q(n2036), .DIN1(g1016), .DIN2(g1008), .DIN3(I5528) );
hi1s1 U2429 ( .Q(n2029), .DIN(n2037) );
nnd3s1 U2430 ( .Q(n1812), .DIN1(g77), .DIN2(n1854), .DIN3(n1873) );
nnd2s1 U2431 ( .Q(n2039), .DIN1(n1435), .DIN2(n2040) );
nnd4s1 U2432 ( .Q(n2040), .DIN1(g55), .DIN2(n1527), .DIN3(n1529), .DIN4(n2041) );
hi1s1 U2433 ( .Q(n1529), .DIN(g42) );
hi1s1 U2434 ( .Q(n1527), .DIN(g41) );
nor2s1 U2435 ( .Q(g8875), .DIN1(n2042), .DIN2(n1994) );
and2s1 U2436 ( .Q(n2042), .DIN1(n2043), .DIN2(n2044) );
nnd3s1 U2437 ( .Q(n2044), .DIN1(g1462), .DIN2(n2045), .DIN3(n2046) );
nnd2s1 U2438 ( .Q(n2043), .DIN1(g1467), .DIN2(n2024) );
hi1s1 U2439 ( .Q(n2024), .DIN(n1996) );
nor2s1 U2440 ( .Q(n1996), .DIN1(n2045), .DIN2(g4659) );
nnd4s1 U2441 ( .Q(n2045), .DIN1(n2047), .DIN2(g1519), .DIN3(g1467), .DIN4(g1462) );
nor2s1 U2442 ( .Q(g8874), .DIN1(g1097), .DIN2(n2048) );
xor2s1 U2443 ( .Q(n2048), .DIN1(g1142), .DIN2(n2049) );
nnd2s1 U2444 ( .Q(g8873), .DIN1(n2050), .DIN2(n2051) );
nnd3s1 U2445 ( .Q(n2051), .DIN1(n2052), .DIN2(n2028), .DIN3(n1915) );
nnd2s1 U2446 ( .Q(n2050), .DIN1(g1053), .DIN2(n2027) );
nnd2s1 U2447 ( .Q(n2027), .DIN1(n2000), .DIN2(n2053) );
nnd2s1 U2448 ( .Q(n2053), .DIN1(n2028), .DIN2(n1920) );
nnd2s1 U2449 ( .Q(n2028), .DIN1(g1053), .DIN2(n2052) );
hi1s1 U2450 ( .Q(n2052), .DIN(n2054) );
nnd2s1 U2451 ( .Q(g8871), .DIN1(n2055), .DIN2(n2056) );
nnd3s1 U2452 ( .Q(n2056), .DIN1(n2057), .DIN2(n2058), .DIN3(g1025) );
and3s1 U2453 ( .Q(g8870), .DIN1(n2059), .DIN2(n1446), .DIN3(n2057) );
nnd2s1 U2454 ( .Q(n2059), .DIN1(n2058), .DIN2(n2060) );
nnd2s1 U2455 ( .Q(n2060), .DIN1(g1021), .DIN2(g1018) );
nnd2s1 U2456 ( .Q(g8869), .DIN1(n2055), .DIN2(n2061) );
nnd2s1 U2457 ( .Q(n2061), .DIN1(n2057), .DIN2(n1433) );
and3s1 U2458 ( .Q(n2057), .DIN1(n2062), .DIN2(g6851), .DIN3(n2063) );
or2s1 U2459 ( .Q(n2063), .DIN1(n2058), .DIN2(g1025) );
or2s1 U2460 ( .Q(n2058), .DIN1(g1021), .DIN2(g1018) );
nnd3s1 U2461 ( .Q(n2055), .DIN1(n2062), .DIN2(g6851), .DIN3(g1029) );
nnd2s1 U2462 ( .Q(n2062), .DIN1(n1401), .DIN2(g6565) );
and4s1 U2463 ( .Q(g8867), .DIN1(g6310), .DIN2(g6309), .DIN3(n2064), .DIN4(n2065) );
and2s1 U2464 ( .Q(n2065), .DIN1(g7105), .DIN2(g1013) );
and4s1 U2465 ( .Q(g8865), .DIN1(n2064), .DIN2(g998), .DIN3(n2033), .DIN4(n2034) );
and2s1 U2466 ( .Q(g8864), .DIN1(g6851), .DIN2(g7071) );
nor2s1 U2467 ( .Q(g8678), .DIN1(n2066), .DIN2(n1994) );
hi1s1 U2468 ( .Q(n2066), .DIN(n2067) );
xor2s1 U2469 ( .Q(n2067), .DIN1(g1462), .DIN2(n2046) );
nor2s1 U2470 ( .Q(n2046), .DIN1(n2068), .DIN2(n1451) );
nor2s1 U2471 ( .Q(g8676), .DIN1(n2069), .DIN2(n1403) );
xor2s1 U2472 ( .Q(n2069), .DIN1(g1360), .DIN2(n2070) );
nnd2s1 U2473 ( .Q(n2070), .DIN1(g1357), .DIN2(n2071) );
hi1s1 U2474 ( .Q(n2071), .DIN(n2072) );
nor2s1 U2475 ( .Q(g8675), .DIN1(n2073), .DIN2(n1403) );
xor2s1 U2476 ( .Q(n2073), .DIN1(g1357), .DIN2(n2072) );
nnd3s1 U2477 ( .Q(g8674), .DIN1(n2074), .DIN2(n1402), .DIN3(n2075) );
nnd2s1 U2478 ( .Q(n2075), .DIN1(g1126), .DIN2(n2049) );
nnd2s1 U2479 ( .Q(n2049), .DIN1(g1148), .DIN2(n2076) );
nnd3s1 U2480 ( .Q(n2074), .DIN1(g1122), .DIN2(n2077), .DIN3(n2078) );
nnd2s1 U2481 ( .Q(g8673), .DIN1(n2079), .DIN2(n2080) );
nnd4s1 U2482 ( .Q(n2080), .DIN1(n1915), .DIN2(g1045), .DIN3(n2081), .DIN4(n2054) );
nnd2s1 U2483 ( .Q(n2079), .DIN1(g1049), .DIN2(n2082) );
nnd2s1 U2484 ( .Q(n2082), .DIN1(n2000), .DIN2(n2083) );
nnd2s1 U2485 ( .Q(n2083), .DIN1(n2054), .DIN2(n1920) );
nnd3s1 U2486 ( .Q(n2054), .DIN1(g1045), .DIN2(n2081), .DIN3(g1049) );
and2s1 U2487 ( .Q(g8672), .DIN1(g6851), .DIN2(g6745) );
nnd2s1 U2488 ( .Q(g8671), .DIN1(n2084), .DIN2(n2085) );
nnd2s1 U2489 ( .Q(n2085), .DIN1(g954), .DIN2(n2086) );
nnd2s1 U2490 ( .Q(n2084), .DIN1(n2087), .DIN2(n1522) );
nnd2s1 U2491 ( .Q(g8670), .DIN1(n2088), .DIN2(n2089) );
nnd2s1 U2492 ( .Q(n2089), .DIN1(g953), .DIN2(n2086) );
nnd2s1 U2493 ( .Q(n2088), .DIN1(n2087), .DIN2(n1501) );
nnd2s1 U2494 ( .Q(g8669), .DIN1(n2090), .DIN2(n2091) );
nnd2s1 U2495 ( .Q(n2091), .DIN1(g952), .DIN2(n2086) );
nnd2s1 U2496 ( .Q(n2090), .DIN1(n2087), .DIN2(n1518) );
nnd2s1 U2497 ( .Q(g8668), .DIN1(n2092), .DIN2(n2093) );
nnd2s1 U2498 ( .Q(n2093), .DIN1(g951), .DIN2(n2086) );
nnd2s1 U2499 ( .Q(n2092), .DIN1(n2087), .DIN2(n1498) );
nnd2s1 U2500 ( .Q(g8667), .DIN1(n2094), .DIN2(n2095) );
nnd2s1 U2501 ( .Q(n2095), .DIN1(g950), .DIN2(n2086) );
nnd2s1 U2502 ( .Q(n2094), .DIN1(n2087), .DIN2(n1386) );
nnd2s1 U2503 ( .Q(g8666), .DIN1(n2096), .DIN2(n2097) );
nnd2s1 U2504 ( .Q(n2097), .DIN1(g949), .DIN2(n2086) );
nnd2s1 U2505 ( .Q(n2096), .DIN1(n2087), .DIN2(n1497) );
nnd2s1 U2506 ( .Q(g8665), .DIN1(n2098), .DIN2(n2099) );
nnd2s1 U2507 ( .Q(n2099), .DIN1(g948), .DIN2(n2086) );
nnd2s1 U2508 ( .Q(n2098), .DIN1(n2087), .DIN2(n1387) );
nnd2s1 U2509 ( .Q(g8664), .DIN1(n2087), .DIN2(n1511) );
nnd2s1 U2510 ( .Q(g8662), .DIN1(g944), .DIN2(n1471) );
nnd2s1 U2511 ( .Q(g8633), .DIN1(g6310), .DIN2(n2100) );
nnd2s1 U2512 ( .Q(n2100), .DIN1(n2101), .DIN2(n1442) );
and4s1 U2513 ( .Q(g8630), .DIN1(g1013), .DIN2(n2064), .DIN3(g6310), .DIN4(g162) );
nnd2s1 U2514 ( .Q(g8627), .DIN1(g6310), .DIN2(n2102) );
nnd3s1 U2515 ( .Q(n2102), .DIN1(n2103), .DIN2(n1442), .DIN3(n2101) );
nnd2s1 U2516 ( .Q(n2103), .DIN1(n2035), .DIN2(g6565) );
hi1s1 U2517 ( .Q(n2035), .DIN(g6309) );
and4s1 U2518 ( .Q(g8625), .DIN1(n2064), .DIN2(g162), .DIN3(g6851), .DIN4(n2033) );
hi1s1 U2519 ( .Q(n2033), .DIN(g1000) );
and4s1 U2520 ( .Q(n2064), .DIN1(n2101), .DIN2(n2104), .DIN3(n2105), .DIN4(n2003) );
nor2s1 U2521 ( .Q(n2105), .DIN1(g4599), .DIN2(g2653) );
nor2s1 U2522 ( .Q(n2101), .DIN1(g8223), .DIN2(g7104) );
nor2s1 U2523 ( .Q(g8227), .DIN1(n2106), .DIN2(n1994) );
xor2s1 U2524 ( .Q(n2106), .DIN1(n2068), .DIN2(g1519) );
nnd2s1 U2525 ( .Q(g8226), .DIN1(n2107), .DIN2(n2108) );
or2s1 U2526 ( .Q(n2108), .DIN1(n2109), .DIN2(g1911) );
nnd2s1 U2527 ( .Q(n2107), .DIN1(n2110), .DIN2(n2109) );
xor2s1 U2528 ( .Q(n2110), .DIN1(g6223), .DIN2(n2111) );
nnd2s1 U2529 ( .Q(g8225), .DIN1(n2112), .DIN2(n1402) );
xor2s1 U2530 ( .Q(n2112), .DIN1(g1122), .DIN2(n2113) );
nnd2s1 U2531 ( .Q(g8224), .DIN1(n2114), .DIN2(n2115) );
nnd2s1 U2532 ( .Q(n2115), .DIN1(g1045), .DIN2(n2116) );
nnd3s1 U2533 ( .Q(n2114), .DIN1(n1915), .DIN2(n2081), .DIN3(n1460) );
hi1s1 U2534 ( .Q(n2081), .DIN(n2117) );
hi1s1 U2535 ( .Q(g8223), .DIN(n1922) );
nnd3s1 U2536 ( .Q(n1922), .DIN1(n2104), .DIN2(g6851), .DIN3(g973) );
or2s1 U2537 ( .Q(n2119), .DIN1(g866), .DIN2(g863) );
and2s1 U2538 ( .Q(n1762), .DIN1(n1853), .DIN2(n1839) );
hi1s1 U2539 ( .Q(n1853), .DIN(n1878) );
nnd2s1 U2540 ( .Q(n1878), .DIN1(n1876), .DIN2(n1898) );
and3s1 U2541 ( .Q(n1876), .DIN1(g80), .DIN2(n1409), .DIN3(g74) );
nor2s1 U2542 ( .Q(g7775), .DIN1(n2122), .DIN2(n1994) );
and2s1 U2543 ( .Q(n2122), .DIN1(n2123), .DIN2(n2124) );
nnd3s1 U2544 ( .Q(n2124), .DIN1(g1509), .DIN2(n2125), .DIN3(n2126) );
nnd2s1 U2545 ( .Q(n2123), .DIN1(g1514), .DIN2(n2068) );
nnd2s1 U2546 ( .Q(n2068), .DIN1(n2047), .DIN2(n1419) );
hi1s1 U2547 ( .Q(n2047), .DIN(n2125) );
nnd4s1 U2548 ( .Q(n2125), .DIN1(g1514), .DIN2(g1509), .DIN3(g1504), .DIN4(n2127) );
hi1s1 U2549 ( .Q(n2127), .DIN(n2128) );
nor2s1 U2550 ( .Q(g7774), .DIN1(n2129), .DIN2(n1994) );
hi1s1 U2551 ( .Q(n2129), .DIN(n2130) );
xor2s1 U2552 ( .Q(n2130), .DIN1(g1509), .DIN2(n2126) );
and2s1 U2553 ( .Q(n2126), .DIN1(n2131), .DIN2(g1504) );
nor2s1 U2554 ( .Q(g7773), .DIN1(n2132), .DIN2(n1994) );
xor2s1 U2555 ( .Q(n2132), .DIN1(n2133), .DIN2(g1504) );
nor2s1 U2556 ( .Q(g7772), .DIN1(n2134), .DIN2(n1994) );
and2s1 U2557 ( .Q(n2134), .DIN1(n2135), .DIN2(n2136) );
nnd3s1 U2558 ( .Q(n2136), .DIN1(g1494), .DIN2(n2128), .DIN3(n2137) );
nnd2s1 U2559 ( .Q(n2135), .DIN1(g1499), .DIN2(n2133) );
hi1s1 U2560 ( .Q(n2133), .DIN(n2131) );
nor2s1 U2561 ( .Q(g7771), .DIN1(n2138), .DIN2(n1994) );
hi1s1 U2562 ( .Q(n2138), .DIN(n2139) );
xor2s1 U2563 ( .Q(n2139), .DIN1(g1494), .DIN2(n2137) );
nor2s1 U2564 ( .Q(n2137), .DIN1(n2140), .DIN2(n1455) );
nor2s1 U2565 ( .Q(g7770), .DIN1(n2141), .DIN2(n1994) );
xor2s1 U2566 ( .Q(n2141), .DIN1(n2140), .DIN2(g1489) );
nnd2s1 U2567 ( .Q(n2140), .DIN1(g1481), .DIN2(n1419) );
nor2s1 U2568 ( .Q(g7769), .DIN1(n1994), .DIN2(n2142) );
xor2s1 U2569 ( .Q(n2142), .DIN1(g4659), .DIN2(g1481) );
nnd2s1 U2570 ( .Q(n1994), .DIN1(n2111), .DIN2(n2143) );
nnd2s1 U2571 ( .Q(n2143), .DIN1(n2144), .DIN2(n2145) );
xor2s1 U2572 ( .Q(n2145), .DIN1(g1911), .DIN2(g1513) );
hi1s1 U2573 ( .Q(n2144), .DIN(n2109) );
or2s1 U2574 ( .Q(n2111), .DIN1(n2146), .DIN2(n2147) );
nnd4s1 U2575 ( .Q(n2147), .DIN1(g1519), .DIN2(g1472), .DIN3(n2148), .DIN4(n2149) );
or2s1 U2576 ( .Q(n2149), .DIN1(g1514), .DIN2(g174) );
nnd2s1 U2577 ( .Q(n2148), .DIN1(g174), .DIN2(n2150) );
nnd2s1 U2578 ( .Q(n2150), .DIN1(g1504), .DIN2(g1477) );
nnd4s1 U2579 ( .Q(n2146), .DIN1(g1467), .DIN2(g1462), .DIN3(n2131), .DIN4(n2109) );
nnd2s1 U2580 ( .Q(n2109), .DIN1(g150), .DIN2(n1401) );
nor2s1 U2581 ( .Q(n2131), .DIN1(n2128), .DIN2(g4659) );
nnd4s1 U2582 ( .Q(n2128), .DIN1(g1499), .DIN2(g1494), .DIN3(g1489), .DIN4(g1481) );
and3s1 U2583 ( .Q(g7768), .DIN1(n2151), .DIN2(n2072), .DIN3(g1247) );
nnd3s1 U2584 ( .Q(n2072), .DIN1(g1351), .DIN2(n2152), .DIN3(g1354) );
nnd2s1 U2585 ( .Q(n2151), .DIN1(n1430), .DIN2(n2153) );
nnd2s1 U2586 ( .Q(n2153), .DIN1(g1351), .DIN2(n2152) );
nnd4s1 U2587 ( .Q(g7767), .DIN1(n2154), .DIN2(DFF_562net787), .DIN3(n2155), .DIN4(DFF_576net801) );
nor2s1 U2588 ( .Q(n2155), .DIN1(g7425), .DIN2(g7424) );
nnd3s1 U2589 ( .Q(g7766), .DIN1(n2156), .DIN2(n2157), .DIN3(n1402) );
or2s1 U2590 ( .Q(n2157), .DIN1(n2158), .DIN2(g1118) );
nnd2s1 U2591 ( .Q(n2156), .DIN1(g1118), .DIN2(n2113) );
hi1s1 U2592 ( .Q(n2113), .DIN(n2078) );
nor2s1 U2593 ( .Q(n2078), .DIN1(n2158), .DIN2(n1453) );
nnd2s1 U2594 ( .Q(g7765), .DIN1(n2159), .DIN2(n2160) );
nnd3s1 U2595 ( .Q(n2160), .DIN1(n2161), .DIN2(n2117), .DIN3(n1915) );
nnd2s1 U2596 ( .Q(n2159), .DIN1(g1041), .DIN2(n2116) );
nnd2s1 U2597 ( .Q(n2116), .DIN1(n2000), .DIN2(n2162) );
nnd2s1 U2598 ( .Q(n2162), .DIN1(n2117), .DIN2(n1920) );
nnd2s1 U2599 ( .Q(n2117), .DIN1(g1041), .DIN2(n2161) );
hi1s1 U2600 ( .Q(n2161), .DIN(n2163) );
hi1s1 U2601 ( .Q(g7764), .DIN(n2003) );
nnd3s1 U2602 ( .Q(n2003), .DIN1(n2104), .DIN2(g6851), .DIN3(g976) );
xor2s1 U2603 ( .Q(g7762), .DIN1(g828), .DIN2(n2164) );
xor2s1 U2604 ( .Q(g7761), .DIN1(g819), .DIN2(g815) );
nor2s1 U2605 ( .Q(g7759), .DIN1(n2165), .DIN2(n2166) );
nor2s1 U2606 ( .Q(n2165), .DIN1(n2167), .DIN2(g775) );
and2s1 U2607 ( .Q(n2167), .DIN1(n2168), .DIN2(g812) );
nor2s1 U2608 ( .Q(g7758), .DIN1(n2169), .DIN2(n2166) );
xor2s1 U2609 ( .Q(n2169), .DIN1(g812), .DIN2(n2170) );
nnd2s1 U2610 ( .Q(g7757), .DIN1(n2171), .DIN2(n2172) );
nnd3s1 U2611 ( .Q(n2172), .DIN1(n2173), .DIN2(g799), .DIN3(n1463) );
nnd2s1 U2612 ( .Q(n2171), .DIN1(g7756), .DIN2(g803) );
nor2s1 U2613 ( .Q(g7756), .DIN1(n2166), .DIN2(g799) );
nnd2s1 U2614 ( .Q(n1864), .DIN1(n2179), .DIN2(n1849) );
nor2s1 U2615 ( .Q(n1849), .DIN1(n1431), .DIN2(g68) );
nnd2s1 U2616 ( .Q(n1865), .DIN1(n2179), .DIN2(n1839) );
nor2s1 U2617 ( .Q(n1839), .DIN1(n1431), .DIN2(n1397) );
nnd2s1 U2618 ( .Q(n1888), .DIN1(n1895), .DIN2(n1874) );
and3s1 U2619 ( .Q(n1895), .DIN1(n1391), .DIN2(n1409), .DIN3(n1908) );
and2s1 U2620 ( .Q(n1908), .DIN1(n1898), .DIN2(n1444) );
nor3s1 U2621 ( .Q(n1898), .DIN1(g83), .DIN2(g86), .DIN3(g52) );
nor2s1 U2622 ( .Q(g7733), .DIN1(n1541), .DIN2(n2195) );
and2s1 U2623 ( .Q(n2195), .DIN1(n2196), .DIN2(n1540) );
and2s1 U2624 ( .Q(n1540), .DIN1(n2197), .DIN2(g47) );
nor2s1 U2625 ( .Q(n1541), .DIN1(n2197), .DIN2(n2198) );
and2s1 U2626 ( .Q(n2198), .DIN1(g47), .DIN2(n2196) );
xor2s1 U2627 ( .Q(n2197), .DIN1(n2199), .DIN2(n2200) );
xor2s1 U2628 ( .Q(n2200), .DIN1(n2201), .DIN2(n2202) );
xor2s1 U2629 ( .Q(n2202), .DIN1(n1387), .DIN2(n1511) );
xor2s1 U2630 ( .Q(n2201), .DIN1(n1386), .DIN2(n1497) );
xor2s1 U2631 ( .Q(n2199), .DIN1(n2203), .DIN2(n2204) );
xor2s1 U2632 ( .Q(n2204), .DIN1(n1520), .DIN2(n1447) );
hi1s1 U2633 ( .Q(n2203), .DIN(n2205) );
xor2s1 U2634 ( .Q(n2205), .DIN1(n1523), .DIN2(n1500) );
and2s1 U2635 ( .Q(g7530), .DIN1(n2206), .DIN2(g1247) );
xor2s1 U2636 ( .Q(n2206), .DIN1(g1351), .DIN2(n2152) );
nor2s1 U2637 ( .Q(n2152), .DIN1(n1424), .DIN2(n2207) );
nor2s1 U2638 ( .Q(g7529), .DIN1(n2208), .DIN2(n1403) );
xor2s1 U2639 ( .Q(n2208), .DIN1(g1348), .DIN2(n2207) );
and3s1 U2640 ( .Q(g7528), .DIN1(n2209), .DIN2(n2207), .DIN3(g1247) );
or2s1 U2641 ( .Q(n2207), .DIN1(n1406), .DIN2(n2210) );
nnd2s1 U2642 ( .Q(n2209), .DIN1(n1406), .DIN2(n2210) );
nnd3s1 U2643 ( .Q(g7527), .DIN1(n2211), .DIN2(n1422), .DIN3(n2212) );
xor2s1 U2644 ( .Q(n2212), .DIN1(g3851), .DIN2(n2213) );
nnd2s1 U2645 ( .Q(n2213), .DIN1(g1307), .DIN2(n2214) );
hi1s1 U2646 ( .Q(g7526), .DIN(n2154) );
nnd2s1 U2647 ( .Q(n2154), .DIN1(g1142), .DIN2(n2076) );
hi1s1 U2648 ( .Q(n2076), .DIN(n2077) );
nnd4s1 U2649 ( .Q(n2077), .DIN1(g1126), .DIN2(g1122), .DIN3(g1118), .DIN4(n2215) );
nnd2s1 U2650 ( .Q(g7525), .DIN1(n2216), .DIN2(n2217) );
nnd2s1 U2651 ( .Q(n2217), .DIN1(g1149), .DIN2(n2218) );
nnd3s1 U2652 ( .Q(n2216), .DIN1(n1915), .DIN2(n2219), .DIN3(n1462) );
nnd2s1 U2653 ( .Q(g7524), .DIN1(n2220), .DIN2(n2221) );
nnd3s1 U2654 ( .Q(n2221), .DIN1(n2222), .DIN2(n2223), .DIN3(n1915) );
nnd2s1 U2655 ( .Q(n2220), .DIN1(g1138), .DIN2(n2218) );
nnd2s1 U2656 ( .Q(n2218), .DIN1(n2000), .DIN2(n2224) );
nnd2s1 U2657 ( .Q(n2224), .DIN1(n2223), .DIN2(n1920) );
nnd2s1 U2658 ( .Q(g7523), .DIN1(n2225), .DIN2(n2226) );
nnd4s1 U2659 ( .Q(n2226), .DIN1(n1915), .DIN2(g1130), .DIN3(g1092), .DIN4(n2227) );
nnd2s1 U2660 ( .Q(n2225), .DIN1(g1134), .DIN2(n2228) );
nnd2s1 U2661 ( .Q(n2228), .DIN1(n2000), .DIN2(n2229) );
nnd2s1 U2662 ( .Q(n2229), .DIN1(n2227), .DIN2(n1920) );
nnd2s1 U2663 ( .Q(g7522), .DIN1(n2230), .DIN2(n2231) );
nnd2s1 U2664 ( .Q(n2231), .DIN1(g1130), .DIN2(n2232) );
nnd2s1 U2665 ( .Q(n2232), .DIN1(n2000), .DIN2(n2233) );
nnd2s1 U2666 ( .Q(n2233), .DIN1(n1920), .DIN2(n1441) );
nnd3s1 U2667 ( .Q(n2230), .DIN1(n1915), .DIN2(g1092), .DIN3(n1461) );
nnd3s1 U2668 ( .Q(g7521), .DIN1(n2234), .DIN2(n1402), .DIN3(n2235) );
nnd2s1 U2669 ( .Q(n2235), .DIN1(g1114), .DIN2(n2158) );
nnd2s1 U2670 ( .Q(n2158), .DIN1(g1148), .DIN2(n2215) );
hi1s1 U2671 ( .Q(n2215), .DIN(n2236) );
nnd3s1 U2672 ( .Q(n2234), .DIN1(g1110), .DIN2(n2236), .DIN3(n2237) );
hi1s1 U2673 ( .Q(n2237), .DIN(n2238) );
nnd3s1 U2674 ( .Q(n2236), .DIN1(g1110), .DIN2(n2239), .DIN3(g1114) );
nnd2s1 U2675 ( .Q(g7520), .DIN1(n2240), .DIN2(n2241) );
nnd2s1 U2676 ( .Q(n2241), .DIN1(n1915), .DIN2(n1441) );
nnd2s1 U2677 ( .Q(n2240), .DIN1(n1912), .DIN2(g1092) );
hi1s1 U2678 ( .Q(n1912), .DIN(n2000) );
nnd2s1 U2679 ( .Q(g7519), .DIN1(n2242), .DIN2(n2243) );
nnd4s1 U2680 ( .Q(n2243), .DIN1(n1915), .DIN2(g1149), .DIN3(n2219), .DIN4(n2163) );
nor2s1 U2681 ( .Q(n1915), .DIN1(n2244), .DIN2(n2245) );
nnd2s1 U2682 ( .Q(n2242), .DIN1(g1037), .DIN2(n2246) );
nnd2s1 U2683 ( .Q(n2246), .DIN1(n2000), .DIN2(n2247) );
nnd2s1 U2684 ( .Q(n2247), .DIN1(n2163), .DIN2(n1920) );
nnd3s1 U2685 ( .Q(n2163), .DIN1(g1037), .DIN2(n2219), .DIN3(g1149) );
hi1s1 U2686 ( .Q(n2219), .DIN(n2223) );
nnd2s1 U2687 ( .Q(n2223), .DIN1(g1138), .DIN2(n2222) );
hi1s1 U2688 ( .Q(n2222), .DIN(n2227) );
nnd3s1 U2689 ( .Q(n2227), .DIN1(g1130), .DIN2(g1092), .DIN3(g1134) );
nnd2s1 U2690 ( .Q(n2000), .DIN1(n1920), .DIN2(n2244) );
nnd2s1 U2691 ( .Q(n2244), .DIN1(g1158), .DIN2(n1419) );
hi1s1 U2692 ( .Q(n1920), .DIN(n2245) );
nor2s1 U2693 ( .Q(n2245), .DIN1(n1396), .DIN2(n1407) );
nor3s1 U2694 ( .Q(g7518), .DIN1(g6565), .DIN2(g146), .DIN3(n1401) );
nor2s1 U2695 ( .Q(g7517), .DIN1(g6851), .DIN2(n2248) );
xor2s1 U2696 ( .Q(n2248), .DIN1(g995), .DIN2(n2249) );
nnd2s1 U2697 ( .Q(n2249), .DIN1(g990), .DIN2(g985) );
nor2s1 U2698 ( .Q(g7516), .DIN1(g6851), .DIN2(n2250) );
xor2s1 U2699 ( .Q(n2250), .DIN1(n1393), .DIN2(g990) );
and3s1 U2700 ( .Q(g7515), .DIN1(I5528), .DIN2(n1393), .DIN3(n2037) );
nnd3s1 U2701 ( .Q(n2037), .DIN1(n1393), .DIN2(n1464), .DIN3(g995) );
nnd2s1 U2702 ( .Q(g7513), .DIN1(n2251), .DIN2(n2252) );
nnd2s1 U2703 ( .Q(n2252), .DIN1(g825), .DIN2(n2253) );
nnd2s1 U2704 ( .Q(n2251), .DIN1(n2254), .DIN2(n2255) );
nnd2s1 U2705 ( .Q(n2255), .DIN1(g825), .DIN2(n2256) );
nnd2s1 U2706 ( .Q(n2256), .DIN1(g786), .DIN2(g828) );
nnd2s1 U2707 ( .Q(g7512), .DIN1(n2257), .DIN2(n2258) );
nnd3s1 U2708 ( .Q(n2258), .DIN1(n2164), .DIN2(g828), .DIN3(g786) );
nnd2s1 U2709 ( .Q(n2257), .DIN1(n2259), .DIN2(n2253) );
nnd2s1 U2710 ( .Q(n2259), .DIN1(n1472), .DIN2(n2260) );
nnd2s1 U2711 ( .Q(n2260), .DIN1(g819), .DIN2(g815) );
nnd2s1 U2712 ( .Q(g7511), .DIN1(n2173), .DIN2(n2261) );
nnd2s1 U2713 ( .Q(n2261), .DIN1(n2262), .DIN2(n2170) );
hi1s1 U2714 ( .Q(n2170), .DIN(n2168) );
nnd2s1 U2715 ( .Q(n2262), .DIN1(n1437), .DIN2(n2263) );
nnd2s1 U2716 ( .Q(g7510), .DIN1(n2264), .DIN2(n2173) );
hi1s1 U2717 ( .Q(n2173), .DIN(n2166) );
nnd2s1 U2718 ( .Q(n2166), .DIN1(g781), .DIN2(n2265) );
xor2s1 U2719 ( .Q(n2264), .DIN1(g806), .DIN2(n2266) );
nnd2s1 U2720 ( .Q(n2266), .DIN1(g803), .DIN2(g799) );
nor4s1 U2721 ( .Q(g7509), .DIN1(n2196), .DIN2(g41), .DIN3(g42), .DIN4(g55) );
nnd2s1 U2722 ( .Q(n2196), .DIN1(g44), .DIN2(n2041) );
xor2s1 U2723 ( .Q(g7322), .DIN1(n2267), .DIN2(g786) );
and2s1 U2724 ( .Q(n2267), .DIN1(n2164), .DIN2(g828) );
and2s1 U2725 ( .Q(n2164), .DIN1(g825), .DIN2(n2254) );
hi1s1 U2726 ( .Q(n2254), .DIN(n2253) );
nnd3s1 U2727 ( .Q(n2253), .DIN1(g819), .DIN2(g815), .DIN3(g822) );
nnd2s1 U2728 ( .Q(g7309), .DIN1(n2268), .DIN2(n2269) );
nnd2s1 U2729 ( .Q(n2269), .DIN1(n2270), .DIN2(n1504) );
xor2s1 U2730 ( .Q(n2270), .DIN1(n2271), .DIN2(n1427) );
nnd2s1 U2731 ( .Q(n2268), .DIN1(g93), .DIN2(n1505) );
nor2s1 U2732 ( .Q(g7308), .DIN1(g1329), .DIN2(n2272) );
nor2s1 U2733 ( .Q(n2272), .DIN1(n2273), .DIN2(g13) );
nor2s1 U2734 ( .Q(n2273), .DIN1(n1427), .DIN2(n2271) );
nnd2s1 U2735 ( .Q(g7307), .DIN1(n2274), .DIN2(n2275) );
nnd3s1 U2736 ( .Q(n2275), .DIN1(n2276), .DIN2(n2271), .DIN3(n1504) );
nnd3s1 U2737 ( .Q(n2271), .DIN1(g1326), .DIN2(n2277), .DIN3(g1327) );
nnd2s1 U2738 ( .Q(n2276), .DIN1(n1473), .DIN2(n2278) );
nnd2s1 U2739 ( .Q(n2278), .DIN1(g1326), .DIN2(n2277) );
nnd2s1 U2740 ( .Q(n2274), .DIN1(g98), .DIN2(n1505) );
nnd2s1 U2741 ( .Q(g7306), .DIN1(n2279), .DIN2(n2280) );
nnd2s1 U2742 ( .Q(n2280), .DIN1(n2281), .DIN2(n1504) );
xor2s1 U2743 ( .Q(n2281), .DIN1(g1326), .DIN2(n2277) );
and2s1 U2744 ( .Q(n2277), .DIN1(g1325), .DIN2(n2282) );
nnd2s1 U2745 ( .Q(n2279), .DIN1(g103), .DIN2(g1329) );
nnd2s1 U2746 ( .Q(g7305), .DIN1(n2283), .DIN2(n2284) );
nnd2s1 U2747 ( .Q(n2284), .DIN1(n2285), .DIN2(n1504) );
xor2s1 U2748 ( .Q(n2285), .DIN1(n2282), .DIN2(g1325) );
nnd2s1 U2749 ( .Q(n2283), .DIN1(g108), .DIN2(g1329) );
nor2s1 U2750 ( .Q(g7304), .DIN1(g1304), .DIN2(n2286) );
xor2s1 U2751 ( .Q(n2286), .DIN1(g3847), .DIN2(n2287) );
nnd2s1 U2752 ( .Q(n2287), .DIN1(n2288), .DIN2(g3848) );
hi1s1 U2753 ( .Q(n2288), .DIN(n2289) );
nor2s1 U2754 ( .Q(g7303), .DIN1(g1304), .DIN2(n2290) );
xor2s1 U2755 ( .Q(n2290), .DIN1(n2289), .DIN2(g3848) );
and2s1 U2756 ( .Q(g7302), .DIN1(n2291), .DIN2(n1422) );
nnd2s1 U2757 ( .Q(n2291), .DIN1(n2292), .DIN2(n2293) );
nnd4s1 U2758 ( .Q(n2293), .DIN1(g1307), .DIN2(g3851), .DIN3(n2214), .DIN4(n2294) );
nnd2s1 U2759 ( .Q(n2292), .DIN1(g3850), .DIN2(n2289) );
nnd2s1 U2760 ( .Q(n2289), .DIN1(g1307), .DIN2(n2295) );
nor2s1 U2761 ( .Q(g7301), .DIN1(g1304), .DIN2(n2296) );
xor2s1 U2762 ( .Q(n2296), .DIN1(g3852), .DIN2(n2297) );
nnd2s1 U2763 ( .Q(n2297), .DIN1(n2298), .DIN2(g3844) );
nnd2s1 U2764 ( .Q(g7300), .DIN1(n1400), .DIN2(n2299) );
nnd2s1 U2765 ( .Q(n2299), .DIN1(g1254), .DIN2(n2300) );
xor2s1 U2766 ( .Q(n2300), .DIN1(n2301), .DIN2(n1480) );
nnd2s1 U2767 ( .Q(g7299), .DIN1(n2302), .DIN2(n1402) );
xor2s1 U2768 ( .Q(n2302), .DIN1(g1110), .DIN2(n2238) );
hi1s1 U2769 ( .Q(g7296), .DIN(n2303) );
xor2s1 U2770 ( .Q(n2303), .DIN1(n2265), .DIN2(g778) );
nnd3s1 U2771 ( .Q(n2265), .DIN1(g775), .DIN2(n2168), .DIN3(g812) );
nor2s1 U2772 ( .Q(n2168), .DIN1(n1437), .DIN2(n2263) );
nnd3s1 U2773 ( .Q(n2263), .DIN1(g803), .DIN2(g799), .DIN3(g806) );
nor2s1 U2774 ( .Q(g7252), .DIN1(g7104), .DIN2(n1401) );
nnd2s1 U2775 ( .Q(g7248), .DIN1(n2041), .DIN2(n2304) );
nnd2s1 U2776 ( .Q(n2304), .DIN1(n1388), .DIN2(n1443) );
hi1s1 U2777 ( .Q(n2041), .DIN(g8955) );
and3s1 U2778 ( .Q(g7119), .DIN1(n2305), .DIN2(n2210), .DIN3(g1247) );
nnd3s1 U2779 ( .Q(n2210), .DIN1(g1339), .DIN2(n2306), .DIN3(g1342) );
nnd2s1 U2780 ( .Q(n2305), .DIN1(n1410), .DIN2(n2307) );
nnd2s1 U2781 ( .Q(n2307), .DIN1(g1339), .DIN2(n2306) );
nnd2s1 U2782 ( .Q(g7118), .DIN1(n2308), .DIN2(n2309) );
nnd3s1 U2783 ( .Q(n2309), .DIN1(n2310), .DIN2(n2311), .DIN3(n1504) );
hi1s1 U2784 ( .Q(n2311), .DIN(n2282) );
nor2s1 U2785 ( .Q(n2282), .DIN1(n1438), .DIN2(n2312) );
nnd2s1 U2786 ( .Q(n2310), .DIN1(n1438), .DIN2(n2312) );
or2s1 U2787 ( .Q(n2312), .DIN1(n1436), .DIN2(n2313) );
nnd2s1 U2788 ( .Q(n2308), .DIN1(g113), .DIN2(n1505) );
nnd2s1 U2789 ( .Q(g7117), .DIN1(n2314), .DIN2(n2315) );
nnd2s1 U2790 ( .Q(n2315), .DIN1(n2316), .DIN2(n1504) );
xor2s1 U2791 ( .Q(n2316), .DIN1(n2313), .DIN2(n1436) );
nnd2s1 U2792 ( .Q(n2313), .DIN1(g1322), .DIN2(n2317) );
nnd2s1 U2793 ( .Q(n2314), .DIN1(g117), .DIN2(g1329) );
nnd2s1 U2794 ( .Q(g7116), .DIN1(n2318), .DIN2(n2319) );
nnd2s1 U2795 ( .Q(n2319), .DIN1(n2320), .DIN2(n1504) );
xor2s1 U2796 ( .Q(n2320), .DIN1(g1322), .DIN2(n2317) );
nnd2s1 U2797 ( .Q(n2318), .DIN1(g121), .DIN2(g1329) );
nnd2s1 U2798 ( .Q(g7115), .DIN1(n2321), .DIN2(n2322) );
nnd3s1 U2799 ( .Q(n2322), .DIN1(n2323), .DIN2(n2324), .DIN3(n1504) );
hi1s1 U2800 ( .Q(n2324), .DIN(n2317) );
nor2s1 U2801 ( .Q(n2317), .DIN1(n1439), .DIN2(n2325) );
nnd2s1 U2802 ( .Q(n2323), .DIN1(n1439), .DIN2(n2325) );
nnd3s1 U2803 ( .Q(n2325), .DIN1(g1319), .DIN2(n2326), .DIN3(g1320) );
nnd2s1 U2804 ( .Q(n2321), .DIN1(g125), .DIN2(g1329) );
nnd2s1 U2805 ( .Q(g7114), .DIN1(n2327), .DIN2(n2328) );
nnd2s1 U2806 ( .Q(n2328), .DIN1(n2329), .DIN2(n1504) );
xor2s1 U2807 ( .Q(n2329), .DIN1(g1320), .DIN2(n2330) );
and2s1 U2808 ( .Q(n2330), .DIN1(n2326), .DIN2(g1319) );
nnd2s1 U2809 ( .Q(n2327), .DIN1(g129), .DIN2(g1329) );
nnd2s1 U2810 ( .Q(g7113), .DIN1(n2331), .DIN2(n2332) );
nnd2s1 U2811 ( .Q(n2332), .DIN1(n2333), .DIN2(n1504) );
xor2s1 U2812 ( .Q(n2333), .DIN1(g1319), .DIN2(n2326) );
hi1s1 U2813 ( .Q(n2326), .DIN(n2334) );
nnd2s1 U2814 ( .Q(n2331), .DIN1(g133), .DIN2(n1505) );
and2s1 U2815 ( .Q(g7112), .DIN1(n1422), .DIN2(n2335) );
xor2s1 U2816 ( .Q(n2335), .DIN1(n2298), .DIN2(g3844) );
nor2s1 U2817 ( .Q(n2298), .DIN1(n2336), .DIN2(n1449) );
nnd2s1 U2818 ( .Q(g7111), .DIN1(g1253), .DIN2(n2337) );
and4s1 U2819 ( .Q(g7110), .DIN1(g1254), .DIN2(n2338), .DIN3(n2301), .DIN4(n1400) );
nnd3s1 U2820 ( .Q(n2301), .DIN1(n1489), .DIN2(n2339), .DIN3(n1507) );
nnd2s1 U2821 ( .Q(n2338), .DIN1(n1488), .DIN2(n2340) );
nnd2s1 U2822 ( .Q(n2340), .DIN1(n1507), .DIN2(n2339) );
nnd2s1 U2823 ( .Q(g7109), .DIN1(n2341), .DIN2(n1400) );
xor2s1 U2824 ( .Q(n2341), .DIN1(n1506), .DIN2(n2339) );
nor2s1 U2825 ( .Q(n2339), .DIN1(n1490), .DIN2(n2342) );
nnd2s1 U2826 ( .Q(g7108), .DIN1(n2343), .DIN2(n1400) );
xor2s1 U2827 ( .Q(n2343), .DIN1(n1491), .DIN2(n2342) );
nnd3s1 U2828 ( .Q(g7107), .DIN1(n2344), .DIN2(n1402), .DIN3(n2345) );
nnd2s1 U2829 ( .Q(n2345), .DIN1(g1106), .DIN2(n2238) );
nnd2s1 U2830 ( .Q(n2238), .DIN1(g1148), .DIN2(n2239) );
hi1s1 U2831 ( .Q(n2239), .DIN(n2346) );
nnd3s1 U2832 ( .Q(n2344), .DIN1(g1102), .DIN2(n2346), .DIN3(n2347) );
nnd4s1 U2833 ( .Q(n2346), .DIN1(g1106), .DIN2(g1102), .DIN3(g1098), .DIN4(g1087) );
xor2s1 U2834 ( .Q(g7106), .DIN1(g2888), .DIN2(n2348) );
nnd2s1 U2835 ( .Q(n2348), .DIN1(n2349), .DIN2(n2350) );
nnd3s1 U2836 ( .Q(n2350), .DIN1(g652), .DIN2(g1158), .DIN3(g1179) );
nor2s1 U2837 ( .Q(g7105), .DIN1(I5528), .DIN2(g162) );
and3s1 U2838 ( .Q(g7104), .DIN1(g6851), .DIN2(n1475), .DIN3(g984) );
nnd2s1 U2839 ( .Q(g7102), .DIN1(n2351), .DIN2(n2352) );
nnd2s1 U2840 ( .Q(n2352), .DIN1(g11), .DIN2(n1469) );
nnd2s1 U2841 ( .Q(n2351), .DIN1(g12), .DIN2(g859) );
nnd3s1 U2842 ( .Q(g7101), .DIN1(n2353), .DIN2(n2354), .DIN3(n2355) );
nnd4s1 U2843 ( .Q(n2354), .DIN1(g889), .DIN2(g887), .DIN3(g874), .DIN4(n1405) );
nnd2s1 U2844 ( .Q(n2353), .DIN1(n2356), .DIN2(n1468) );
nnd2s1 U2845 ( .Q(n2356), .DIN1(n2357), .DIN2(n2358) );
or4s1 U2846 ( .Q(n2358), .DIN1(n1405), .DIN2(n2359), .DIN3(g866), .DIN4(g875) );
nnd2s1 U2847 ( .Q(n2357), .DIN1(n2360), .DIN2(n2361) );
nnd2s1 U2848 ( .Q(n2361), .DIN1(n1417), .DIN2(n2362) );
nnd2s1 U2849 ( .Q(n2362), .DIN1(n2363), .DIN2(n2364) );
nnd2s1 U2850 ( .Q(n2363), .DIN1(n1465), .DIN2(n2365) );
nnd3s1 U2851 ( .Q(g7100), .DIN1(n2366), .DIN2(n2367), .DIN3(n2355) );
nnd2s1 U2852 ( .Q(n2355), .DIN1(g4302), .DIN2(n2364) );
nnd3s1 U2853 ( .Q(n2367), .DIN1(n2360), .DIN2(g889), .DIN3(g866) );
nnd3s1 U2854 ( .Q(n2366), .DIN1(n2368), .DIN2(n2369), .DIN3(n2370) );
nnd2s1 U2855 ( .Q(n2369), .DIN1(g4316), .DIN2(n1405) );
nnd2s1 U2856 ( .Q(n2368), .DIN1(g875), .DIN2(g888) );
nnd3s1 U2857 ( .Q(g7099), .DIN1(n2371), .DIN2(n2359), .DIN3(n2372) );
nnd2s1 U2858 ( .Q(n2372), .DIN1(g887), .DIN2(n2364) );
hi1s1 U2859 ( .Q(n2359), .DIN(n2370) );
nnd2s1 U2860 ( .Q(n2371), .DIN1(n2373), .DIN2(n1405) );
nnd3s1 U2861 ( .Q(n2373), .DIN1(n2374), .DIN2(n1432), .DIN3(n2375) );
nnd2s1 U2862 ( .Q(n2375), .DIN1(g3855), .DIN2(n2376) );
nnd2s1 U2863 ( .Q(n2376), .DIN1(g4654), .DIN2(n1417) );
nnd4s1 U2864 ( .Q(n2374), .DIN1(g866), .DIN2(n2365), .DIN3(n2364), .DIN4(n1417) );
or2s1 U2865 ( .Q(n2365), .DIN1(n2377), .DIN2(n2378) );
nnd4s1 U2866 ( .Q(n2378), .DIN1(n1423), .DIN2(n1395), .DIN3(n1383), .DIN4(n1380) );
nnd4s1 U2867 ( .Q(n2377), .DIN1(n1421), .DIN2(n1394), .DIN3(n1382), .DIN4(n1379) );
nor2s1 U2868 ( .Q(g7071), .DIN1(n2034), .DIN2(n2104) );
hi1s1 U2869 ( .Q(n2034), .DIN(g6310) );
nnd2s1 U2870 ( .Q(g6952), .DIN1(n2379), .DIN2(n2380) );
nnd2s1 U2871 ( .Q(n2380), .DIN1(g31), .DIN2(n2381) );
hi1s1 U2872 ( .Q(n2381), .DIN(g32) );
nnd2s1 U2873 ( .Q(n2379), .DIN1(g30), .DIN2(g32) );
xor2s1 U2874 ( .Q(g6891), .DIN1(g611), .DIN2(n1507) );
xor2s1 U2875 ( .Q(g6890), .DIN1(g612), .DIN2(n1491) );
xor2s1 U2876 ( .Q(g6889), .DIN1(g613), .DIN2(n1478) );
xor2s1 U2877 ( .Q(g6888), .DIN1(g614), .DIN2(n1483) );
xor2s1 U2878 ( .Q(g6887), .DIN1(g615), .DIN2(n1509) );
xor2s1 U2879 ( .Q(g6886), .DIN1(g616), .DIN2(n1493) );
xor2s1 U2880 ( .Q(g6885), .DIN1(g617), .DIN2(n1503) );
xor2s1 U2881 ( .Q(g6884), .DIN1(g618), .DIN2(n1487) );
xor2s1 U2882 ( .Q(g6883), .DIN1(g619), .DIN2(n1485) );
xor2s1 U2883 ( .Q(g6882), .DIN1(g621), .DIN2(n1514) );
xor2s1 U2884 ( .Q(g6881), .DIN1(g620), .DIN2(n1495) );
xor2s1 U2885 ( .Q(g6880), .DIN1(g610), .DIN2(n1489) );
xor2s1 U2886 ( .Q(g6879), .DIN1(g609), .DIN2(n1481) );
xor2s1 U2887 ( .Q(g6878), .DIN1(g598), .DIN2(n1507) );
xor2s1 U2888 ( .Q(g6877), .DIN1(g599), .DIN2(n1491) );
xor2s1 U2889 ( .Q(g6876), .DIN1(g600), .DIN2(n1478) );
xor2s1 U2890 ( .Q(g6875), .DIN1(g601), .DIN2(n1483) );
xor2s1 U2891 ( .Q(g6874), .DIN1(g602), .DIN2(n1509) );
xor2s1 U2892 ( .Q(g6873), .DIN1(g603), .DIN2(n1493) );
xor2s1 U2893 ( .Q(g6872), .DIN1(g604), .DIN2(n1503) );
xor2s1 U2894 ( .Q(g6871), .DIN1(g605), .DIN2(n1487) );
xor2s1 U2895 ( .Q(g6870), .DIN1(g606), .DIN2(n1485) );
xor2s1 U2896 ( .Q(g6869), .DIN1(g608), .DIN2(n1514) );
xor2s1 U2897 ( .Q(g6868), .DIN1(g607), .DIN2(n1495) );
xor2s1 U2898 ( .Q(g6867), .DIN1(g597), .DIN2(n1489) );
xor2s1 U2899 ( .Q(g6866), .DIN1(g596), .DIN2(n1481) );
nnd2s1 U2900 ( .Q(g6865), .DIN1(n2382), .DIN2(n2383) );
nnd3s1 U2901 ( .Q(n2383), .DIN1(g1247), .DIN2(n2306), .DIN3(n1408) );
nnd2s1 U2902 ( .Q(n2382), .DIN1(n2384), .DIN2(g1339) );
nor2s1 U2903 ( .Q(g6864), .DIN1(n2385), .DIN2(n2386) );
hi1s1 U2904 ( .Q(n2386), .DIN(n2384) );
nor2s1 U2905 ( .Q(n2384), .DIN1(n1403), .DIN2(n2306) );
and3s1 U2906 ( .Q(n2306), .DIN1(g1333), .DIN2(g1330), .DIN3(g1336) );
nor2s1 U2907 ( .Q(n2385), .DIN1(n2387), .DIN2(g1336) );
nor2s1 U2908 ( .Q(n2387), .DIN1(n1411), .DIN2(n1390) );
nnd2s1 U2909 ( .Q(g6863), .DIN1(n2388), .DIN2(n2389) );
nnd3s1 U2910 ( .Q(n2389), .DIN1(g1247), .DIN2(g1330), .DIN3(n1390) );
nnd2s1 U2911 ( .Q(n2388), .DIN1(g6862), .DIN2(g1333) );
nor2s1 U2912 ( .Q(g6862), .DIN1(n1403), .DIN2(g1330) );
nnd2s1 U2913 ( .Q(g6861), .DIN1(n2390), .DIN2(n2391) );
nnd3s1 U2914 ( .Q(n2391), .DIN1(n2392), .DIN2(n2334), .DIN3(n1504) );
nnd3s1 U2915 ( .Q(n2334), .DIN1(g1317), .DIN2(g1313), .DIN3(g1318) );
nnd2s1 U2916 ( .Q(n2392), .DIN1(n1474), .DIN2(n2393) );
nnd2s1 U2917 ( .Q(n2393), .DIN1(g1317), .DIN2(g1313) );
nnd2s1 U2918 ( .Q(n2390), .DIN1(g137), .DIN2(g1329) );
hi1s1 U2919 ( .Q(g6860), .DIN(n2337) );
nnd2s1 U2920 ( .Q(n2337), .DIN1(g1247), .DIN2(n2394) );
nnd2s1 U2921 ( .Q(n2394), .DIN1(n2395), .DIN2(n2396) );
or2s1 U2922 ( .Q(n2396), .DIN1(g1257), .DIN2(g1263) );
nnd2s1 U2923 ( .Q(g6859), .DIN1(n1400), .DIN2(n2397) );
nnd2s1 U2924 ( .Q(n2397), .DIN1(n2398), .DIN2(n2342) );
or2s1 U2925 ( .Q(n2342), .DIN1(n1477), .DIN2(n2399) );
nnd2s1 U2926 ( .Q(n2398), .DIN1(n1477), .DIN2(n2399) );
nnd4s1 U2927 ( .Q(n2399), .DIN1(n1514), .DIN2(n1495), .DIN3(n2400), .DIN4(n2401) );
nnd2s1 U2928 ( .Q(g6858), .DIN1(n2402), .DIN2(n1400) );
xor2s1 U2929 ( .Q(n2402), .DIN1(n1483), .DIN2(n2403) );
nnd2s1 U2930 ( .Q(n2403), .DIN1(n2404), .DIN2(n1509) );
hi1s1 U2931 ( .Q(n2404), .DIN(n2405) );
nnd2s1 U2932 ( .Q(g6857), .DIN1(n2406), .DIN2(n1400) );
xor2s1 U2933 ( .Q(n2406), .DIN1(n1509), .DIN2(n2405) );
nnd2s1 U2934 ( .Q(g6856), .DIN1(n2349), .DIN2(n2407) );
nnd3s1 U2935 ( .Q(n2407), .DIN1(g652), .DIN2(g1158), .DIN3(g1176) );
nnd2s1 U2936 ( .Q(n2349), .DIN1(g2888), .DIN2(g1077) );
and2s1 U2937 ( .Q(g6855), .DIN1(n1402), .DIN2(n2408) );
xor2s1 U2938 ( .Q(n2408), .DIN1(n2347), .DIN2(g1102) );
nor2s1 U2939 ( .Q(n2347), .DIN1(n2409), .DIN2(n1454) );
nor2s1 U2940 ( .Q(g6854), .DIN1(g1097), .DIN2(n2410) );
xor2s1 U2941 ( .Q(n2410), .DIN1(g1098), .DIN2(n2409) );
nnd2s1 U2942 ( .Q(n2409), .DIN1(g1148), .DIN2(g1087) );
and2s1 U2943 ( .Q(g6853), .DIN1(n1402), .DIN2(n2411) );
xor2s1 U2944 ( .Q(n2411), .DIN1(g1148), .DIN2(g1087) );
nnd2s1 U2945 ( .Q(g6852), .DIN1(n2412), .DIN2(n2413) );
or2s1 U2946 ( .Q(n2413), .DIN1(n1445), .DIN2(g1176) );
nnd2s1 U2947 ( .Q(n2412), .DIN1(g1080), .DIN2(n1445) );
nor2s1 U2948 ( .Q(g6745), .DIN1(n2104), .DIN2(g6310) );
nor4s1 U2949 ( .Q(n2104), .DIN1(g962), .DIN2(g1871), .DIN3(g1870), .DIN4(n2414) );
nnd4s1 U2950 ( .Q(n2414), .DIN1(DFF_144net369), .DIN2(DFF_622net847), .DIN3(DFF_381net606), .DIN4(DFF_371net596) );
nnd3s1 U2951 ( .Q(g6565), .DIN1(g6851), .DIN2(n1446), .DIN3(g1033) );
and2s1 U2952 ( .Q(n1671), .DIN1(n2179), .DIN2(n1874) );
nor2s1 U2953 ( .Q(n1874), .DIN1(g68), .DIN2(g71) );
nnd2s1 U2954 ( .Q(n1866), .DIN1(n2179), .DIN2(n1854) );
nor2s1 U2955 ( .Q(n1854), .DIN1(n1397), .DIN2(g71) );
and2s1 U2956 ( .Q(n2179), .DIN1(n1873), .DIN2(n1409) );
and4s1 U2957 ( .Q(n1873), .DIN1(g86), .DIN2(g83), .DIN3(n2415), .DIN4(g52) );
nor2s1 U2958 ( .Q(n2415), .DIN1(g74), .DIN2(n1444) );
or2s1 U2959 ( .Q(g6392), .DIN1(n2416), .DIN2(n2417) );
or4s1 U2960 ( .Q(n2417), .DIN1(n2418), .DIN2(n2419), .DIN3(n2420), .DIN4(n2421) );
xor2s1 U2961 ( .Q(n2421), .DIN1(g3848), .DIN2(g768) );
xor2s1 U2962 ( .Q(n2420), .DIN1(g769), .DIN2(g3850) );
xor2s1 U2963 ( .Q(n2419), .DIN1(g3851), .DIN2(g770) );
xor2s1 U2964 ( .Q(n2418), .DIN1(g771), .DIN2(g3852) );
or4s1 U2965 ( .Q(n2416), .DIN1(n2422), .DIN2(n2423), .DIN3(n2424), .DIN4(n2425) );
xor2s1 U2966 ( .Q(n2425), .DIN1(g3844), .DIN2(g772) );
xor2s1 U2967 ( .Q(n2424), .DIN1(g3845), .DIN2(g773) );
xor2s1 U2968 ( .Q(n2423), .DIN1(g3846), .DIN2(g774) );
xor2s1 U2969 ( .Q(n2422), .DIN1(g767), .DIN2(g3847) );
or4s1 U2970 ( .Q(g6391), .DIN1(n2426), .DIN2(n2427), .DIN3(n2428), .DIN4(n2429) );
nnd4s1 U2971 ( .Q(n2429), .DIN1(n1411), .DIN2(n1390), .DIN3(n2430), .DIN4(n2431) );
and3s1 U2972 ( .Q(n2431), .DIN1(n2432), .DIN2(n2433), .DIN3(n2434) );
xor2s1 U2973 ( .Q(n2434), .DIN1(n1410), .DIN2(g764) );
xor2s1 U2974 ( .Q(n2433), .DIN1(n1406), .DIN2(g763) );
xor2s1 U2975 ( .Q(n2432), .DIN1(n1408), .DIN2(g765) );
xor2s1 U2976 ( .Q(n2430), .DIN1(n1420), .DIN2(g766) );
nnd3s1 U2977 ( .Q(n2428), .DIN1(n2435), .DIN2(n2436), .DIN3(n2437) );
xor2s1 U2978 ( .Q(n2437), .DIN1(g1351), .DIN2(n1425) );
xor2s1 U2979 ( .Q(n2436), .DIN1(n1430), .DIN2(g760) );
xor2s1 U2980 ( .Q(n2435), .DIN1(n1424), .DIN2(g762) );
xor2s1 U2981 ( .Q(n2427), .DIN1(g758), .DIN2(g1360) );
xor2s1 U2982 ( .Q(n2426), .DIN1(g759), .DIN2(g1357) );
or4s1 U2983 ( .Q(g6386), .DIN1(n2438), .DIN2(n2439), .DIN3(n2440), .DIN4(n2441) );
nnd4s1 U2984 ( .Q(n2441), .DIN1(n2442), .DIN2(n2443), .DIN3(n2444), .DIN4(n2445) );
and3s1 U2985 ( .Q(n2445), .DIN1(n2446), .DIN2(n2447), .DIN3(n2448) );
xor2s1 U2986 ( .Q(n2448), .DIN1(n1390), .DIN2(g631) );
xor2s1 U2987 ( .Q(n2447), .DIN1(n1420), .DIN2(g630) );
xor2s1 U2988 ( .Q(n2446), .DIN1(n1411), .DIN2(g632) );
xor2s1 U2989 ( .Q(n2444), .DIN1(n1410), .DIN2(g628) );
xor2s1 U2990 ( .Q(n2443), .DIN1(n1406), .DIN2(g627) );
xor2s1 U2991 ( .Q(n2442), .DIN1(n1408), .DIN2(g629) );
or3s1 U2992 ( .Q(n2440), .DIN1(n2449), .DIN2(n2450), .DIN3(n2451) );
xor2s1 U2993 ( .Q(n2451), .DIN1(g1351), .DIN2(g625) );
xor2s1 U2994 ( .Q(n2450), .DIN1(g1354), .DIN2(g624) );
xor2s1 U2995 ( .Q(n2449), .DIN1(g1348), .DIN2(g626) );
xor2s1 U2996 ( .Q(n2439), .DIN1(g622), .DIN2(g1360) );
xor2s1 U2997 ( .Q(n2438), .DIN1(g623), .DIN2(g1357) );
nnd2s1 U2998 ( .Q(g6385), .DIN1(DFF_373net598), .DIN2(n2452) );
nor2s1 U2999 ( .Q(g6384), .DIN1(g1304), .DIN2(n2453) );
xor2s1 U3000 ( .Q(n2453), .DIN1(g3845), .DIN2(n2336) );
nnd2s1 U3001 ( .Q(n2336), .DIN1(g1307), .DIN2(g3846) );
and2s1 U3002 ( .Q(g6383), .DIN1(n1422), .DIN2(n2454) );
xor2s1 U3003 ( .Q(n2454), .DIN1(g3846), .DIN2(g1307) );
nnd2s1 U3004 ( .Q(g6382), .DIN1(g1266), .DIN2(n2395) );
nnd2s1 U3005 ( .Q(g6381), .DIN1(g1257), .DIN2(n2395) );
nnd2s1 U3006 ( .Q(g6380), .DIN1(g1263), .DIN2(n2395) );
and4s1 U3007 ( .Q(n2395), .DIN1(n2401), .DIN2(n1488), .DIN3(n1478), .DIN4(n2455) );
and3s1 U3008 ( .Q(n2455), .DIN1(n1507), .DIN2(n1491), .DIN3(n1481) );
and3s1 U3009 ( .Q(n2401), .DIN1(n1509), .DIN2(n1483), .DIN3(n1493) );
nnd2s1 U3010 ( .Q(g6379), .DIN1(n1400), .DIN2(n2456) );
nnd2s1 U3011 ( .Q(n2456), .DIN1(n2457), .DIN2(n2405) );
nnd3s1 U3012 ( .Q(n2405), .DIN1(n1493), .DIN2(n2458), .DIN3(n2459) );
nnd2s1 U3013 ( .Q(n2457), .DIN1(n1492), .DIN2(n2460) );
nnd2s1 U3014 ( .Q(n2460), .DIN1(n2459), .DIN2(n2458) );
nnd2s1 U3015 ( .Q(g6378), .DIN1(n2461), .DIN2(n1400) );
xor2s1 U3016 ( .Q(n2461), .DIN1(n1503), .DIN2(n2462) );
nnd2s1 U3017 ( .Q(n2462), .DIN1(n2459), .DIN2(n1487) );
nnd2s1 U3018 ( .Q(g6377), .DIN1(n2463), .DIN2(n1400) );
xor2s1 U3019 ( .Q(n2463), .DIN1(n1486), .DIN2(n2459) );
hi1s1 U3020 ( .Q(n2459), .DIN(n2464) );
nnd2s1 U3021 ( .Q(g6372), .DIN1(n2086), .DIN2(n2465) );
nnd2s1 U3022 ( .Q(n2465), .DIN1(g2801), .DIN2(DFF_605net830) );
or4s1 U3023 ( .Q(g6371), .DIN1(n2466), .DIN2(n2467), .DIN3(n2468), .DIN4(n2469) );
nnd3s1 U3024 ( .Q(n2469), .DIN1(n2470), .DIN2(n2471), .DIN3(n2472) );
nnd2s1 U3025 ( .Q(n2472), .DIN1(g652), .DIN2(g677) );
nnd2s1 U3026 ( .Q(n2471), .DIN1(g647), .DIN2(g681) );
nnd2s1 U3027 ( .Q(n2470), .DIN1(g648), .DIN2(g685) );
nnd4s1 U3028 ( .Q(n2468), .DIN1(n2473), .DIN2(n2474), .DIN3(n2475), .DIN4(n2476) );
nnd2s1 U3029 ( .Q(n2476), .DIN1(g633), .DIN2(g661) );
nnd2s1 U3030 ( .Q(n2475), .DIN1(g634), .DIN2(g665) );
nnd2s1 U3031 ( .Q(n2474), .DIN1(g635), .DIN2(g669) );
nnd2s1 U3032 ( .Q(n2473), .DIN1(g645), .DIN2(g673) );
nnd3s1 U3033 ( .Q(n2467), .DIN1(n2477), .DIN2(n2478), .DIN3(n2479) );
nnd2s1 U3034 ( .Q(n2479), .DIN1(g723), .DIN2(g730) );
nnd2s1 U3035 ( .Q(n2478), .DIN1(g702), .DIN2(g718) );
nnd2s1 U3036 ( .Q(n2477), .DIN1(g722), .DIN2(g734) );
nnd3s1 U3037 ( .Q(n2466), .DIN1(n2480), .DIN2(n2481), .DIN3(n2482) );
nnd2s1 U3038 ( .Q(n2482), .DIN1(g698), .DIN2(g714) );
nnd2s1 U3039 ( .Q(n2481), .DIN1(g690), .DIN2(g706) );
nnd2s1 U3040 ( .Q(n2480), .DIN1(g694), .DIN2(g710) );
nnd2s1 U3041 ( .Q(g6370), .DIN1(n2483), .DIN2(n2484) );
nnd2s1 U3042 ( .Q(n2484), .DIN1(g560), .DIN2(n2485) );
nnd2s1 U3043 ( .Q(n2483), .DIN1(g587), .DIN2(n2486) );
nnd2s1 U3044 ( .Q(g6369), .DIN1(n2487), .DIN2(n2488) );
nnd2s1 U3045 ( .Q(n2488), .DIN1(g584), .DIN2(n2485) );
nnd2s1 U3046 ( .Q(n2487), .DIN1(g583), .DIN2(n2486) );
nnd2s1 U3047 ( .Q(g6368), .DIN1(n2489), .DIN2(n2490) );
nnd2s1 U3048 ( .Q(n2490), .DIN1(g580), .DIN2(n2485) );
nnd2s1 U3049 ( .Q(n2489), .DIN1(g579), .DIN2(n2486) );
nnd2s1 U3050 ( .Q(g6367), .DIN1(n2491), .DIN2(n2492) );
nnd2s1 U3051 ( .Q(n2492), .DIN1(g567), .DIN2(n2485) );
nnd2s1 U3052 ( .Q(n2491), .DIN1(g566), .DIN2(n2486) );
nnd2s1 U3053 ( .Q(g6366), .DIN1(n2493), .DIN2(n2494) );
nnd2s1 U3054 ( .Q(n2494), .DIN1(g557), .DIN2(n2485) );
nnd2s1 U3055 ( .Q(n2493), .DIN1(g556), .DIN2(n2486) );
nnd2s1 U3056 ( .Q(g6365), .DIN1(n2495), .DIN2(n2496) );
nnd2s1 U3057 ( .Q(n2496), .DIN1(g544), .DIN2(n2485) );
nnd2s1 U3058 ( .Q(n2495), .DIN1(g543), .DIN2(n2486) );
nnd2s1 U3059 ( .Q(g6364), .DIN1(n2497), .DIN2(n2498) );
nnd2s1 U3060 ( .Q(n2498), .DIN1(g540), .DIN2(n2485) );
nnd2s1 U3061 ( .Q(n2497), .DIN1(g539), .DIN2(n2486) );
nnd2s1 U3062 ( .Q(g6363), .DIN1(n2499), .DIN2(n2500) );
nnd2s1 U3063 ( .Q(n2500), .DIN1(g536), .DIN2(n2485) );
nnd2s1 U3064 ( .Q(n2499), .DIN1(g535), .DIN2(n2486) );
hi1s1 U3065 ( .Q(n2486), .DIN(n2485) );
nnd2s1 U3066 ( .Q(n2485), .DIN1(g595), .DIN2(DFF_550net775) );
nnd2s1 U3067 ( .Q(g6362), .DIN1(n2501), .DIN2(n2502) );
nnd2s1 U3068 ( .Q(n2502), .DIN1(g521), .DIN2(n2503) );
nnd2s1 U3069 ( .Q(n2501), .DIN1(g517), .DIN2(n2504) );
nnd2s1 U3070 ( .Q(g6361), .DIN1(n2505), .DIN2(n2506) );
nnd2s1 U3071 ( .Q(n2506), .DIN1(g518), .DIN2(n2503) );
nnd2s1 U3072 ( .Q(n2505), .DIN1(g516), .DIN2(n2504) );
nnd2s1 U3073 ( .Q(g6360), .DIN1(n2507), .DIN2(n2508) );
nnd2s1 U3074 ( .Q(n2508), .DIN1(g495), .DIN2(n2503) );
nnd2s1 U3075 ( .Q(n2507), .DIN1(g479), .DIN2(n2504) );
nnd2s1 U3076 ( .Q(g6359), .DIN1(n2509), .DIN2(n2510) );
nnd2s1 U3077 ( .Q(n2510), .DIN1(g492), .DIN2(n2503) );
nnd2s1 U3078 ( .Q(n2509), .DIN1(g478), .DIN2(n2504) );
nnd2s1 U3079 ( .Q(g6358), .DIN1(n2511), .DIN2(n2512) );
nnd2s1 U3080 ( .Q(n2512), .DIN1(g489), .DIN2(n2503) );
nnd2s1 U3081 ( .Q(n2511), .DIN1(g477), .DIN2(n2504) );
nnd2s1 U3082 ( .Q(g6357), .DIN1(n2513), .DIN2(n2514) );
nnd2s1 U3083 ( .Q(n2514), .DIN1(g486), .DIN2(n2503) );
nnd2s1 U3084 ( .Q(n2513), .DIN1(g476), .DIN2(n2504) );
nnd2s1 U3085 ( .Q(g6356), .DIN1(n2515), .DIN2(n2516) );
nnd2s1 U3086 ( .Q(n2516), .DIN1(g483), .DIN2(n2503) );
nnd2s1 U3087 ( .Q(n2515), .DIN1(g475), .DIN2(n2504) );
nnd2s1 U3088 ( .Q(g6355), .DIN1(n2517), .DIN2(n2518) );
nnd2s1 U3089 ( .Q(n2518), .DIN1(g480), .DIN2(n2503) );
nnd2s1 U3090 ( .Q(n2517), .DIN1(g474), .DIN2(n2504) );
nnd2s1 U3091 ( .Q(g6354), .DIN1(n2519), .DIN2(n2520) );
nnd2s1 U3092 ( .Q(n2520), .DIN1(g471), .DIN2(n2503) );
nnd2s1 U3093 ( .Q(n2519), .DIN1(g458), .DIN2(n2504) );
nnd2s1 U3094 ( .Q(g6353), .DIN1(n2521), .DIN2(n2522) );
nnd2s1 U3095 ( .Q(n2522), .DIN1(g468), .DIN2(n2503) );
nnd2s1 U3096 ( .Q(n2521), .DIN1(g457), .DIN2(n2504) );
nnd2s1 U3097 ( .Q(g6352), .DIN1(n2523), .DIN2(n2524) );
nnd2s1 U3098 ( .Q(n2524), .DIN1(g465), .DIN2(n2503) );
nnd2s1 U3099 ( .Q(n2523), .DIN1(g456), .DIN2(n2504) );
nnd2s1 U3100 ( .Q(g6351), .DIN1(n2525), .DIN2(n2526) );
nnd2s1 U3101 ( .Q(n2526), .DIN1(g462), .DIN2(n2503) );
nnd2s1 U3102 ( .Q(n2525), .DIN1(g455), .DIN2(n2504) );
nnd2s1 U3103 ( .Q(g6350), .DIN1(n2527), .DIN2(n2528) );
nnd2s1 U3104 ( .Q(n2528), .DIN1(g459), .DIN2(n2503) );
nnd2s1 U3105 ( .Q(n2527), .DIN1(g454), .DIN2(n2504) );
hi1s1 U3106 ( .Q(n2504), .DIN(n2503) );
nnd2s1 U3107 ( .Q(n2503), .DIN1(g533), .DIN2(DFF_286net511) );
nnd2s1 U3108 ( .Q(g6349), .DIN1(n2529), .DIN2(n2530) );
nnd2s1 U3109 ( .Q(n2530), .DIN1(g440), .DIN2(n2531) );
nnd2s1 U3110 ( .Q(n2529), .DIN1(g436), .DIN2(n2532) );
nnd2s1 U3111 ( .Q(g6348), .DIN1(n2533), .DIN2(n2534) );
nnd2s1 U3112 ( .Q(n2534), .DIN1(g437), .DIN2(n2531) );
nnd2s1 U3113 ( .Q(n2533), .DIN1(g435), .DIN2(n2532) );
nnd2s1 U3114 ( .Q(g6347), .DIN1(n2535), .DIN2(n2536) );
nnd2s1 U3115 ( .Q(n2536), .DIN1(g414), .DIN2(n2531) );
nnd2s1 U3116 ( .Q(n2535), .DIN1(g398), .DIN2(n2532) );
nnd2s1 U3117 ( .Q(g6346), .DIN1(n2537), .DIN2(n2538) );
nnd2s1 U3118 ( .Q(n2538), .DIN1(g411), .DIN2(n2531) );
nnd2s1 U3119 ( .Q(n2537), .DIN1(g397), .DIN2(n2532) );
nnd2s1 U3120 ( .Q(g6345), .DIN1(n2539), .DIN2(n2540) );
nnd2s1 U3121 ( .Q(n2540), .DIN1(g408), .DIN2(n2531) );
nnd2s1 U3122 ( .Q(n2539), .DIN1(g396), .DIN2(n2532) );
nnd2s1 U3123 ( .Q(g6344), .DIN1(n2541), .DIN2(n2542) );
nnd2s1 U3124 ( .Q(n2542), .DIN1(g405), .DIN2(n2531) );
nnd2s1 U3125 ( .Q(n2541), .DIN1(g395), .DIN2(n2532) );
nnd2s1 U3126 ( .Q(g6343), .DIN1(n2543), .DIN2(n2544) );
nnd2s1 U3127 ( .Q(n2544), .DIN1(g402), .DIN2(n2531) );
nnd2s1 U3128 ( .Q(n2543), .DIN1(g394), .DIN2(n2532) );
nnd2s1 U3129 ( .Q(g6342), .DIN1(n2545), .DIN2(n2546) );
nnd2s1 U3130 ( .Q(n2546), .DIN1(g399), .DIN2(n2531) );
nnd2s1 U3131 ( .Q(n2545), .DIN1(g393), .DIN2(n2532) );
nnd2s1 U3132 ( .Q(g6341), .DIN1(n2547), .DIN2(n2548) );
nnd2s1 U3133 ( .Q(n2548), .DIN1(g390), .DIN2(n2531) );
nnd2s1 U3134 ( .Q(n2547), .DIN1(g377), .DIN2(n2532) );
nnd2s1 U3135 ( .Q(g6340), .DIN1(n2549), .DIN2(n2550) );
nnd2s1 U3136 ( .Q(n2550), .DIN1(g387), .DIN2(n2531) );
nnd2s1 U3137 ( .Q(n2549), .DIN1(g376), .DIN2(n2532) );
nnd2s1 U3138 ( .Q(g6339), .DIN1(n2551), .DIN2(n2552) );
nnd2s1 U3139 ( .Q(n2552), .DIN1(g384), .DIN2(n2531) );
nnd2s1 U3140 ( .Q(n2551), .DIN1(g375), .DIN2(n2532) );
nnd2s1 U3141 ( .Q(g6338), .DIN1(n2553), .DIN2(n2554) );
nnd2s1 U3142 ( .Q(n2554), .DIN1(g381), .DIN2(n2531) );
nnd2s1 U3143 ( .Q(n2553), .DIN1(g374), .DIN2(n2532) );
nnd2s1 U3144 ( .Q(g6337), .DIN1(n2555), .DIN2(n2556) );
nnd2s1 U3145 ( .Q(n2556), .DIN1(g378), .DIN2(n2531) );
nnd2s1 U3146 ( .Q(n2555), .DIN1(g373), .DIN2(n2532) );
hi1s1 U3147 ( .Q(n2532), .DIN(n2531) );
nnd2s1 U3148 ( .Q(n2531), .DIN1(g452), .DIN2(DFF_171net396) );
nnd2s1 U3149 ( .Q(g6336), .DIN1(n2557), .DIN2(n2558) );
nnd2s1 U3150 ( .Q(n2558), .DIN1(g359), .DIN2(n2559) );
nnd2s1 U3151 ( .Q(n2557), .DIN1(g355), .DIN2(n2560) );
nnd2s1 U3152 ( .Q(g6335), .DIN1(n2561), .DIN2(n2562) );
nnd2s1 U3153 ( .Q(n2562), .DIN1(g356), .DIN2(n2559) );
nnd2s1 U3154 ( .Q(n2561), .DIN1(g354), .DIN2(n2560) );
nnd2s1 U3155 ( .Q(g6334), .DIN1(n2563), .DIN2(n2564) );
nnd2s1 U3156 ( .Q(n2564), .DIN1(g333), .DIN2(n2559) );
nnd2s1 U3157 ( .Q(n2563), .DIN1(g317), .DIN2(n2560) );
nnd2s1 U3158 ( .Q(g6333), .DIN1(n2565), .DIN2(n2566) );
nnd2s1 U3159 ( .Q(n2566), .DIN1(g330), .DIN2(n2559) );
nnd2s1 U3160 ( .Q(n2565), .DIN1(g316), .DIN2(n2560) );
nnd2s1 U3161 ( .Q(g6332), .DIN1(n2567), .DIN2(n2568) );
nnd2s1 U3162 ( .Q(n2568), .DIN1(g327), .DIN2(n2559) );
nnd2s1 U3163 ( .Q(n2567), .DIN1(g315), .DIN2(n2560) );
nnd2s1 U3164 ( .Q(g6331), .DIN1(n2569), .DIN2(n2570) );
nnd2s1 U3165 ( .Q(n2570), .DIN1(g324), .DIN2(n2559) );
nnd2s1 U3166 ( .Q(n2569), .DIN1(g314), .DIN2(n2560) );
nnd2s1 U3167 ( .Q(g6330), .DIN1(n2571), .DIN2(n2572) );
nnd2s1 U3168 ( .Q(n2572), .DIN1(g321), .DIN2(n2559) );
nnd2s1 U3169 ( .Q(n2571), .DIN1(g313), .DIN2(n2560) );
nnd2s1 U3170 ( .Q(g6329), .DIN1(n2573), .DIN2(n2574) );
nnd2s1 U3171 ( .Q(n2574), .DIN1(g318), .DIN2(n2559) );
nnd2s1 U3172 ( .Q(n2573), .DIN1(g312), .DIN2(n2560) );
nnd2s1 U3173 ( .Q(g6328), .DIN1(n2575), .DIN2(n2576) );
nnd2s1 U3174 ( .Q(n2576), .DIN1(g309), .DIN2(n2559) );
nnd2s1 U3175 ( .Q(n2575), .DIN1(g296), .DIN2(n2560) );
nnd2s1 U3176 ( .Q(g6327), .DIN1(n2577), .DIN2(n2578) );
nnd2s1 U3177 ( .Q(n2578), .DIN1(g306), .DIN2(n2559) );
nnd2s1 U3178 ( .Q(n2577), .DIN1(g295), .DIN2(n2560) );
nnd2s1 U3179 ( .Q(g6326), .DIN1(n2579), .DIN2(n2580) );
nnd2s1 U3180 ( .Q(n2580), .DIN1(g303), .DIN2(n2559) );
nnd2s1 U3181 ( .Q(n2579), .DIN1(g294), .DIN2(n2560) );
nnd2s1 U3182 ( .Q(g6325), .DIN1(n2581), .DIN2(n2582) );
nnd2s1 U3183 ( .Q(n2582), .DIN1(g300), .DIN2(n2559) );
nnd2s1 U3184 ( .Q(n2581), .DIN1(g293), .DIN2(n2560) );
nnd2s1 U3185 ( .Q(g6324), .DIN1(n2583), .DIN2(n2584) );
nnd2s1 U3186 ( .Q(n2584), .DIN1(g297), .DIN2(n2559) );
nnd2s1 U3187 ( .Q(n2583), .DIN1(g292), .DIN2(n2560) );
hi1s1 U3188 ( .Q(n2560), .DIN(n2559) );
nnd2s1 U3189 ( .Q(n2559), .DIN1(g371), .DIN2(DFF_365net590) );
nnd2s1 U3190 ( .Q(g6323), .DIN1(n2585), .DIN2(n2586) );
nnd2s1 U3191 ( .Q(n2586), .DIN1(g278), .DIN2(n2587) );
nnd2s1 U3192 ( .Q(n2585), .DIN1(g274), .DIN2(n2588) );
nnd2s1 U3193 ( .Q(g6322), .DIN1(n2589), .DIN2(n2590) );
nnd2s1 U3194 ( .Q(n2590), .DIN1(g275), .DIN2(n2587) );
nnd2s1 U3195 ( .Q(n2589), .DIN1(g273), .DIN2(n2588) );
nnd2s1 U3196 ( .Q(g6321), .DIN1(n2591), .DIN2(n2592) );
nnd2s1 U3197 ( .Q(n2592), .DIN1(g252), .DIN2(n2587) );
nnd2s1 U3198 ( .Q(n2591), .DIN1(g236), .DIN2(n2588) );
nnd2s1 U3199 ( .Q(g6320), .DIN1(n2593), .DIN2(n2594) );
nnd2s1 U3200 ( .Q(n2594), .DIN1(g249), .DIN2(n2587) );
nnd2s1 U3201 ( .Q(n2593), .DIN1(g235), .DIN2(n2588) );
nnd2s1 U3202 ( .Q(g6319), .DIN1(n2595), .DIN2(n2596) );
nnd2s1 U3203 ( .Q(n2596), .DIN1(g246), .DIN2(n2587) );
nnd2s1 U3204 ( .Q(n2595), .DIN1(g234), .DIN2(n2588) );
nnd2s1 U3205 ( .Q(g6318), .DIN1(n2597), .DIN2(n2598) );
nnd2s1 U3206 ( .Q(n2598), .DIN1(g243), .DIN2(n2587) );
nnd2s1 U3207 ( .Q(n2597), .DIN1(g233), .DIN2(n2588) );
nnd2s1 U3208 ( .Q(g6317), .DIN1(n2599), .DIN2(n2600) );
nnd2s1 U3209 ( .Q(n2600), .DIN1(g240), .DIN2(n2587) );
nnd2s1 U3210 ( .Q(n2599), .DIN1(g232), .DIN2(n2588) );
nnd2s1 U3211 ( .Q(g6316), .DIN1(n2601), .DIN2(n2602) );
nnd2s1 U3212 ( .Q(n2602), .DIN1(g237), .DIN2(n2587) );
nnd2s1 U3213 ( .Q(n2601), .DIN1(g231), .DIN2(n2588) );
nnd2s1 U3214 ( .Q(g6315), .DIN1(n2603), .DIN2(n2604) );
nnd2s1 U3215 ( .Q(n2604), .DIN1(g228), .DIN2(n2587) );
nnd2s1 U3216 ( .Q(n2603), .DIN1(g215), .DIN2(n2588) );
nnd2s1 U3217 ( .Q(g6314), .DIN1(n2605), .DIN2(n2606) );
nnd2s1 U3218 ( .Q(n2606), .DIN1(g225), .DIN2(n2587) );
nnd2s1 U3219 ( .Q(n2605), .DIN1(g214), .DIN2(n2588) );
nnd2s1 U3220 ( .Q(g6313), .DIN1(n2607), .DIN2(n2608) );
nnd2s1 U3221 ( .Q(n2608), .DIN1(g222), .DIN2(n2587) );
nnd2s1 U3222 ( .Q(n2607), .DIN1(g213), .DIN2(n2588) );
nnd2s1 U3223 ( .Q(g6312), .DIN1(n2609), .DIN2(n2610) );
nnd2s1 U3224 ( .Q(n2610), .DIN1(g219), .DIN2(n2587) );
nnd2s1 U3225 ( .Q(n2609), .DIN1(g212), .DIN2(n2588) );
nnd2s1 U3226 ( .Q(g6311), .DIN1(n2611), .DIN2(n2612) );
nnd2s1 U3227 ( .Q(n2612), .DIN1(g216), .DIN2(n2587) );
nnd2s1 U3228 ( .Q(n2611), .DIN1(g211), .DIN2(n2588) );
hi1s1 U3229 ( .Q(n2588), .DIN(n2587) );
nnd2s1 U3230 ( .Q(n2587), .DIN1(g290), .DIN2(DFF_342net567) );
nor4s1 U3231 ( .Q(g6056), .DIN1(g889), .DIN2(g778), .DIN3(n2613), .DIN4(n2614) );
hi1s1 U3232 ( .Q(n2614), .DIN(n2360) );
nor2s1 U3233 ( .Q(n2360), .DIN1(g887), .DIN2(g888) );
nor2s1 U3234 ( .Q(n2613), .DIN1(n2615), .DIN2(n2616) );
nnd4s1 U3235 ( .Q(n2616), .DIN1(n2617), .DIN2(n2618), .DIN3(n2619), .DIN4(n2620) );
xor2s1 U3236 ( .Q(n2620), .DIN1(g840), .DIN2(n1421) );
xor2s1 U3237 ( .Q(n2619), .DIN1(g837), .DIN2(n1394) );
xor2s1 U3238 ( .Q(n2618), .DIN1(g834), .DIN2(n1382) );
xor2s1 U3239 ( .Q(n2617), .DIN1(g831), .DIN2(n1379) );
nnd4s1 U3240 ( .Q(n2615), .DIN1(n2621), .DIN2(n2622), .DIN3(n2623), .DIN4(n2624) );
xor2s1 U3241 ( .Q(n2624), .DIN1(g852), .DIN2(n1423) );
xor2s1 U3242 ( .Q(n2623), .DIN1(g849), .DIN2(n1395) );
xor2s1 U3243 ( .Q(n2622), .DIN1(g846), .DIN2(n1383) );
xor2s1 U3244 ( .Q(n2621), .DIN1(g843), .DIN2(n1380) );
nnd2s1 U3245 ( .Q(g5746), .DIN1(n2625), .DIN2(n1389) );
xor2s1 U3246 ( .Q(n2625), .DIN1(n2626), .DIN2(DFF_166net391) );
nor2s1 U3247 ( .Q(n2626), .DIN1(g33), .DIN2(n2627) );
nnd2s1 U3248 ( .Q(g5745), .DIN1(g5180), .DIN2(n2628) );
or3s1 U3249 ( .Q(n2628), .DIN1(g1430), .DIN2(g1431), .DIN3(n1466) );
nnd2s1 U3250 ( .Q(g5744), .DIN1(g5177), .DIN2(n2629) );
or3s1 U3251 ( .Q(n2629), .DIN1(g1428), .DIN2(g1429), .DIN3(n1467) );
nnd2s1 U3252 ( .Q(g5743), .DIN1(n2630), .DIN2(n2631) );
nnd2s1 U3253 ( .Q(n2631), .DIN1(n2632), .DIN2(n1504) );
xor2s1 U3254 ( .Q(n2632), .DIN1(g1317), .DIN2(g1313) );
nnd2s1 U3255 ( .Q(n2630), .DIN1(g141), .DIN2(g1329) );
nnd2s1 U3256 ( .Q(g5742), .DIN1(n2633), .DIN2(n2634) );
nnd2s1 U3257 ( .Q(n2634), .DIN1(g145), .DIN2(g1329) );
or2s1 U3258 ( .Q(n2633), .DIN1(g1313), .DIN2(n1505) );
hi1s1 U3259 ( .Q(g5741), .DIN(n2211) );
nnd3s1 U3260 ( .Q(n2211), .DIN1(g3847), .DIN2(n2295), .DIN3(g3848) );
hi1s1 U3261 ( .Q(n2295), .DIN(n2294) );
nnd3s1 U3262 ( .Q(n2294), .DIN1(g3850), .DIN2(n2214), .DIN3(g3851) );
and4s1 U3263 ( .Q(n2214), .DIN1(g3852), .DIN2(g3846), .DIN3(g3845), .DIN4(g3844) );
nnd4s1 U3264 ( .Q(g5740), .DIN1(n1495), .DIN2(n1485), .DIN3(n1502), .DIN4(n1486) );
and3s1 U3265 ( .Q(g5739), .DIN1(n1494), .DIN2(n1513), .DIN3(n2400) );
and3s1 U3266 ( .Q(g5738), .DIN1(n2400), .DIN2(n1494), .DIN3(n1514) );
and3s1 U3267 ( .Q(g5737), .DIN1(n2400), .DIN2(n1513), .DIN3(n1495) );
and2s1 U3268 ( .Q(n2400), .DIN1(n1485), .DIN2(n2458) );
nor2s1 U3269 ( .Q(n2458), .DIN1(n1486), .DIN2(n1502) );
and3s1 U3270 ( .Q(g5736), .DIN1(n2635), .DIN2(n2464), .DIN3(g1254) );
nnd3s1 U3271 ( .Q(n2464), .DIN1(n1495), .DIN2(n1485), .DIN3(n1514) );
nnd2s1 U3272 ( .Q(n2635), .DIN1(n2636), .DIN2(n2637) );
or2s1 U3273 ( .Q(n2637), .DIN1(n1494), .DIN2(g5173) );
nnd2s1 U3274 ( .Q(n2636), .DIN1(n1485), .DIN2(n1400) );
nor2s1 U3275 ( .Q(g5735), .DIN1(n2638), .DIN2(n2639) );
hi1s1 U3276 ( .Q(n2639), .DIN(g2801) );
nor2s1 U3277 ( .Q(g5733), .DIN1(n2640), .DIN2(n1404) );
nor2s1 U3278 ( .Q(n2640), .DIN1(g5161), .DIN2(n2641) );
xor2s1 U3279 ( .Q(n2641), .DIN1(g3849), .DIN2(g210) );
nor2s1 U3280 ( .Q(g5732), .DIN1(n2642), .DIN2(n1404) );
nor2s1 U3281 ( .Q(n2642), .DIN1(g5160), .DIN2(n2643) );
xor2s1 U3282 ( .Q(n2643), .DIN1(g3842), .DIN2(g205) );
nor2s1 U3283 ( .Q(g5731), .DIN1(n2644), .DIN2(n1404) );
nor2s1 U3284 ( .Q(n2644), .DIN1(g5159), .DIN2(n2645) );
xor2s1 U3285 ( .Q(n2645), .DIN1(g3836), .DIN2(g195) );
nor2s1 U3286 ( .Q(g5730), .DIN1(n2646), .DIN2(n1404) );
nor2s1 U3287 ( .Q(n2646), .DIN1(g5158), .DIN2(n2647) );
xor2s1 U3288 ( .Q(n2647), .DIN1(g3838), .DIN2(g186) );
nnd2s1 U3289 ( .Q(g5187), .DIN1(n2648), .DIN2(n2649) );
nnd3s1 U3290 ( .Q(n2649), .DIN1(n2650), .DIN2(n1392), .DIN3(g1454) );
nnd2s1 U3291 ( .Q(n2648), .DIN1(g1450), .DIN2(n2651) );
nnd2s1 U3292 ( .Q(g5186), .DIN1(n2652), .DIN2(n2653) );
nnd2s1 U3293 ( .Q(n2653), .DIN1(n2651), .DIN2(n1415) );
hi1s1 U3294 ( .Q(n2651), .DIN(g5185) );
nnd4s1 U3295 ( .Q(n2652), .DIN1(n1452), .DIN2(n1392), .DIN3(n2650), .DIN4(g1450) );
nnd3s1 U3296 ( .Q(g5185), .DIN1(n2650), .DIN2(n1392), .DIN3(g1444) );
nnd2s1 U3297 ( .Q(n2650), .DIN1(g1454), .DIN2(g1450) );
nnd2s1 U3298 ( .Q(g5184), .DIN1(n2654), .DIN2(n1389) );
xor2s1 U3299 ( .Q(n2654), .DIN1(g33), .DIN2(n2627) );
nnd2s1 U3300 ( .Q(g5183), .DIN1(n2655), .DIN2(n2656) );
nnd3s1 U3301 ( .Q(n2656), .DIN1(g1432), .DIN2(n1389), .DIN3(n2627) );
nnd2s1 U3302 ( .Q(n2655), .DIN1(g1439), .DIN2(n2657) );
hi1s1 U3303 ( .Q(n2657), .DIN(g5181) );
nnd2s1 U3304 ( .Q(g5182), .DIN1(n2658), .DIN2(n2659) );
or2s1 U3305 ( .Q(n2659), .DIN1(g5181), .DIN2(g1439) );
nnd4s1 U3306 ( .Q(n2658), .DIN1(n1458), .DIN2(n1389), .DIN3(n2627), .DIN4(g1439) );
nnd3s1 U3307 ( .Q(g5181), .DIN1(n2627), .DIN2(n1389), .DIN3(g1435) );
nnd2s1 U3308 ( .Q(n2627), .DIN1(g1439), .DIN2(g1432) );
or3s1 U3309 ( .Q(g5180), .DIN1(g1430), .DIN2(g1431), .DIN3(g1412) );
and3s1 U3310 ( .Q(g5179), .DIN1(n1448), .DIN2(n1399), .DIN3(g1416) );
nnd2s1 U3311 ( .Q(g5178), .DIN1(n2660), .DIN2(n2661) );
nnd2s1 U3312 ( .Q(n2661), .DIN1(g1409), .DIN2(g1416) );
nnd2s1 U3313 ( .Q(n2660), .DIN1(g2474), .DIN2(n1398) );
or3s1 U3314 ( .Q(g5177), .DIN1(g1428), .DIN2(g1429), .DIN3(g1405) );
hi1s1 U3315 ( .Q(g5176), .DIN(n2452) );
nnd2s1 U3316 ( .Q(n2452), .DIN1(g154), .DIN2(n1401) );
or2s1 U3317 ( .Q(g5175), .DIN1(n2662), .DIN2(n2663) );
nnd4s1 U3318 ( .Q(n2663), .DIN1(n1480), .DIN2(n1488), .DIN3(n1506), .DIN4(n1490) );
or4s1 U3319 ( .Q(n2662), .DIN1(n1478), .DIN2(n1483), .DIN3(n1509), .DIN4(n1493) );
nnd2s1 U3320 ( .Q(g5174), .DIN1(n2664), .DIN2(n1400) );
xor2s1 U3321 ( .Q(n2664), .DIN1(n1494), .DIN2(n1514) );
nnd2s1 U3322 ( .Q(g5173), .DIN1(n1514), .DIN2(n1400) );
nnd4s1 U3323 ( .Q(g5172), .DIN1(n1396), .DIN2(DFF_630net855), .DIN3(n1456), .DIN4(n2665) );
and3s1 U3324 ( .Q(n2665), .DIN1(DFF_66net291), .DIN2(DFF_517net742), .DIN3(DFF_313net538) );
nor2s1 U3325 ( .Q(g5170), .DIN1(n2638), .DIN2(n2666) );
nor2s1 U3326 ( .Q(n2666), .DIN1(n2667), .DIN2(g945) );
and2s1 U3327 ( .Q(n2667), .DIN1(g955), .DIN2(g959) );
and3s1 U3328 ( .Q(n2638), .DIN1(g945), .DIN2(g955), .DIN3(g959) );
xor2s1 U3329 ( .Q(g5169), .DIN1(g959), .DIN2(g955) );
nor2s1 U3330 ( .Q(g5168), .DIN1(n2668), .DIN2(DFF_391net616) );
and2s1 U3331 ( .Q(n2668), .DIN1(n1426), .DIN2(g940) );
nor2s1 U3332 ( .Q(g5167), .DIN1(g4654), .DIN2(n2669) );
nor2s1 U3333 ( .Q(n2669), .DIN1(n2670), .DIN2(g871) );
and2s1 U3334 ( .Q(n2670), .DIN1(g929), .DIN2(g933) );
xor2s1 U3335 ( .Q(g5166), .DIN1(g933), .DIN2(g929) );
and3s1 U3336 ( .Q(g5165), .DIN1(g888), .DIN2(n2370), .DIN3(g4316) );
nor2s1 U3337 ( .Q(n2370), .DIN1(n1432), .DIN2(g889) );
nor2s1 U3338 ( .Q(g5163), .DIN1(g4316), .DIN2(n1457) );
and3s1 U3339 ( .Q(g4669), .DIN1(g1454), .DIN2(n1415), .DIN3(g1444) );
nor3s1 U3340 ( .Q(g4668), .DIN1(g1444), .DIN2(g1454), .DIN3(n1415) );
nnd2s1 U3341 ( .Q(g4665), .DIN1(n1399), .DIN2(n2671) );
nnd2s1 U3342 ( .Q(n2671), .DIN1(n1398), .DIN2(n1448) );
nor4s1 U3343 ( .Q(g4658), .DIN1(n2672), .DIN2(n2673), .DIN3(n2674), .DIN4(n2675) );
nnd3s1 U3344 ( .Q(n2675), .DIN1(DFF_422net647), .DIN2(DFF_63net288), .DIN3(DFF_412net637) );
nnd3s1 U3345 ( .Q(n2674), .DIN1(DFF_601net826), .DIN2(DFF_215net440), .DIN3(DFF_635net860) );
nnd3s1 U3346 ( .Q(n2673), .DIN1(DFF_260net485), .DIN2(DFF_24net249), .DIN3(DFF_68net293) );
nnd4s1 U3347 ( .Q(n2672), .DIN1(DFF_140net365), .DIN2(DFF_518net743), .DIN3(DFF_527net752), .DIN4(DFF_180net405) );
nor2s1 U3348 ( .Q(g4656), .DIN1(g1269), .DIN2(g1268) );
hi1s1 U3349 ( .Q(g4654), .DIN(n2364) );
nnd3s1 U3350 ( .Q(n2364), .DIN1(g871), .DIN2(g929), .DIN3(g933) );
and3s1 U3351 ( .Q(g4302), .DIN1(g889), .DIN2(g887), .DIN3(g888) );
nnd2s1 U3352 ( .Q(g3861), .DIN1(DFF_175net400), .DIN2(DFF_98net323) );
hi1s1 U3353 ( .Q(g3856), .DIN(g929) );
nor2s1 U3354 ( .Q(g3555), .DIN1(g1398), .DIN2(DFF_218net443) );
nor2s1 U3355 ( .Q(g3528), .DIN1(g1391), .DIN2(DFF_402net627) );
nor2s1 U3356 ( .Q(g3516), .DIN1(g1401), .DIN2(DFF_252net477) );
nor2s1 U3357 ( .Q(g3505), .DIN1(g1395), .DIN2(DFF_377net602) );
nor4s1 U3358 ( .Q(g3504), .DIN1(n2676), .DIN2(n2677), .DIN3(n2678), .DIN4(n2679) );
nnd3s1 U3359 ( .Q(n2679), .DIN1(DFF_84net309), .DIN2(DFF_200net425), .DIN3(DFF_314net539) );
nnd3s1 U3360 ( .Q(n2678), .DIN1(DFF_578net803), .DIN2(DFF_236net461), .DIN3(DFF_564net789) );
nnd3s1 U3361 ( .Q(n2677), .DIN1(DFF_521net746), .DIN2(DFF_101net326), .DIN3(DFF_159net384) );
nnd4s1 U3362 ( .Q(n2676), .DIN1(DFF_619net844), .DIN2(DFF_155net380), .DIN3(DFF_597net822), .DIN4(DFF_20net245) );
hi1s1 U3363 ( .Q(g3084), .DIN(g955) );
nnd2s1 U3364 ( .Q(g2801), .DIN1(n2086), .DIN2(n2680) );
nnd2s1 U3365 ( .Q(n2680), .DIN1(g940), .DIN2(n1426) );
hi1s1 U3366 ( .Q(n2086), .DIN(n2087) );
nor2s1 U3367 ( .Q(n2087), .DIN1(n1426), .DIN2(g940) );
nnd2s1 U3368 ( .Q(g2474), .DIN1(g1412), .DIN2(g1405) );
hi1s1 U3369 ( .Q(g1683), .DIN(g795) );
hi1s1 U3370 ( .Q(I5528), .DIN(g6851) );
hi1s1 U3499 ( .Q(n1431), .DIN(g71) );
hi1s1 U3500 ( .Q(n1456), .DIN(g1179) );
hi1s1 U3501 ( .Q(n1415), .DIN(g1450) );
hi1s1 U3502 ( .Q(DFF_630net855), .DIN(g4370) );
hi1s1 U3503 ( .Q(n1465), .DIN(g866) );
hi1s1 U3504 ( .Q(n1407), .DIN(g1158) );
hi1s1 U3505 ( .Q(n1451), .DIN(g1519) );
hi1s1 U3506 ( .Q(n1459), .DIN(g1057) );
hi1s1 U3507 ( .Q(n1474), .DIN(g1318) );
hi1s1 U3508 ( .Q(DFF_576net801), .DIN(g7423) );
hi1s1 U3509 ( .Q(n1453), .DIN(g1118) );
hi1s1 U3510 ( .Q(n1429), .DIN(n1387) );
hi1s1 U3511 ( .Q(g3863), .DIN(g2661) );
hi1s1 U3512 ( .Q(n1424), .DIN(g1348) );
hi1s1 U3513 ( .Q(n1411), .DIN(g1330) );
hi1s1 U3514 ( .Q(n1461), .DIN(g1130) );
hi1s1 U3515 ( .Q(DFF_550net775), .DIN(g2844) );
hi1s1 U3516 ( .Q(n1419), .DIN(g4659) );
hi1s1 U3517 ( .Q(n1398), .DIN(g1416) );
hi1s1 U3518 ( .Q(n1492), .DIN(g4646) );
hi1s1 U3519 ( .Q(DFF_517net742), .DIN(g4373) );
hi1s1 U3520 ( .Q(n1494), .DIN(g4650) );
hi1s1 U3521 ( .Q(n1462), .DIN(g1149) );
hi1s1 U3522 ( .Q(n1504), .DIN(g1329) );
hi1s1 U3523 ( .Q(n1457), .DIN(g874) );
hi1s1 U3524 ( .Q(n1430), .DIN(g1354) );
hi1s1 U3525 ( .Q(n1402), .DIN(g1097) );
hi1s1 U3526 ( .Q(n1445), .DIN(g1944) );
hi1s1 U3527 ( .Q(n1410), .DIN(g1342) );
hi1s1 U3528 ( .Q(n1480), .DIN(g4639) );
hi1s1 U3529 ( .Q(n1506), .DIN(g4641) );
hi1s1 U3530 ( .Q(n1440), .DIN(g1065) );
hi1s1 U3531 ( .Q(n1420), .DIN(g1336) );
hi1s1 U3532 ( .Q(n1383), .DIN(g2646) );
hi1s1 U3533 ( .Q(n1513), .DIN(g4651) );
hi1s1 U3534 ( .Q(n1405), .DIN(g888) );
hi1s1 U3535 ( .Q(n1470), .DIN(g1069) );
hi1s1 U3536 ( .Q(n1396), .DIN(g4267) );
hi1s1 U3537 ( .Q(n1482), .DIN(g4644) );
hi1s1 U3538 ( .Q(n1394), .DIN(g2649) );
hi1s1 U3539 ( .Q(DFF_404net629), .DIN(g5146) );
hi1s1 U3540 ( .Q(n1488), .DIN(g4640) );
hi1s1 U3541 ( .Q(n1423), .DIN(g2644) );
hi1s1 U3542 ( .Q(n1455), .DIN(g1489) );
hi1s1 U3543 ( .Q(n1382), .DIN(g2650) );
hi1s1 U3544 ( .Q(DFF_373net598), .DIN(g5571) );
hi1s1 U3545 ( .Q(n1484), .DIN(g4649) );
hi1s1 U3546 ( .Q(n1471), .DIN(g855) );
hi1s1 U3547 ( .Q(DFF_365net590), .DIN(g3130) );
hi1s1 U3548 ( .Q(n1468), .DIN(g3855) );
hi1s1 U3549 ( .Q(n1458), .DIN(g1435) );
hi1s1 U3550 ( .Q(n1432), .DIN(g887) );
hi1s1 U3551 ( .Q(n1511), .DIN(g6841) );
hi1s1 U3552 ( .Q(n1508), .DIN(g4645) );
hi1s1 U3553 ( .Q(DFF_342net567), .DIN(g3096) );
hi1s1 U3554 ( .Q(n1414), .DIN(n1385) );
hi1s1 U3555 ( .Q(n1449), .DIN(g3845) );
hi1s1 U3556 ( .Q(n1475), .DIN(g2653) );
hi1s1 U3557 ( .Q(n1397), .DIN(g68) );
hi1s1 U3558 ( .Q(g6675), .DIN(g1432) );
hi1s1 U3559 ( .Q(DFF_313net538), .DIN(g4371) );
hi1s1 U3560 ( .Q(n1391), .DIN(g74) );
hi1s1 U3561 ( .Q(n1416), .DIN(g815) );
hi1s1 U3562 ( .Q(n1388), .DIN(g62) );
hi1s1 U3563 ( .Q(n1496), .DIN(g6843) );
hi1s1 U3564 ( .Q(DFF_286net511), .DIN(g3191) );
hi1s1 U3565 ( .Q(n1401), .DIN(g4599) );
hi1s1 U3566 ( .Q(n1469), .DIN(g859) );
hi1s1 U3567 ( .Q(DFF_270net495), .DIN(g5145) );
hi1s1 U3568 ( .Q(n1473), .DIN(g1327) );
hi1s1 U3569 ( .Q(n1409), .DIN(g77) );
hi1s1 U3570 ( .Q(n1418), .DIN(g158) );
hi1s1 U3571 ( .Q(n1502), .DIN(g4647) );
hi1s1 U3572 ( .Q(n1464), .DIN(g990) );
hi1s1 U3573 ( .Q(n1433), .DIN(g1018) );
hi1s1 U3574 ( .Q(n1390), .DIN(g1333) );
hi1s1 U3575 ( .Q(n1486), .DIN(g4648) );
hi1s1 U3576 ( .Q(n1403), .DIN(g1247) );
hi1s1 U3577 ( .Q(DFF_175net400), .DIN(g2664) );
hi1s1 U3578 ( .Q(DFF_171net396), .DIN(g3159) );
hi1s1 U3579 ( .Q(n1490), .DIN(g4642) );
hi1s1 U3580 ( .Q(DFF_166net391), .DIN(g38) );
hi1s1 U3581 ( .Q(n1460), .DIN(g1045) );
hi1s1 U3582 ( .Q(n1477), .DIN(g4643) );
hi1s1 U3583 ( .Q(n1380), .DIN(g2647) );
hi1s1 U3584 ( .Q(n1472), .DIN(g822) );
hi1s1 U3585 ( .Q(n1428), .DIN(n1384) );
hi1s1 U3586 ( .Q(n1454), .DIN(g1098) );
hi1s1 U3587 ( .Q(n1417), .DIN(g889) );
hi1s1 U3588 ( .Q(n1393), .DIN(g985) );
hi1s1 U3589 ( .Q(n1446), .DIN(g1029) );
hi1s1 U3590 ( .Q(n1412), .DIN(n1386) );
hi1s1 U3591 ( .Q(n1413), .DIN(n1381) );
hi1s1 U3592 ( .Q(DFF_66net291), .DIN(g4372) );
hi1s1 U3593 ( .Q(n1379), .DIN(g2651) );
hi1s1 U3594 ( .Q(n1421), .DIN(g2648) );
hi1s1 U3595 ( .Q(n1463), .DIN(g803) );
hi1s1 U3596 ( .Q(n1452), .DIN(g1444) );
hi1s1 U3597 ( .Q(n1444), .DIN(g80) );
hi1s1 U3598 ( .Q(n1422), .DIN(g1304) );
hi1s1 U3599 ( .Q(n1395), .DIN(g2645) );
hi1s1 U3600 ( .Q(n1400), .DIN(g2659) );
hi1s1 U3601 ( .Q(n1399), .DIN(g2672) );
hi1s1 U3602 ( .Q(n1408), .DIN(g1339) );
hi1s1 U3603 ( .Q(n1441), .DIN(g1092) );
endmodule